
library work;
use work.extra_types.all;
use work.dpath_components.all;

entity start_dp is
  port(
    ip : in  bit_vector(276 downto 1);
    op : out bit_vector(273 downto 1) := (others => '0');

    load_reqs : out bit_vector(23 downto 0) := (others => '0');
    load_acks : in bit_vector(23 downto 0);
    load_addr : out MemoryBusVectorType(23 downto 0);
    load_data : in  MemoryBusVectorType(23 downto 0);

    store_reqs : out bit_vector(15 downto 0) := (others => '0');
    store_acks : in bit_vector(15 downto 0);
    store_addr : out MemoryBusVectorType(15 downto 0);
    store_data : out MemoryBusVectorType(15 downto 0);

    reset : in bit;
    clk   : in  bit);
end start_dp;

architecture Behavioral of start_dp is

  signal cst_0_uint_d_wire : bit_vector(31 downto 0);
  signal cst_10_uint_d_wire : bit_vector(31 downto 0);
  signal cst_11_int_d_wire : bit_vector(31 downto 0);
  signal cst_12_uint_d_wire : bit_vector(31 downto 0);
  signal cst_13_uint_d_wire : bit_vector(31 downto 0);
  signal cst_14_int_d_wire : bit_vector(31 downto 0);
  signal cst_15_int_d_wire : bit_vector(31 downto 0);
  signal cst_16_uint_d_wire : bit_vector(31 downto 0);
  signal cst_17_int_d_wire : bit_vector(31 downto 0);
  signal cst_18_int_d_wire : bit_vector(31 downto 0);
  signal cst_19_uint_d_wire : bit_vector(31 downto 0);
  signal cst_1_uint_d_wire : bit_vector(31 downto 0);
  signal cst_20_uint_d_wire : bit_vector(31 downto 0);
  signal cst_21_uint_d_wire : bit_vector(31 downto 0);
  signal cst_22_int_d_wire : bit_vector(31 downto 0);
  signal cst_23_int_d_wire : bit_vector(31 downto 0);
  signal cst_24_uint_d_wire : bit_vector(31 downto 0);
  signal cst_25_uint_d_wire : bit_vector(31 downto 0);
  signal cst_26_uint_d_wire : bit_vector(31 downto 0);
  signal cst_27_uint_d_wire : bit_vector(31 downto 0);
  signal cst_28_uint_d_wire : bit_vector(31 downto 0);
  signal cst_29_uint_d_wire : bit_vector(31 downto 0);
  signal cst_2_uint_d_wire : bit_vector(31 downto 0);
  signal cst_30_int_d_wire : bit_vector(31 downto 0);
  signal cst_31_uint_d_wire : bit_vector(31 downto 0);
  signal cst_32_uint_d_wire : bit_vector(31 downto 0);
  signal cst_33_uint_d_wire : bit_vector(31 downto 0);
  signal cst_34_int_d_wire : bit_vector(31 downto 0);
  signal cst_35_uint_d_wire : bit_vector(31 downto 0);
  signal cst_36_int_d_wire : bit_vector(31 downto 0);
  signal cst_37_int_d_wire : bit_vector(31 downto 0);
  signal cst_38_uint_d_wire : bit_vector(31 downto 0);
  signal cst_39_uint_d_wire : bit_vector(31 downto 0);
  signal cst_3_float_d_wire : bit_vector(31 downto 0);
  signal cst_40_int_d_wire : bit_vector(31 downto 0);
  signal cst_41_int_d_wire : bit_vector(31 downto 0);
  signal cst_42_uint_d_wire : bit_vector(31 downto 0);
  signal cst_43_uint_d_wire : bit_vector(31 downto 0);
  signal cst_44_uint_d_wire : bit_vector(31 downto 0);
  signal cst_45_uint_d_wire : bit_vector(31 downto 0);
  signal cst_46_uint_d_wire : bit_vector(31 downto 0);
  signal cst_47_int_d_wire : bit_vector(31 downto 0);
  signal cst_48_int_d_wire : bit_vector(31 downto 0);
  signal cst_49_uint_d_wire : bit_vector(31 downto 0);
  signal cst_4_uint_d_wire : bit_vector(31 downto 0);
  signal cst_50_uint_d_wire : bit_vector(31 downto 0);
  signal cst_51_uint_d_wire : bit_vector(31 downto 0);
  signal cst_52_int_d_wire : bit_vector(31 downto 0);
  signal cst_53_uint_d_wire : bit_vector(31 downto 0);
  signal cst_54_uint_d_wire : bit_vector(31 downto 0);
  signal cst_55_uint_d_wire : bit_vector(31 downto 0);
  signal cst_56_float_d_wire : bit_vector(31 downto 0);
  signal cst_57_int_d_wire : bit_vector(31 downto 0);
  signal cst_58_int_d_wire : bit_vector(31 downto 0);
  signal cst_59_uint_d_wire : bit_vector(31 downto 0);
  signal cst_5_uint_d_wire : bit_vector(31 downto 0);
  signal cst_60_float_d_wire : bit_vector(31 downto 0);
  signal cst_61_uint_d_wire : bit_vector(31 downto 0);
  signal cst_62_uint_d_wire : bit_vector(31 downto 0);
  signal cst_63_int_d_wire : bit_vector(31 downto 0);
  signal cst_64_int_d_wire : bit_vector(31 downto 0);
  signal cst_65_float_d_wire : bit_vector(31 downto 0);
  signal cst_66_uint_d_wire : bit_vector(31 downto 0);
  signal cst_67_uint_d_wire : bit_vector(31 downto 0);
  signal cst_68_int_d_wire : bit_vector(31 downto 0);
  signal cst_69_int_d_wire : bit_vector(31 downto 0);
  signal cst_6_uint_d_wire : bit_vector(31 downto 0);
  signal cst_70_uint_d_wire : bit_vector(31 downto 0);
  signal cst_71_uint_d_wire : bit_vector(31 downto 0);
  signal cst_72_uint_d_wire : bit_vector(31 downto 0);
  signal cst_73_int_d_wire : bit_vector(31 downto 0);
  signal cst_74_uint_d_wire : bit_vector(31 downto 0);
  signal cst_75_uint_d_wire : bit_vector(31 downto 0);
  signal cst_76_uint_d_wire : bit_vector(31 downto 0);
  signal cst_77_int_d_wire : bit_vector(31 downto 0);
  signal cst_78_uint_d_wire : bit_vector(31 downto 0);
  signal cst_79_int_d_wire : bit_vector(31 downto 0);
  signal cst_7_uint_d_wire : bit_vector(31 downto 0);
  signal cst_80_uint_d_wire : bit_vector(31 downto 0);
  signal cst_81_uint_d_wire : bit_vector(31 downto 0);
  signal cst_82_uint_d_wire : bit_vector(31 downto 0);
  signal cst_83_int_d_wire : bit_vector(31 downto 0);
  signal cst_84_int_d_wire : bit_vector(31 downto 0);
  signal cst_85_uint_d_wire : bit_vector(31 downto 0);
  signal cst_86_uint_d_wire : bit_vector(31 downto 0);
  signal cst_87_int_d_wire : bit_vector(31 downto 0);
  signal cst_88_int_d_wire : bit_vector(31 downto 0);
  signal cst_89_uint_d_wire : bit_vector(31 downto 0);
  signal cst_8_int_d_wire : bit_vector(31 downto 0);
  signal cst_90_int_d_wire : bit_vector(31 downto 0);
  signal cst_91_uint_d_wire : bit_vector(31 downto 0);
  signal cst_92_uint_d_wire : bit_vector(31 downto 0);
  signal cst_9_uint_d_wire : bit_vector(31 downto 0);
  signal indvar118_d_ph_d_ph_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar121_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar123_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar126_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar129_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar132_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar134_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar138_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar143_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar146_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar148_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar151_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar153_mux_1_d_wire : bit_vector(31 downto 0);
  signal indvar_mux_1_d_wire : bit_vector(31 downto 0);
  signal j_d_3_d_in_d_ph_mux_1_d_wire : bit_vector(31 downto 0);
  signal j_d_3_d_in_mux_1_d_wire : bit_vector(31 downto 0);
  signal j_d_9_d_2_d_be_mux_1_d_wire : bit_vector(31 downto 0);
  signal j_d_9_d_2_d_be_mux_2_d_wire : bit_vector(31 downto 0);
  signal j_d_9_d_2_mux_1_d_wire : bit_vector(31 downto 0);
  signal k_d_1_d_in_d_ph_mux_1_d_wire : bit_vector(31 downto 0);
  signal k_d_2_d_3_mux_1_d_wire : bit_vector(31 downto 0);
  signal k_d_3_d_0_mux_1_d_wire : bit_vector(31 downto 0);
  signal k_d_4_d_3_mux_1_d_wire : bit_vector(31 downto 0);
  signal k_d_5_d_0_mux_1_d_wire : bit_vector(31 downto 0);
  signal load_A_d_wire : bit_vector(31 downto 0);
  signal load_ccoeff_d_wire : bit_vector(31 downto 0);
  signal load_l_array_d_wire : bit_vector(31 downto 0);
  signal load_noofelem_d_wire : bit_vector(31 downto 0);
  signal load_rcoeff_d_wire : bit_vector(31 downto 0);
  signal load_start_call_divide_0_return_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_103_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_108_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_123_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_128_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_133_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_159_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_180_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_193_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_211_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_21_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_230_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_26_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_31_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_48_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_53_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_66_d_wire : bit_vector(31 downto 0);
  signal load_tmp_d_75_d_wire : bit_vector(31 downto 0);
  signal load_u_array_d_wire : bit_vector(31 downto 0);
  signal location_start_B_d_wire : bit_vector(31 downto 0);
  signal location_start_L_d_wire : bit_vector(31 downto 0);
  signal location_start_U_d_wire : bit_vector(31 downto 0);
  signal location_start_call_divide_0_actual_0_d_wire : bit_vector(31 downto 0);
  signal location_start_call_divide_0_actual_1_d_wire : bit_vector(31 downto 0);
  signal location_start_call_divide_0_return_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_0_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_1_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_2_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_3_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_4_d_wire : bit_vector(31 downto 0);
  signal location_start_formal_5_d_wire : bit_vector(31 downto 0);
  signal maxcoeff_d_2_d_2_mux_1_d_wire : bit_vector(31 downto 0);
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_wire : bit_vector(31 downto 0);
  signal maxcoeff_d_2_d_ph_mux_1_d_wire : bit_vector(31 downto 0);
  signal maxcoeff_d_2_mux_1_d_wire : bit_vector(31 downto 0);
  signal oper_exitcond120_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond128_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond131_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond142_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond145_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond150_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond158_bool_d_wire : bit_vector(0 downto 0);
  signal oper_exitcond_bool_d_wire : bit_vector(0 downto 0);
  signal oper_inc_d_11_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_12_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_14_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_15_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_2_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_5_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_960_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_976_int_d_wire : bit_vector(31 downto 0);
  signal oper_inc_d_9_int_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next119_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next122_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next124_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next127_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next130_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next133_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next139_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next144_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next147_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next149_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next152_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next157_uint_d_wire : bit_vector(31 downto 0);
  signal oper_indvar_d_next_uint_d_wire : bit_vector(31 downto 0);
  signal oper_j_d_321_int_d_wire : bit_vector(31 downto 0);
  signal oper_j_d_3_int_d_wire : bit_vector(31 downto 0);
  signal oper_j_d_746_int_d_wire : bit_vector(31 downto 0);
  signal oper_j_d_7_int_d_wire : bit_vector(31 downto 0);
  signal oper_k_d_1_d_in_int_d_wire : bit_vector(31 downto 0);
  signal oper_k_d_1_int_d_wire : bit_vector(31 downto 0);
  signal oper_k_d_2_d_2_int_d_wire : bit_vector(31 downto 0);
  signal oper_k_d_4_d_2_int_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_107_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_11348_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_113_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_11_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_125_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_132_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_134_float_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_135_float_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_136_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_137_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_14574_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_14578_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_14580_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_149_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_155_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_158_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_1614_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_166_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_16_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_175_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_179_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_188_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_192_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_20299_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_202_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_210_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_221111_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_221_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_229_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_27_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_4223_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_42_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_52_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_54_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_74_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_92_bool_d_wire : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_id_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_wire : bit_vector(31 downto 0);
  signal oper_tmp_d_uint_d_wire : bit_vector(31 downto 0);
  signal tc_i_d_1_d_0_d_wire : bit_vector(31 downto 0);
  signal tc_i_d_2_d_0_d_ph_d_wire : bit_vector(31 downto 0);
  signal tc_i_d_3_d_0_d_ph_d_wire : bit_vector(31 downto 0);
  signal tc_i_d_4_d_0_d_wire : bit_vector(31 downto 0);
  signal tc_i_d_5_d_0_d_wire : bit_vector(31 downto 0);
  signal tc_indvar138_d_wire : bit_vector(31 downto 0);
  signal tc_indvar151_d_wire : bit_vector(31 downto 0);
  signal tc_j_d_11_d_2_d_wire : bit_vector(31 downto 0);
  signal tc_j_d_13_d_2_d_wire : bit_vector(31 downto 0);
  signal tc_j_d_3_d_2_d_wire : bit_vector(31 downto 0);
  signal tc_j_d_3_d_in_d_wire : bit_vector(31 downto 0);
  signal tc_j_d_7_d_1_d_wire : bit_vector(31 downto 0);
  signal tc_p_d_0_d_0_d_ph_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_wire : bit_vector(31 downto 0);
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_wire : bit_vector(31 downto 0);

begin

  cbr_10_oper_tmp_d_42_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_42_bool_d_wire -- in
    , req0 => ip(58)
    , ack0 => op(55)
    , ack1 => op(54)
    , reset => reset
    , clk => clk);

  cbr_11_oper_tmp_d_54_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_54_bool_d_wire -- in
    , req0 => ip(73)
    , ack0 => op(69)
    , ack1 => op(68)
    , reset => reset
    , clk => clk);

  cbr_12_oper_tmp_d_4223_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_4223_bool_d_wire -- in
    , req0 => ip(77)
    , ack0 => op(74)
    , ack1 => op(73)
    , reset => reset
    , clk => clk);

  cbr_13_oper_exitcond128_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond128_bool_d_wire -- in
    , req0 => ip(95)
    , ack0 => op(91)
    , ack1 => op(90)
    , reset => reset
    , clk => clk);

  cbr_14_oper_exitcond131_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond131_bool_d_wire -- in
    , req0 => ip(99)
    , ack0 => op(96)
    , ack1 => op(95)
    , reset => reset
    , clk => clk);

  cbr_15_oper_tmp_d_92_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_92_bool_d_wire -- in
    , req0 => ip(117)
    , ack0 => op(112)
    , ack1 => op(111)
    , reset => reset
    , clk => clk);

  cbr_16_oper_tmp_d_11348_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_11348_bool_d_wire -- in
    , req0 => ip(128)
    , ack0 => op(124)
    , ack1 => op(123)
    , reset => reset
    , clk => clk);

  cbr_17_oper_tmp_d_113_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_113_bool_d_wire -- in
    , req0 => ip(150)
    , ack0 => op(146)
    , ack1 => op(145)
    , reset => reset
    , clk => clk);

  cbr_18_oper_exitcond142_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond142_bool_d_wire -- in
    , req0 => ip(152)
    , ack0 => op(149)
    , ack1 => op(148)
    , reset => reset
    , clk => clk);

  cbr_19_oper_tmp_d_149_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_149_bool_d_wire -- in
    , req0 => ip(159)
    , ack0 => op(155)
    , ack1 => op(154)
    , reset => reset
    , clk => clk);

  cbr_20_oper_tmp_d_14574_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_14574_bool_d_wire -- in
    , req0 => ip(177)
    , ack0 => op(174)
    , ack1 => op(173)
    , reset => reset
    , clk => clk);

  cbr_21_oper_tmp_d_166_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_166_bool_d_wire -- in
    , req0 => ip(187)
    , ack0 => op(183)
    , ack1 => op(182)
    , reset => reset
    , clk => clk);

  cbr_22_oper_tmp_d_14578_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_14578_bool_d_wire -- in
    , req0 => ip(201)
    , ack0 => op(198)
    , ack1 => op(197)
    , reset => reset
    , clk => clk);

  cbr_23_oper_tmp_d_14580_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_14580_bool_d_wire -- in
    , req0 => ip(215)
    , ack0 => op(213)
    , ack1 => op(212)
    , reset => reset
    , clk => clk);

  cbr_24_oper_exitcond145_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond145_bool_d_wire -- in
    , req0 => ip(218)
    , ack0 => op(217)
    , ack1 => op(216)
    , reset => reset
    , clk => clk);

  cbr_25_oper_tmp_d_202_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_202_bool_d_wire -- in
    , req0 => ip(225)
    , ack0 => op(223)
    , ack1 => op(222)
    , reset => reset
    , clk => clk);

  cbr_26_oper_tmp_d_20299_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_20299_bool_d_wire -- in
    , req0 => ip(240)
    , ack0 => op(238)
    , ack1 => op(237)
    , reset => reset
    , clk => clk);

  cbr_27_oper_exitcond150_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond150_bool_d_wire -- in
    , req0 => ip(246)
    , ack0 => op(244)
    , ack1 => op(243)
    , reset => reset
    , clk => clk);

  cbr_28_oper_tmp_d_221_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_221_bool_d_wire -- in
    , req0 => ip(253)
    , ack0 => op(250)
    , ack1 => op(249)
    , reset => reset
    , clk => clk);

  cbr_29_oper_tmp_d_221111_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_221111_bool_d_wire -- in
    , req0 => ip(270)
    , ack0 => op(267)
    , ack1 => op(266)
    , reset => reset
    , clk => clk);

  cbr_30_oper_exitcond158_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond158_bool_d_wire -- in
    , req0 => ip(276)
    , ack0 => op(273)
    , ack1 => op(272)
    , reset => reset
    , clk => clk);

  cbr_6_oper_exitcond_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond_bool_d_wire -- in
    , req0 => ip(17)
    , ack0 => op(16)
    , ack1 => op(15)
    , reset => reset
    , clk => clk);

  cbr_7_oper_exitcond120_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_exitcond120_bool_d_wire -- in
    , req0 => ip(20)
    , ack0 => op(20)
    , ack1 => op(19)
    , reset => reset
    , clk => clk);

  cbr_8_oper_tmp_d_16_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_16_bool_d_wire -- in
    , req0 => ip(22)
    , ack0 => op(23)
    , ack1 => op(22)
    , reset => reset
    , clk => clk);

  cbr_9_oper_tmp_d_1614_bool : libdec
  generic map(
     ip_wd => 1)
  port map(
    ip => oper_tmp_d_1614_bool_d_wire -- in
    , req0 => ip(41)
    , ack0 => op(42)
    , ack1 => op(41)
    , reset => reset
    , clk => clk);

  indvar118_d_ph_d_ph_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => cst_0_uint_d_wire -- in
    , ip1 => oper_indvar_d_next119_uint_d_wire -- in
    , op => indvar118_d_ph_d_ph_mux_1_d_wire -- out
    , req0 => ip(7)
    , req1 => ip(8)
    , ack0 => op(7)
    , reset => reset
    , clk => clk);

  indvar121_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next122_uint_d_wire -- in
    , ip1 => cst_9_uint_d_wire -- in
    , op => indvar121_mux_1_d_wire -- out
    , req0 => ip(23)
    , req1 => ip(24)
    , ack0 => op(24)
    , reset => reset
    , clk => clk);

  indvar123_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => cst_20_uint_d_wire -- in
    , ip1 => oper_indvar_d_next124_uint_d_wire -- in
    , op => indvar123_mux_1_d_wire -- out
    , req0 => ip(62)
    , req1 => ip(63)
    , ack0 => op(59)
    , reset => reset
    , clk => clk);

  indvar126_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next127_uint_d_wire -- in
    , ip1 => cst_25_uint_d_wire -- in
    , op => indvar126_mux_1_d_wire -- out
    , req0 => ip(80)
    , req1 => ip(81)
    , ack0 => op(76)
    , reset => reset
    , clk => clk);

  indvar129_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next130_uint_d_wire -- in
    , ip1 => cst_13_uint_d_wire -- in
    , op => indvar129_mux_1_d_wire -- out
    , req0 => ip(42)
    , req1 => ip(43)
    , ack0 => op(43)
    , reset => reset
    , clk => clk);

  indvar132_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next133_uint_d_wire -- in
    , ip1 => cst_44_uint_d_wire -- in
    , op => indvar132_mux_1_d_wire -- out
    , req0 => ip(130)
    , req1 => ip(131)
    , ack0 => op(126)
    , reset => reset
    , clk => clk);

  indvar134_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_136_uint_d_wire -- in
    , ip1 => cst_33_uint_d_wire -- in
    , op => indvar134_mux_1_d_wire -- out
    , req0 => ip(100)
    , req1 => ip(101)
    , ack0 => op(97)
    , reset => reset
    , clk => clk);

  indvar138_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => cst_39_uint_d_wire -- in
    , ip1 => oper_indvar_d_next139_uint_d_wire -- in
    , op => indvar138_mux_1_d_wire -- out
    , req0 => ip(111)
    , req1 => ip(112)
    , ack0 => op(106)
    , reset => reset
    , clk => clk);

  indvar143_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next144_uint_d_wire -- in
    , ip1 => cst_51_uint_d_wire -- in
    , op => indvar143_mux_1_d_wire -- out
    , req0 => ip(153)
    , req1 => ip(154)
    , ack0 => op(150)
    , reset => reset
    , clk => clk);

  indvar146_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next147_uint_d_wire -- in
    , ip1 => cst_75_uint_d_wire -- in
    , op => indvar146_mux_1_d_wire -- out
    , req0 => ip(226)
    , req1 => ip(227)
    , ack0 => op(224)
    , reset => reset
    , clk => clk);

  indvar148_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next149_uint_d_wire -- in
    , ip1 => cst_72_uint_d_wire -- in
    , op => indvar148_mux_1_d_wire -- out
    , req0 => ip(219)
    , req1 => ip(220)
    , ack0 => op(218)
    , reset => reset
    , clk => clk);

  indvar151_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next152_uint_d_wire -- in
    , ip1 => cst_85_uint_d_wire -- in
    , op => indvar151_mux_1_d_wire -- out
    , req0 => ip(254)
    , req1 => ip(255)
    , ack0 => op(251)
    , reset => reset
    , clk => clk);

  indvar153_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next157_uint_d_wire -- in
    , ip1 => cst_82_uint_d_wire -- in
    , op => indvar153_mux_1_d_wire -- out
    , req0 => ip(247)
    , req1 => ip(248)
    , ack0 => op(245)
    , reset => reset
    , clk => clk);

  indvar_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_indvar_d_next_uint_d_wire -- in
    , ip1 => cst_1_uint_d_wire -- in
    , op => indvar_mux_1_d_wire -- out
    , req0 => ip(9)
    , req1 => ip(10)
    , ack0 => op(8)
    , reset => reset
    , clk => clk);

  j_d_3_d_in_d_ph_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_inc_d_5_int_d_wire -- in
    , ip1 => cst_14_int_d_wire -- in
    , op => j_d_3_d_in_d_ph_mux_1_d_wire -- out
    , req0 => ip(44)
    , req1 => ip(45)
    , ack0 => op(44)
    , reset => reset
    , clk => clk);

  j_d_3_d_in_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_3_d_in_d_ph_mux_1_d_wire -- in
    , ip1 => tc_j_d_3_d_2_d_wire -- in
    , op => j_d_3_d_in_mux_1_d_wire -- out
    , req0 => ip(52)
    , req1 => ip(53)
    , ack0 => op(50)
    , reset => reset
    , clk => clk);

  j_d_9_d_2_d_be_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_inc_d_960_int_d_wire -- in
    , ip1 => oper_inc_d_976_int_d_wire -- in
    , op => j_d_9_d_2_d_be_mux_1_d_wire -- out
    , req0 => ip(180)
    , req1 => ip(181)
    , ack0 => op(176)
    , reset => reset
    , clk => clk);

  j_d_9_d_2_d_be_mux_2 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_9_d_2_d_be_mux_1_d_wire -- in
    , ip1 => oper_inc_d_9_int_d_wire -- in
    , op => j_d_9_d_2_d_be_mux_2_d_wire -- out
    , req0 => ip(178)
    , req1 => ip(179)
    , ack0 => op(175)
    , reset => reset
    , clk => clk);

  j_d_9_d_2_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => cst_52_int_d_wire -- in
    , ip1 => j_d_9_d_2_d_be_mux_2_d_wire -- in
    , op => j_d_9_d_2_mux_1_d_wire -- out
    , req0 => ip(156)
    , req1 => ip(157)
    , ack0 => op(152)
    , reset => reset
    , clk => clk);

  k_d_1_d_in_d_ph_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_j_d_746_int_d_wire -- in
    , ip1 => cst_34_int_d_wire -- in
    , op => k_d_1_d_in_d_ph_mux_1_d_wire -- out
    , req0 => ip(102)
    , req1 => ip(103)
    , ack0 => op(98)
    , reset => reset
    , clk => clk);

  k_d_2_d_3_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => k_d_3_d_0_mux_1_d_wire -- in
    , ip1 => oper_inc_d_11_int_d_wire -- in
    , op => k_d_2_d_3_mux_1_d_wire -- out
    , req0 => ip(242)
    , req1 => ip(243)
    , ack0 => op(240)
    , reset => reset
    , clk => clk);

  k_d_3_d_0_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => k_d_2_d_3_mux_1_d_wire -- in
    , ip1 => cst_73_int_d_wire -- in
    , op => k_d_3_d_0_mux_1_d_wire -- out
    , req0 => ip(221)
    , req1 => ip(222)
    , ack0 => op(219)
    , reset => reset
    , clk => clk);

  k_d_4_d_3_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => k_d_5_d_0_mux_1_d_wire -- in
    , ip1 => oper_inc_d_14_int_d_wire -- in
    , op => k_d_4_d_3_mux_1_d_wire -- out
    , req0 => ip(272)
    , req1 => ip(273)
    , ack0 => op(269)
    , reset => reset
    , clk => clk);

  k_d_5_d_0_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => k_d_4_d_3_mux_1_d_wire -- in
    , ip1 => cst_83_int_d_wire -- in
    , op => k_d_5_d_0_mux_1_d_wire -- out
    , req0 => ip(249)
    , req1 => ip(250)
    , ack0 => op(246)
    , reset => reset
    , clk => clk);

  load_A : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_1_d_wire -- in
    , dp => load_A_d_wire -- out
    , req0 => ip(2)
    , ack0 => op(2)
    , mreq => load_reqs(0)
    , mack => load_acks(0)
    , maddr => load_addr(0)
    , mdata => load_data(0)
    , reset => reset
    , clk => clk);

  load_ccoeff : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_3_d_wire -- in
    , dp => load_ccoeff_d_wire -- out
    , req0 => ip(4)
    , ack0 => op(4)
    , mreq => load_reqs(1)
    , mack => load_acks(1)
    , maddr => load_addr(1)
    , mdata => load_data(1)
    , reset => reset
    , clk => clk);

  load_l_array : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_4_d_wire -- in
    , dp => load_l_array_d_wire -- out
    , req0 => ip(5)
    , ack0 => op(5)
    , mreq => load_reqs(2)
    , mack => load_acks(2)
    , maddr => load_addr(2)
    , mdata => load_data(2)
    , reset => reset
    , clk => clk);

  load_noofelem : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_0_d_wire -- in
    , dp => load_noofelem_d_wire -- out
    , req0 => ip(1)
    , ack0 => op(1)
    , mreq => load_reqs(3)
    , mack => load_acks(3)
    , maddr => load_addr(3)
    , mdata => load_data(3)
    , reset => reset
    , clk => clk);

  load_rcoeff : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_2_d_wire -- in
    , dp => load_rcoeff_d_wire -- out
    , req0 => ip(3)
    , ack0 => op(3)
    , mreq => load_reqs(4)
    , mack => load_acks(4)
    , maddr => load_addr(4)
    , mdata => load_data(4)
    , reset => reset
    , clk => clk);

  load_start_call_divide_0_return : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_call_divide_0_return_d_wire -- in
    , dp => load_start_call_divide_0_return_d_wire -- out
    , req0 => ip(126)
    , ack0 => op(121)
    , mreq => load_reqs(5)
    , mack => load_acks(5)
    , maddr => load_addr(5)
    , mdata => load_data(5)
    , reset => reset
    , clk => clk);

  load_tmp_d_103 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_97_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_103_d_wire -- out
    , req0 => ip(122)
    , ack0 => op(117)
    , mreq => load_reqs(6)
    , mack => load_acks(6)
    , maddr => load_addr(6)
    , mdata => load_data(6)
    , reset => reset
    , clk => clk);

  load_tmp_d_108 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_107_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_108_d_wire -- out
    , req0 => ip(123)
    , ack0 => op(118)
    , mreq => load_reqs(7)
    , mack => load_acks(7)
    , maddr => load_addr(7)
    , mdata => load_data(7)
    , reset => reset
    , clk => clk);

  load_tmp_d_123 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_118_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_123_d_wire -- out
    , req0 => ip(138)
    , ack0 => op(133)
    , mreq => load_reqs(8)
    , mack => load_acks(8)
    , maddr => load_addr(8)
    , mdata => load_data(8)
    , reset => reset
    , clk => clk);

  load_tmp_d_128 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_97_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_128_d_wire -- out
    , req0 => ip(139)
    , ack0 => op(134)
    , mreq => load_reqs(9)
    , mack => load_acks(9)
    , maddr => load_addr(9)
    , mdata => load_data(9)
    , reset => reset
    , clk => clk);

  load_tmp_d_133 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_132_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_133_d_wire -- out
    , req0 => ip(143)
    , ack0 => op(138)
    , mreq => load_reqs(10)
    , mack => load_acks(10)
    , maddr => load_addr(10)
    , mdata => load_data(10)
    , reset => reset
    , clk => clk);

  load_tmp_d_159 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_158_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_159_d_wire -- out
    , req0 => ip(168)
    , ack0 => op(164)
    , mreq => load_reqs(11)
    , mack => load_acks(11)
    , maddr => load_addr(11)
    , mdata => load_data(11)
    , reset => reset
    , clk => clk);

  load_tmp_d_180 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_179_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_180_d_wire -- out
    , req0 => ip(197)
    , ack0 => op(193)
    , mreq => load_reqs(12)
    , mack => load_acks(12)
    , maddr => load_addr(12)
    , mdata => load_data(12)
    , reset => reset
    , clk => clk);

  load_tmp_d_193 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_192_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_193_d_wire -- out
    , req0 => ip(211)
    , ack0 => op(208)
    , mreq => load_reqs(13)
    , mack => load_acks(13)
    , maddr => load_addr(13)
    , mdata => load_data(13)
    , reset => reset
    , clk => clk);

  load_tmp_d_21 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_20_d_lvl_d_0_uint_d_wire -- in
    , dp => load_tmp_d_21_d_wire -- out
    , req0 => ip(27)
    , ack0 => op(27)
    , mreq => load_reqs(14)
    , mack => load_acks(14)
    , maddr => load_addr(14)
    , mdata => load_data(14)
    , reset => reset
    , clk => clk);

  load_tmp_d_211 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_210_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_211_d_wire -- out
    , req0 => ip(235)
    , ack0 => op(232)
    , mreq => load_reqs(15)
    , mack => load_acks(15)
    , maddr => load_addr(15)
    , mdata => load_data(15)
    , reset => reset
    , clk => clk);

  load_tmp_d_230 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_229_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_230_d_wire -- out
    , req0 => ip(265)
    , ack0 => op(261)
    , mreq => load_reqs(16)
    , mack => load_acks(16)
    , maddr => load_addr(16)
    , mdata => load_data(16)
    , reset => reset
    , clk => clk);

  load_tmp_d_26 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_25_d_lvl_d_0_uint_d_wire -- in
    , dp => load_tmp_d_26_d_wire -- out
    , req0 => ip(29)
    , ack0 => op(29)
    , mreq => load_reqs(17)
    , mack => load_acks(17)
    , maddr => load_addr(17)
    , mdata => load_data(17)
    , reset => reset
    , clk => clk);

  load_tmp_d_31 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_30_d_lvl_d_0_uint_d_wire -- in
    , dp => load_tmp_d_31_d_wire -- out
    , req0 => ip(36)
    , ack0 => op(36)
    , mreq => load_reqs(18)
    , mack => load_acks(18)
    , maddr => load_addr(18)
    , mdata => load_data(18)
    , reset => reset
    , clk => clk);

  load_tmp_d_48 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_47_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_48_d_wire -- out
    , req0 => ip(71)
    , ack0 => op(66)
    , mreq => load_reqs(19)
    , mack => load_acks(19)
    , maddr => load_addr(19)
    , mdata => load_data(19)
    , reset => reset
    , clk => clk);

  load_tmp_d_53 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_52_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_53_d_wire -- out
    , req0 => ip(60)
    , ack0 => op(57)
    , mreq => load_reqs(20)
    , mack => load_acks(20)
    , maddr => load_addr(20)
    , mdata => load_data(20)
    , reset => reset
    , clk => clk);

  load_tmp_d_66 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_65_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_66_d_wire -- out
    , req0 => ip(85)
    , ack0 => op(80)
    , mreq => load_reqs(21)
    , mack => load_acks(21)
    , maddr => load_addr(21)
    , mdata => load_data(21)
    , reset => reset
    , clk => clk);

  load_tmp_d_75 : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_74_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_75_d_wire -- out
    , req0 => ip(90)
    , ack0 => op(85)
    , mreq => load_reqs(22)
    , mack => load_acks(22)
    , maddr => load_addr(22)
    , mdata => load_data(22)
    , reset => reset
    , clk => clk);

  load_u_array : liblod
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_formal_5_d_wire -- in
    , dp => load_u_array_d_wire -- out
    , req0 => ip(6)
    , ack0 => op(6)
    , mreq => load_reqs(23)
    , mack => load_acks(23)
    , maddr => load_addr(23)
    , mdata => load_data(23)
    , reset => reset
    , clk => clk);

  maxcoeff_d_2_d_2_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => maxcoeff_d_2_mux_1_d_wire -- in
    , ip1 => tc_j_d_3_d_2_d_wire -- in
    , op => maxcoeff_d_2_d_2_mux_1_d_wire -- out
    , req0 => ip(64)
    , req1 => ip(65)
    , ack0 => op(60)
    , reset => reset
    , clk => clk);

  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => maxcoeff_d_2_mux_1_d_wire -- in
    , ip1 => tc_j_d_3_d_2_d_wire -- in
    , op => maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_wire -- out
    , req0 => ip(78)
    , req1 => ip(79)
    , ack0 => op(75)
    , reset => reset
    , clk => clk);

  maxcoeff_d_2_d_ph_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_inc_d_5_int_d_wire -- in
    , ip1 => cst_15_int_d_wire -- in
    , op => maxcoeff_d_2_d_ph_mux_1_d_wire -- out
    , req0 => ip(46)
    , req1 => ip(47)
    , ack0 => op(45)
    , reset => reset
    , clk => clk);

  maxcoeff_d_2_mux_1 : libmux
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => maxcoeff_d_2_d_ph_mux_1_d_wire -- in
    , ip1 => maxcoeff_d_2_d_2_mux_1_d_wire -- in
    , op => maxcoeff_d_2_mux_1_d_wire -- out
    , req0 => ip(54)
    , req1 => ip(55)
    , ack0 => op(51)
    , reset => reset
    , clk => clk);

  oper_exitcond120_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next119_uint_d_wire -- in
    , ip1 => cst_7_uint_d_wire -- in
    , op => oper_exitcond120_bool_d_wire -- out
    , req0 => ip(19)
    , ack0 => op(18)
    , reset => reset
    , clk => clk);

  oper_exitcond128_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next127_uint_d_wire -- in
    , ip1 => cst_29_uint_d_wire -- in
    , op => oper_exitcond128_bool_d_wire -- out
    , req0 => ip(94)
    , ack0 => op(89)
    , reset => reset
    , clk => clk);

  oper_exitcond131_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next130_uint_d_wire -- in
    , ip1 => cst_32_uint_d_wire -- in
    , op => oper_exitcond131_bool_d_wire -- out
    , req0 => ip(98)
    , ack0 => op(94)
    , reset => reset
    , clk => clk);

  oper_exitcond142_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_tmp_d_136_uint_d_wire -- in
    , ip1 => cst_50_uint_d_wire -- in
    , op => oper_exitcond142_bool_d_wire -- out
    , req0 => ip(151)
    , ack0 => op(147)
    , reset => reset
    , clk => clk);

  oper_exitcond145_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next144_uint_d_wire -- in
    , ip1 => cst_71_uint_d_wire -- in
    , op => oper_exitcond145_bool_d_wire -- out
    , req0 => ip(217)
    , ack0 => op(215)
    , reset => reset
    , clk => clk);

  oper_exitcond150_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next149_uint_d_wire -- in
    , ip1 => cst_81_uint_d_wire -- in
    , op => oper_exitcond150_bool_d_wire -- out
    , req0 => ip(245)
    , ack0 => op(242)
    , reset => reset
    , clk => clk);

  oper_exitcond158_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next157_uint_d_wire -- in
    , ip1 => cst_92_uint_d_wire -- in
    , op => oper_exitcond158_bool_d_wire -- out
    , req0 => ip(275)
    , ack0 => op(271)
    , reset => reset
    , clk => clk);

  oper_exitcond_bool : libeq_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_indvar_d_next_uint_d_wire -- in
    , ip1 => cst_5_uint_d_wire -- in
    , op => oper_exitcond_bool_d_wire -- out
    , req0 => ip(16)
    , ack0 => op(14)
    , reset => reset
    , clk => clk);

  oper_inc_d_11_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_k_d_2_d_2_int_d_wire -- in
    , ip1 => cst_79_int_d_wire -- in
    , op => oper_inc_d_11_int_d_wire -- out
    , req0 => ip(241)
    , ack0 => op(239)
    , reset => reset
    , clk => clk);

  oper_inc_d_12_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_11_d_2_d_wire -- in
    , ip1 => cst_77_int_d_wire -- in
    , op => oper_inc_d_12_int_d_wire -- out
    , req0 => ip(237)
    , ack0 => op(234)
    , reset => reset
    , clk => clk);

  oper_inc_d_14_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_k_d_4_d_2_int_d_wire -- in
    , ip1 => cst_90_int_d_wire -- in
    , op => oper_inc_d_14_int_d_wire -- out
    , req0 => ip(271)
    , ack0 => op(268)
    , reset => reset
    , clk => clk);

  oper_inc_d_15_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_13_d_2_d_wire -- in
    , ip1 => cst_87_int_d_wire -- in
    , op => oper_inc_d_15_int_d_wire -- out
    , req0 => ip(267)
    , ack0 => op(263)
    , reset => reset
    , clk => clk);

  oper_inc_d_2_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_i_d_1_d_0_d_wire -- in
    , ip1 => cst_11_int_d_wire -- in
    , op => oper_inc_d_2_int_d_wire -- out
    , req0 => ip(38)
    , ack0 => op(38)
    , reset => reset
    , clk => clk);

  oper_inc_d_5_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_i_d_2_d_0_d_ph_d_wire -- in
    , ip1 => cst_30_int_d_wire -- in
    , op => oper_inc_d_5_int_d_wire -- out
    , req0 => ip(96)
    , ack0 => op(92)
    , reset => reset
    , clk => clk);

  oper_inc_d_960_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_9_d_2_mux_1_d_wire -- in
    , ip1 => cst_57_int_d_wire -- in
    , op => oper_inc_d_960_int_d_wire -- out
    , req0 => ip(175)
    , ack0 => op(171)
    , reset => reset
    , clk => clk);

  oper_inc_d_976_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_9_d_2_mux_1_d_wire -- in
    , ip1 => cst_63_int_d_wire -- in
    , op => oper_inc_d_976_int_d_wire -- out
    , req0 => ip(199)
    , ack0 => op(195)
    , reset => reset
    , clk => clk);

  oper_inc_d_9_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_9_d_2_mux_1_d_wire -- in
    , ip1 => cst_68_int_d_wire -- in
    , op => oper_inc_d_9_int_d_wire -- out
    , req0 => ip(213)
    , ack0 => op(210)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next119_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar118_d_ph_d_ph_mux_1_d_wire -- in
    , ip1 => cst_6_uint_d_wire -- in
    , op => oper_indvar_d_next119_uint_d_wire -- out
    , req0 => ip(18)
    , ack0 => op(17)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next122_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar121_mux_1_d_wire -- in
    , ip1 => cst_12_uint_d_wire -- in
    , op => oper_indvar_d_next122_uint_d_wire -- out
    , req0 => ip(40)
    , ack0 => op(40)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next124_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar123_mux_1_d_wire -- in
    , ip1 => cst_24_uint_d_wire -- in
    , op => oper_indvar_d_next124_uint_d_wire -- out
    , req0 => ip(76)
    , ack0 => op(72)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next127_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar126_mux_1_d_wire -- in
    , ip1 => cst_28_uint_d_wire -- in
    , op => oper_indvar_d_next127_uint_d_wire -- out
    , req0 => ip(93)
    , ack0 => op(88)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next130_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar129_mux_1_d_wire -- in
    , ip1 => cst_31_uint_d_wire -- in
    , op => oper_indvar_d_next130_uint_d_wire -- out
    , req0 => ip(97)
    , ack0 => op(93)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next133_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar132_mux_1_d_wire -- in
    , ip1 => cst_49_uint_d_wire -- in
    , op => oper_indvar_d_next133_uint_d_wire -- out
    , req0 => ip(149)
    , ack0 => op(144)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next139_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar138_mux_1_d_wire -- in
    , ip1 => cst_43_uint_d_wire -- in
    , op => oper_indvar_d_next139_uint_d_wire -- out
    , req0 => ip(129)
    , ack0 => op(125)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next144_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_70_uint_d_wire -- in
    , op => oper_indvar_d_next144_uint_d_wire -- out
    , req0 => ip(216)
    , ack0 => op(214)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next147_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar146_mux_1_d_wire -- in
    , ip1 => cst_78_uint_d_wire -- in
    , op => oper_indvar_d_next147_uint_d_wire -- out
    , req0 => ip(239)
    , ack0 => op(236)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next149_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar148_mux_1_d_wire -- in
    , ip1 => cst_80_uint_d_wire -- in
    , op => oper_indvar_d_next149_uint_d_wire -- out
    , req0 => ip(244)
    , ack0 => op(241)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next152_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar151_mux_1_d_wire -- in
    , ip1 => cst_89_uint_d_wire -- in
    , op => oper_indvar_d_next152_uint_d_wire -- out
    , req0 => ip(269)
    , ack0 => op(265)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next157_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar153_mux_1_d_wire -- in
    , ip1 => cst_91_uint_d_wire -- in
    , op => oper_indvar_d_next157_uint_d_wire -- out
    , req0 => ip(274)
    , ack0 => op(270)
    , reset => reset
    , clk => clk);

  oper_indvar_d_next_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar_mux_1_d_wire -- in
    , ip1 => cst_4_uint_d_wire -- in
    , op => oper_indvar_d_next_uint_d_wire -- out
    , req0 => ip(15)
    , ack0 => op(13)
    , reset => reset
    , clk => clk);

  oper_j_d_321_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_3_d_2_d_wire -- in
    , ip1 => cst_22_int_d_wire -- in
    , op => oper_j_d_321_int_d_wire -- out
    , req0 => ip(74)
    , ack0 => op(70)
    , reset => reset
    , clk => clk);

  oper_j_d_3_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => j_d_3_d_in_mux_1_d_wire -- in
    , ip1 => cst_17_int_d_wire -- in
    , op => oper_j_d_3_int_d_wire -- out
    , req0 => ip(56)
    , ack0 => op(52)
    , reset => reset
    , clk => clk);

  oper_j_d_746_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_p_d_0_d_0_d_ph_d_wire -- in
    , ip1 => cst_36_int_d_wire -- in
    , op => oper_j_d_746_int_d_wire -- out
    , req0 => ip(108)
    , ack0 => op(103)
    , reset => reset
    , clk => clk);

  oper_j_d_7_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_7_d_1_d_wire -- in
    , ip1 => cst_47_int_d_wire -- in
    , op => oper_j_d_7_int_d_wire -- out
    , req0 => ip(147)
    , ack0 => op(142)
    , reset => reset
    , clk => clk);

  oper_k_d_1_d_in_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_indvar138_d_wire -- in
    , ip1 => k_d_1_d_in_d_ph_mux_1_d_wire -- in
    , op => oper_k_d_1_d_in_int_d_wire -- out
    , req0 => ip(114)
    , ack0 => op(108)
    , reset => reset
    , clk => clk);

  oper_k_d_1_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_k_d_1_d_in_int_d_wire -- in
    , ip1 => cst_40_int_d_wire -- in
    , op => oper_k_d_1_int_d_wire -- out
    , req0 => ip(115)
    , ack0 => op(109)
    , reset => reset
    , clk => clk);

  oper_k_d_2_d_2_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_11_d_2_d_wire -- in
    , ip1 => k_d_3_d_0_mux_1_d_wire -- in
    , op => oper_k_d_2_d_2_int_d_wire -- out
    , req0 => ip(229)
    , ack0 => op(226)
    , reset => reset
    , clk => clk);

  oper_k_d_4_d_2_int : libadd_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_indvar151_d_wire -- in
    , ip1 => k_d_5_d_0_mux_1_d_wire -- in
    , op => oper_k_d_4_d_2_int_d_wire -- out
    , req0 => ip(259)
    , ack0 => op(255)
    , reset => reset
    , clk => clk);

  oper_tmp_d_107_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar134_mux_1_d_wire -- in
    , ip1 => cst_35_uint_d_wire -- in
    , op => oper_tmp_d_107_d_id_d_1_uint_d_wire -- out
    , req0 => ip(105)
    , ack0 => op(100)
    , reset => reset
    , clk => clk);

  oper_tmp_d_107_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_107_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_107_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(106)
    , ack0 => op(101)
    , reset => reset
    , clk => clk);

  oper_tmp_d_107_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_107_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar134_mux_1_d_wire -- in
    , op => oper_tmp_d_107_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(107)
    , ack0 => op(102)
    , reset => reset
    , clk => clk);

  oper_tmp_d_11348_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_j_d_746_int_d_wire -- in
    , ip1 => cst_37_int_d_wire -- in
    , op => oper_tmp_d_11348_bool_d_wire -- out
    , req0 => ip(109)
    , ack0 => op(104)
    , reset => reset
    , clk => clk);

  oper_tmp_d_113_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_j_d_7_int_d_wire -- in
    , ip1 => cst_48_int_d_wire -- in
    , op => oper_tmp_d_113_bool_d_wire -- out
    , req0 => ip(148)
    , ack0 => op(143)
    , reset => reset
    , clk => clk);

  oper_tmp_d_118_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_tmp_d_118_d_id_d_1_d_cast_d_wire -- in
    , ip1 => cst_45_uint_d_wire -- in
    , op => oper_tmp_d_118_d_id_d_1_uint_d_wire -- out
    , req0 => ip(135)
    , ack0 => op(130)
    , reset => reset
    , clk => clk);

  oper_tmp_d_118_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_118_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_118_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(136)
    , ack0 => op(131)
    , reset => reset
    , clk => clk);

  oper_tmp_d_118_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_118_d_lvl_d_1_uint_d_wire -- in
    , ip1 => oper_tmp_d_137_uint_d_wire -- in
    , op => oper_tmp_d_118_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(137)
    , ack0 => op(132)
    , reset => reset
    , clk => clk);

  oper_tmp_d_11_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar118_d_ph_d_ph_mux_1_d_wire -- in
    , ip1 => cst_2_uint_d_wire -- in
    , op => oper_tmp_d_11_d_id_d_1_uint_d_wire -- out
    , req0 => ip(11)
    , ack0 => op(9)
    , reset => reset
    , clk => clk);

  oper_tmp_d_11_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_11_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_11_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(12)
    , ack0 => op(10)
    , reset => reset
    , clk => clk);

  oper_tmp_d_11_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_11_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar_mux_1_d_wire -- in
    , op => oper_tmp_d_11_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(13)
    , ack0 => op(11)
    , reset => reset
    , clk => clk);

  oper_tmp_d_125_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar123_mux_1_d_wire -- in
    , ip1 => oper_tmp_d_uint_d_wire -- in
    , op => oper_tmp_d_125_uint_d_wire -- out
    , req0 => ip(66)
    , ack0 => op(61)
    , reset => reset
    , clk => clk);

  oper_tmp_d_132_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar134_mux_1_d_wire -- in
    , ip1 => cst_46_uint_d_wire -- in
    , op => oper_tmp_d_132_d_id_d_1_uint_d_wire -- out
    , req0 => ip(140)
    , ack0 => op(135)
    , reset => reset
    , clk => clk);

  oper_tmp_d_132_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_132_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_132_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(141)
    , ack0 => op(136)
    , reset => reset
    , clk => clk);

  oper_tmp_d_132_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_132_d_lvl_d_1_uint_d_wire -- in
    , ip1 => oper_tmp_d_137_uint_d_wire -- in
    , op => oper_tmp_d_132_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(142)
    , ack0 => op(137)
    , reset => reset
    , clk => clk);

  oper_tmp_d_134_float : libmul_float
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_tmp_d_128_d_wire -- in
    , ip1 => load_tmp_d_133_d_wire -- in
    , op => oper_tmp_d_134_float_d_wire -- out
    , req0 => ip(144)
    , ack0 => op(139)
    , reset => reset
    , clk => clk);

  oper_tmp_d_135_float : libsub_float
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_tmp_d_123_d_wire -- in
    , ip1 => oper_tmp_d_134_float_d_wire -- in
    , op => oper_tmp_d_135_float_d_wire -- out
    , req0 => ip(145)
    , ack0 => op(140)
    , reset => reset
    , clk => clk);

  oper_tmp_d_136_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar134_mux_1_d_wire -- in
    , ip1 => cst_38_uint_d_wire -- in
    , op => oper_tmp_d_136_uint_d_wire -- out
    , req0 => ip(110)
    , ack0 => op(105)
    , reset => reset
    , clk => clk);

  oper_tmp_d_137_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar132_mux_1_d_wire -- in
    , ip1 => oper_tmp_d_136_uint_d_wire -- in
    , op => oper_tmp_d_137_uint_d_wire -- out
    , req0 => ip(132)
    , ack0 => op(127)
    , reset => reset
    , clk => clk);

  oper_tmp_d_14574_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_960_int_d_wire -- in
    , ip1 => cst_58_int_d_wire -- in
    , op => oper_tmp_d_14574_bool_d_wire -- out
    , req0 => ip(176)
    , ack0 => op(172)
    , reset => reset
    , clk => clk);

  oper_tmp_d_14578_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_976_int_d_wire -- in
    , ip1 => cst_64_int_d_wire -- in
    , op => oper_tmp_d_14578_bool_d_wire -- out
    , req0 => ip(200)
    , ack0 => op(196)
    , reset => reset
    , clk => clk);

  oper_tmp_d_14580_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_9_int_d_wire -- in
    , ip1 => cst_69_int_d_wire -- in
    , op => oper_tmp_d_14580_bool_d_wire -- out
    , req0 => ip(214)
    , ack0 => op(211)
    , reset => reset
    , clk => clk);

  oper_tmp_d_149_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => j_d_9_d_2_mux_1_d_wire -- in
    , ip1 => tc_i_d_3_d_0_d_ph_d_wire -- in
    , op => oper_tmp_d_149_bool_d_wire -- out
    , req0 => ip(158)
    , ack0 => op(153)
    , reset => reset
    , clk => clk);

  oper_tmp_d_154_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_53_uint_d_wire -- in
    , op => oper_tmp_d_154_d_id_d_1_uint_d_wire -- out
    , req0 => ip(160)
    , ack0 => op(156)
    , reset => reset
    , clk => clk);

  oper_tmp_d_154_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_L_d_wire -- in
    , ip1 => oper_tmp_d_154_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_154_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(161)
    , ack0 => op(157)
    , reset => reset
    , clk => clk);

  oper_tmp_d_154_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_154_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_154_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_154_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(163)
    , ack0 => op(159)
    , reset => reset
    , clk => clk);

  oper_tmp_d_155_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar151_mux_1_d_wire -- in
    , ip1 => indvar153_mux_1_d_wire -- in
    , op => oper_tmp_d_155_uint_d_wire -- out
    , req0 => ip(257)
    , ack0 => op(253)
    , reset => reset
    , clk => clk);

  oper_tmp_d_158_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_54_uint_d_wire -- in
    , op => oper_tmp_d_158_d_id_d_1_uint_d_wire -- out
    , req0 => ip(164)
    , ack0 => op(160)
    , reset => reset
    , clk => clk);

  oper_tmp_d_158_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_158_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_158_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(165)
    , ack0 => op(161)
    , reset => reset
    , clk => clk);

  oper_tmp_d_158_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_158_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_158_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_158_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(167)
    , ack0 => op(163)
    , reset => reset
    , clk => clk);

  oper_tmp_d_1614_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_2_int_d_wire -- in
    , ip1 => load_noofelem_d_wire -- in
    , op => oper_tmp_d_1614_bool_d_wire -- out
    , req0 => ip(39)
    , ack0 => op(39)
    , reset => reset
    , clk => clk);

  oper_tmp_d_163_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_55_uint_d_wire -- in
    , op => oper_tmp_d_163_d_id_d_1_uint_d_wire -- out
    , req0 => ip(170)
    , ack0 => op(166)
    , reset => reset
    , clk => clk);

  oper_tmp_d_163_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_U_d_wire -- in
    , ip1 => oper_tmp_d_163_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_163_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(171)
    , ack0 => op(167)
    , reset => reset
    , clk => clk);

  oper_tmp_d_163_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_163_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_163_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_163_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(173)
    , ack0 => op(169)
    , reset => reset
    , clk => clk);

  oper_tmp_d_166_bool : libeq_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => j_d_9_d_2_mux_1_d_wire -- in
    , ip1 => tc_i_d_3_d_0_d_ph_d_wire -- in
    , op => oper_tmp_d_166_bool_d_wire -- out
    , req0 => ip(182)
    , ack0 => op(177)
    , reset => reset
    , clk => clk);

  oper_tmp_d_16_bool : libgt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => load_noofelem_d_wire -- in
    , ip1 => cst_8_int_d_wire -- in
    , op => oper_tmp_d_16_bool_d_wire -- out
    , req0 => ip(21)
    , ack0 => op(21)
    , reset => reset
    , clk => clk);

  oper_tmp_d_171_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_59_uint_d_wire -- in
    , op => oper_tmp_d_171_d_id_d_1_uint_d_wire -- out
    , req0 => ip(183)
    , ack0 => op(178)
    , reset => reset
    , clk => clk);

  oper_tmp_d_171_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_L_d_wire -- in
    , ip1 => oper_tmp_d_171_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_171_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(184)
    , ack0 => op(179)
    , reset => reset
    , clk => clk);

  oper_tmp_d_171_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_171_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_171_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_171_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(186)
    , ack0 => op(181)
    , reset => reset
    , clk => clk);

  oper_tmp_d_175_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_61_uint_d_wire -- in
    , op => oper_tmp_d_175_d_id_d_1_uint_d_wire -- out
    , req0 => ip(189)
    , ack0 => op(185)
    , reset => reset
    , clk => clk);

  oper_tmp_d_175_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_U_d_wire -- in
    , ip1 => oper_tmp_d_175_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_175_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(190)
    , ack0 => op(186)
    , reset => reset
    , clk => clk);

  oper_tmp_d_175_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_175_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_175_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_175_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(192)
    , ack0 => op(188)
    , reset => reset
    , clk => clk);

  oper_tmp_d_179_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_62_uint_d_wire -- in
    , op => oper_tmp_d_179_d_id_d_1_uint_d_wire -- out
    , req0 => ip(193)
    , ack0 => op(189)
    , reset => reset
    , clk => clk);

  oper_tmp_d_179_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_179_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_179_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(194)
    , ack0 => op(190)
    , reset => reset
    , clk => clk);

  oper_tmp_d_179_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_179_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_179_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_179_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(196)
    , ack0 => op(192)
    , reset => reset
    , clk => clk);

  oper_tmp_d_188_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_66_uint_d_wire -- in
    , op => oper_tmp_d_188_d_id_d_1_uint_d_wire -- out
    , req0 => ip(203)
    , ack0 => op(200)
    , reset => reset
    , clk => clk);

  oper_tmp_d_188_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_U_d_wire -- in
    , ip1 => oper_tmp_d_188_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_188_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(204)
    , ack0 => op(201)
    , reset => reset
    , clk => clk);

  oper_tmp_d_188_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_188_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_188_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_188_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(206)
    , ack0 => op(203)
    , reset => reset
    , clk => clk);

  oper_tmp_d_192_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar143_mux_1_d_wire -- in
    , ip1 => cst_67_uint_d_wire -- in
    , op => oper_tmp_d_192_d_id_d_1_uint_d_wire -- out
    , req0 => ip(207)
    , ack0 => op(204)
    , reset => reset
    , clk => clk);

  oper_tmp_d_192_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_192_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_192_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(208)
    , ack0 => op(205)
    , reset => reset
    , clk => clk);

  oper_tmp_d_192_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_192_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_192_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_192_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(210)
    , ack0 => op(207)
    , reset => reset
    , clk => clk);

  oper_tmp_d_20299_bool : libgt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_12_int_d_wire -- in
    , ip1 => tc_i_d_4_d_0_d_wire -- in
    , op => oper_tmp_d_20299_bool_d_wire -- out
    , req0 => ip(238)
    , ack0 => op(235)
    , reset => reset
    , clk => clk);

  oper_tmp_d_202_bool : libgt_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => indvar148_mux_1_d_wire -- in
    , ip1 => cst_74_uint_d_wire -- in
    , op => oper_tmp_d_202_bool_d_wire -- out
    , req0 => ip(224)
    , ack0 => op(221)
    , reset => reset
    , clk => clk);

  oper_tmp_d_206_d_lvl_d_0_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_l_array_d_wire -- in
    , ip1 => tc_tmp_d_206_d_id_d_0_d_cast_d_wire -- in
    , op => oper_tmp_d_206_d_lvl_d_0_uint_d_wire -- out
    , req0 => ip(231)
    , ack0 => op(228)
    , reset => reset
    , clk => clk);

  oper_tmp_d_20_d_lvl_d_0_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_rcoeff_d_wire -- in
    , ip1 => indvar121_mux_1_d_wire -- in
    , op => oper_tmp_d_20_d_lvl_d_0_uint_d_wire -- out
    , req0 => ip(26)
    , ack0 => op(26)
    , reset => reset
    , clk => clk);

  oper_tmp_d_210_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar148_mux_1_d_wire -- in
    , ip1 => cst_76_uint_d_wire -- in
    , op => oper_tmp_d_210_d_id_d_1_uint_d_wire -- out
    , req0 => ip(232)
    , ack0 => op(229)
    , reset => reset
    , clk => clk);

  oper_tmp_d_210_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_L_d_wire -- in
    , ip1 => oper_tmp_d_210_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_210_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(233)
    , ack0 => op(230)
    , reset => reset
    , clk => clk);

  oper_tmp_d_210_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_210_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar146_mux_1_d_wire -- in
    , op => oper_tmp_d_210_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(234)
    , ack0 => op(231)
    , reset => reset
    , clk => clk);

  oper_tmp_d_221111_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_inc_d_15_int_d_wire -- in
    , ip1 => cst_88_int_d_wire -- in
    , op => oper_tmp_d_221111_bool_d_wire -- out
    , req0 => ip(268)
    , ack0 => op(264)
    , reset => reset
    , clk => clk);

  oper_tmp_d_221_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => tc_i_d_5_d_0_d_wire -- in
    , ip1 => cst_84_int_d_wire -- in
    , op => oper_tmp_d_221_bool_d_wire -- out
    , req0 => ip(252)
    , ack0 => op(248)
    , reset => reset
    , clk => clk);

  oper_tmp_d_225_d_lvl_d_0_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_u_array_d_wire -- in
    , ip1 => tc_tmp_d_225_d_id_d_0_d_cast_d_wire -- in
    , op => oper_tmp_d_225_d_lvl_d_0_uint_d_wire -- out
    , req0 => ip(261)
    , ack0 => op(257)
    , reset => reset
    , clk => clk);

  oper_tmp_d_229_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar153_mux_1_d_wire -- in
    , ip1 => cst_86_uint_d_wire -- in
    , op => oper_tmp_d_229_d_id_d_1_uint_d_wire -- out
    , req0 => ip(262)
    , ack0 => op(258)
    , reset => reset
    , clk => clk);

  oper_tmp_d_229_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_U_d_wire -- in
    , ip1 => oper_tmp_d_229_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_229_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(263)
    , ack0 => op(259)
    , reset => reset
    , clk => clk);

  oper_tmp_d_229_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_229_d_lvl_d_1_uint_d_wire -- in
    , ip1 => oper_tmp_d_155_uint_d_wire -- in
    , op => oper_tmp_d_229_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(264)
    , ack0 => op(260)
    , reset => reset
    , clk => clk);

  oper_tmp_d_25_d_lvl_d_0_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_ccoeff_d_wire -- in
    , ip1 => indvar121_mux_1_d_wire -- in
    , op => oper_tmp_d_25_d_lvl_d_0_uint_d_wire -- out
    , req0 => ip(28)
    , ack0 => op(28)
    , reset => reset
    , clk => clk);

  oper_tmp_d_27_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_tmp_d_27_d_id_d_1_d_cast_d_wire -- in
    , ip1 => cst_10_uint_d_wire -- in
    , op => oper_tmp_d_27_d_id_d_1_uint_d_wire -- out
    , req0 => ip(31)
    , ack0 => op(31)
    , reset => reset
    , clk => clk);

  oper_tmp_d_27_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_27_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_27_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(32)
    , ack0 => op(32)
    , reset => reset
    , clk => clk);

  oper_tmp_d_27_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_27_d_lvl_d_1_uint_d_wire -- in
    , ip1 => tc_tmp_d_27_d_id_d_2_d_cast_d_wire -- in
    , op => oper_tmp_d_27_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(34)
    , ack0 => op(34)
    , reset => reset
    , clk => clk);

  oper_tmp_d_30_d_lvl_d_0_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => load_A_d_wire -- in
    , ip1 => indvar121_mux_1_d_wire -- in
    , op => oper_tmp_d_30_d_lvl_d_0_uint_d_wire -- out
    , req0 => ip(35)
    , ack0 => op(35)
    , reset => reset
    , clk => clk);

  oper_tmp_d_4223_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_j_d_321_int_d_wire -- in
    , ip1 => cst_23_int_d_wire -- in
    , op => oper_tmp_d_4223_bool_d_wire -- out
    , req0 => ip(75)
    , ack0 => op(71)
    , reset => reset
    , clk => clk);

  oper_tmp_d_42_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_j_d_3_int_d_wire -- in
    , ip1 => cst_18_int_d_wire -- in
    , op => oper_tmp_d_42_bool_d_wire -- out
    , req0 => ip(57)
    , ack0 => op(53)
    , reset => reset
    , clk => clk);

  oper_tmp_d_47_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_125_uint_d_wire -- in
    , ip1 => cst_21_uint_d_wire -- in
    , op => oper_tmp_d_47_d_id_d_1_uint_d_wire -- out
    , req0 => ip(68)
    , ack0 => op(63)
    , reset => reset
    , clk => clk);

  oper_tmp_d_47_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_47_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_47_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(69)
    , ack0 => op(64)
    , reset => reset
    , clk => clk);

  oper_tmp_d_47_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_47_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar129_mux_1_d_wire -- in
    , op => oper_tmp_d_47_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(70)
    , ack0 => op(65)
    , reset => reset
    , clk => clk);

  oper_tmp_d_52_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar129_mux_1_d_wire -- in
    , ip1 => cst_16_uint_d_wire -- in
    , op => oper_tmp_d_52_d_id_d_1_uint_d_wire -- out
    , req0 => ip(49)
    , ack0 => op(47)
    , reset => reset
    , clk => clk);

  oper_tmp_d_52_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_52_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_52_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(50)
    , ack0 => op(48)
    , reset => reset
    , clk => clk);

  oper_tmp_d_52_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_52_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar129_mux_1_d_wire -- in
    , op => oper_tmp_d_52_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(51)
    , ack0 => op(49)
    , reset => reset
    , clk => clk);

  oper_tmp_d_54_bool : libgt_float
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => load_tmp_d_48_d_wire -- in
    , ip1 => load_tmp_d_53_d_wire -- in
    , op => oper_tmp_d_54_bool_d_wire -- out
    , req0 => ip(72)
    , ack0 => op(67)
    , reset => reset
    , clk => clk);

  oper_tmp_d_65_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => indvar129_mux_1_d_wire -- in
    , ip1 => cst_26_uint_d_wire -- in
    , op => oper_tmp_d_65_d_id_d_1_uint_d_wire -- out
    , req0 => ip(82)
    , ack0 => op(77)
    , reset => reset
    , clk => clk);

  oper_tmp_d_65_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_65_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_65_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(83)
    , ack0 => op(78)
    , reset => reset
    , clk => clk);

  oper_tmp_d_65_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_65_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar126_mux_1_d_wire -- in
    , op => oper_tmp_d_65_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(84)
    , ack0 => op(79)
    , reset => reset
    , clk => clk);

  oper_tmp_d_74_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_tmp_d_74_d_id_d_1_d_cast_d_wire -- in
    , ip1 => cst_27_uint_d_wire -- in
    , op => oper_tmp_d_74_d_id_d_1_uint_d_wire -- out
    , req0 => ip(87)
    , ack0 => op(82)
    , reset => reset
    , clk => clk);

  oper_tmp_d_74_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_74_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_74_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(88)
    , ack0 => op(83)
    , reset => reset
    , clk => clk);

  oper_tmp_d_74_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_74_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar126_mux_1_d_wire -- in
    , op => oper_tmp_d_74_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(89)
    , ack0 => op(84)
    , reset => reset
    , clk => clk);

  oper_tmp_d_92_bool : liblt_int
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 1)
  port map(
    ip0 => oper_k_d_1_int_d_wire -- in
    , ip1 => cst_41_int_d_wire -- in
    , op => oper_tmp_d_92_bool_d_wire -- out
    , req0 => ip(116)
    , ack0 => op(110)
    , reset => reset
    , clk => clk);

  oper_tmp_d_97_d_id_d_1_uint : libmul_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_tmp_d_97_d_id_d_1_d_cast_d_wire -- in
    , ip1 => cst_42_uint_d_wire -- in
    , op => oper_tmp_d_97_d_id_d_1_uint_d_wire -- out
    , req0 => ip(119)
    , ack0 => op(114)
    , reset => reset
    , clk => clk);

  oper_tmp_d_97_d_lvl_d_1_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => location_start_B_d_wire -- in
    , ip1 => oper_tmp_d_97_d_id_d_1_uint_d_wire -- in
    , op => oper_tmp_d_97_d_lvl_d_1_uint_d_wire -- out
    , req0 => ip(120)
    , ack0 => op(115)
    , reset => reset
    , clk => clk);

  oper_tmp_d_97_d_lvl_d_2_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => oper_tmp_d_97_d_lvl_d_1_uint_d_wire -- in
    , ip1 => indvar134_mux_1_d_wire -- in
    , op => oper_tmp_d_97_d_lvl_d_2_uint_d_wire -- out
    , req0 => ip(121)
    , ack0 => op(116)
    , reset => reset
    , clk => clk);

  oper_tmp_d_uint : libadd_uint
  generic map(
     ip0_wd => 32
    , ip1_wd => 32
    , op_wd => 32)
  port map(
    ip0 => tc_j_d_3_d_in_d_wire -- in
    , ip1 => cst_19_uint_d_wire -- in
    , op => oper_tmp_d_uint_d_wire -- out
    , req0 => ip(61)
    , ack0 => op(58)
    , reset => reset
    , clk => clk);

  start_call_divide_0_actual_0_wr : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_call_divide_0_actual_0_d_wire -- in
    , dp => load_tmp_d_103_d_wire -- in
    , req0 => ip(124)
    , ack0 => op(119)
    , mreq => store_reqs(0)
    , mack => store_acks(0)
    , maddr => store_addr(0)
    , mdata => store_data(0)
    , reset => reset
    , clk => clk);

  start_call_divide_0_actual_1_wr : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => location_start_call_divide_0_actual_1_d_wire -- in
    , dp => load_tmp_d_108_d_wire -- in
    , req0 => ip(125)
    , ack0 => op(120)
    , mreq => store_reqs(1)
    , mack => store_acks(1)
    , maddr => store_addr(1)
    , mdata => store_data(1)
    , reset => reset
    , clk => clk);

  store_0 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_11_d_lvl_d_2_uint_d_wire -- in
    , dp => cst_3_float_d_wire -- in
    , req0 => ip(14)
    , ack0 => op(12)
    , mreq => store_reqs(2)
    , mack => store_acks(2)
    , maddr => store_addr(2)
    , mdata => store_data(2)
    , reset => reset
    , clk => clk);

  store_1 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_27_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_31_d_wire -- in
    , req0 => ip(37)
    , ack0 => op(37)
    , mreq => store_reqs(3)
    , mack => store_acks(3)
    , maddr => store_addr(3)
    , mdata => store_data(3)
    , reset => reset
    , clk => clk);

  store_10 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_171_d_lvl_d_2_uint_d_wire -- in
    , dp => cst_65_float_d_wire -- in
    , req0 => ip(202)
    , ack0 => op(199)
    , mreq => store_reqs(4)
    , mack => store_acks(4)
    , maddr => store_addr(4)
    , mdata => store_data(4)
    , reset => reset
    , clk => clk);

  store_11 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_188_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_193_d_wire -- in
    , req0 => ip(212)
    , ack0 => op(209)
    , mreq => store_reqs(5)
    , mack => store_acks(5)
    , maddr => store_addr(5)
    , mdata => store_data(5)
    , reset => reset
    , clk => clk);

  store_12 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_206_d_lvl_d_0_uint_d_wire -- in
    , dp => load_tmp_d_211_d_wire -- in
    , req0 => ip(236)
    , ack0 => op(233)
    , mreq => store_reqs(6)
    , mack => store_acks(6)
    , maddr => store_addr(6)
    , mdata => store_data(6)
    , reset => reset
    , clk => clk);

  store_13 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_225_d_lvl_d_0_uint_d_wire -- in
    , dp => load_tmp_d_230_d_wire -- in
    , req0 => ip(266)
    , ack0 => op(262)
    , mreq => store_reqs(7)
    , mack => store_acks(7)
    , maddr => store_addr(7)
    , mdata => store_data(7)
    , reset => reset
    , clk => clk);

  store_2 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_65_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_75_d_wire -- in
    , req0 => ip(91)
    , ack0 => op(86)
    , mreq => store_reqs(8)
    , mack => store_acks(8)
    , maddr => store_addr(8)
    , mdata => store_data(8)
    , reset => reset
    , clk => clk);

  store_3 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_74_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_66_d_wire -- in
    , req0 => ip(92)
    , ack0 => op(87)
    , mreq => store_reqs(9)
    , mack => store_acks(9)
    , maddr => store_addr(9)
    , mdata => store_data(9)
    , reset => reset
    , clk => clk);

  store_4 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_97_d_lvl_d_2_uint_d_wire -- in
    , dp => load_start_call_divide_0_return_d_wire -- in
    , req0 => ip(127)
    , ack0 => op(122)
    , mreq => store_reqs(10)
    , mack => store_acks(10)
    , maddr => store_addr(10)
    , mdata => store_data(10)
    , reset => reset
    , clk => clk);

  store_5 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_118_d_lvl_d_2_uint_d_wire -- in
    , dp => oper_tmp_d_135_float_d_wire -- in
    , req0 => ip(146)
    , ack0 => op(141)
    , mreq => store_reqs(11)
    , mack => store_acks(11)
    , maddr => store_addr(11)
    , mdata => store_data(11)
    , reset => reset
    , clk => clk);

  store_6 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_154_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_159_d_wire -- in
    , req0 => ip(169)
    , ack0 => op(165)
    , mreq => store_reqs(12)
    , mack => store_acks(12)
    , maddr => store_addr(12)
    , mdata => store_data(12)
    , reset => reset
    , clk => clk);

  store_7 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_163_d_lvl_d_2_uint_d_wire -- in
    , dp => cst_56_float_d_wire -- in
    , req0 => ip(174)
    , ack0 => op(170)
    , mreq => store_reqs(13)
    , mack => store_acks(13)
    , maddr => store_addr(13)
    , mdata => store_data(13)
    , reset => reset
    , clk => clk);

  store_8 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_171_d_lvl_d_2_uint_d_wire -- in
    , dp => cst_60_float_d_wire -- in
    , req0 => ip(188)
    , ack0 => op(184)
    , mreq => store_reqs(14)
    , mack => store_acks(14)
    , maddr => store_addr(14)
    , mdata => store_data(14)
    , reset => reset
    , clk => clk);

  store_9 : libsto
  generic map(
     ap_wd => 32
    , dp_wd => 32)
  port map(
    ap => oper_tmp_d_175_d_lvl_d_2_uint_d_wire -- in
    , dp => load_tmp_d_180_d_wire -- in
    , req0 => ip(198)
    , ack0 => op(194)
    , mreq => store_reqs(15)
    , mack => store_acks(15)
    , maddr => store_addr(15)
    , mdata => store_data(15)
    , reset => reset
    , clk => clk);

  tc_i_d_1_d_0 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar121_mux_1_d_wire -- in
    , op => tc_i_d_1_d_0_d_wire -- out
    , req0 => ip(25)
    , ack0 => op(25)
    , reset => reset
    , clk => clk);

  tc_i_d_2_d_0_d_ph : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar129_mux_1_d_wire -- in
    , op => tc_i_d_2_d_0_d_ph_d_wire -- out
    , req0 => ip(48)
    , ack0 => op(46)
    , reset => reset
    , clk => clk);

  tc_i_d_3_d_0_d_ph : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar143_mux_1_d_wire -- in
    , op => tc_i_d_3_d_0_d_ph_d_wire -- out
    , req0 => ip(155)
    , ack0 => op(151)
    , reset => reset
    , clk => clk);

  tc_i_d_4_d_0 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar148_mux_1_d_wire -- in
    , op => tc_i_d_4_d_0_d_wire -- out
    , req0 => ip(223)
    , ack0 => op(220)
    , reset => reset
    , clk => clk);

  tc_i_d_5_d_0 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar153_mux_1_d_wire -- in
    , op => tc_i_d_5_d_0_d_wire -- out
    , req0 => ip(251)
    , ack0 => op(247)
    , reset => reset
    , clk => clk);

  tc_indvar138 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar138_mux_1_d_wire -- in
    , op => tc_indvar138_d_wire -- out
    , req0 => ip(113)
    , ack0 => op(107)
    , reset => reset
    , clk => clk);

  tc_indvar151 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar151_mux_1_d_wire -- in
    , op => tc_indvar151_d_wire -- out
    , req0 => ip(256)
    , ack0 => op(252)
    , reset => reset
    , clk => clk);

  tc_j_d_11_d_2 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar146_mux_1_d_wire -- in
    , op => tc_j_d_11_d_2_d_wire -- out
    , req0 => ip(228)
    , ack0 => op(225)
    , reset => reset
    , clk => clk);

  tc_j_d_13_d_2 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_tmp_d_155_uint_d_wire -- in
    , op => tc_j_d_13_d_2_d_wire -- out
    , req0 => ip(258)
    , ack0 => op(254)
    , reset => reset
    , clk => clk);

  tc_j_d_3_d_2 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_tmp_d_125_uint_d_wire -- in
    , op => tc_j_d_3_d_2_d_wire -- out
    , req0 => ip(67)
    , ack0 => op(62)
    , reset => reset
    , clk => clk);

  tc_j_d_3_d_in : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_3_d_in_mux_1_d_wire -- in
    , op => tc_j_d_3_d_in_d_wire -- out
    , req0 => ip(59)
    , ack0 => op(56)
    , reset => reset
    , clk => clk);

  tc_j_d_7_d_1 : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_tmp_d_137_uint_d_wire -- in
    , op => tc_j_d_7_d_1_d_wire -- out
    , req0 => ip(133)
    , ack0 => op(128)
    , reset => reset
    , clk => clk);

  tc_p_d_0_d_0_d_ph : libcast_uint_to_int
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => indvar134_mux_1_d_wire -- in
    , op => tc_p_d_0_d_0_d_ph_d_wire -- out
    , req0 => ip(104)
    , ack0 => op(99)
    , reset => reset
    , clk => clk);

  tc_tmp_d_118_d_id_d_1_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_k_d_1_int_d_wire -- in
    , op => tc_tmp_d_118_d_id_d_1_d_cast_d_wire -- out
    , req0 => ip(134)
    , ack0 => op(129)
    , reset => reset
    , clk => clk);

  tc_tmp_d_154_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_154_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(162)
    , ack0 => op(158)
    , reset => reset
    , clk => clk);

  tc_tmp_d_158_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_158_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(166)
    , ack0 => op(162)
    , reset => reset
    , clk => clk);

  tc_tmp_d_163_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_163_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(172)
    , ack0 => op(168)
    , reset => reset
    , clk => clk);

  tc_tmp_d_171_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_171_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(185)
    , ack0 => op(180)
    , reset => reset
    , clk => clk);

  tc_tmp_d_175_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_175_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(191)
    , ack0 => op(187)
    , reset => reset
    , clk => clk);

  tc_tmp_d_179_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_179_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(195)
    , ack0 => op(191)
    , reset => reset
    , clk => clk);

  tc_tmp_d_188_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_188_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(205)
    , ack0 => op(202)
    , reset => reset
    , clk => clk);

  tc_tmp_d_192_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => j_d_9_d_2_mux_1_d_wire -- in
    , op => tc_tmp_d_192_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(209)
    , ack0 => op(206)
    , reset => reset
    , clk => clk);

  tc_tmp_d_206_d_id_d_0_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_k_d_2_d_2_int_d_wire -- in
    , op => tc_tmp_d_206_d_id_d_0_d_cast_d_wire -- out
    , req0 => ip(230)
    , ack0 => op(227)
    , reset => reset
    , clk => clk);

  tc_tmp_d_225_d_id_d_0_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_k_d_4_d_2_int_d_wire -- in
    , op => tc_tmp_d_225_d_id_d_0_d_cast_d_wire -- out
    , req0 => ip(260)
    , ack0 => op(256)
    , reset => reset
    , clk => clk);

  tc_tmp_d_27_d_id_d_1_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => load_tmp_d_21_d_wire -- in
    , op => tc_tmp_d_27_d_id_d_1_d_cast_d_wire -- out
    , req0 => ip(30)
    , ack0 => op(30)
    , reset => reset
    , clk => clk);

  tc_tmp_d_27_d_id_d_2_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => load_tmp_d_26_d_wire -- in
    , op => tc_tmp_d_27_d_id_d_2_d_cast_d_wire -- out
    , req0 => ip(33)
    , ack0 => op(33)
    , reset => reset
    , clk => clk);

  tc_tmp_d_74_d_id_d_1_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_wire -- in
    , op => tc_tmp_d_74_d_id_d_1_d_cast_d_wire -- out
    , req0 => ip(86)
    , ack0 => op(81)
    , reset => reset
    , clk => clk);

  tc_tmp_d_97_d_id_d_1_d_cast : libcast_int_to_uint
  generic map(
     ip_wd => 32
    , op_wd => 32)
  port map(
    ip => oper_k_d_1_int_d_wire -- in
    , op => tc_tmp_d_97_d_id_d_1_d_cast_d_wire -- out
    , req0 => ip(118)
    , ack0 => op(113)
    , reset => reset
    , clk => clk);

  cst_0_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_0_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_10_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_10_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_11_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_11_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_12_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_12_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_13_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_13_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_14_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_14_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_15_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_15_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_16_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_16_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_17_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_17_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_18_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_18_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_19_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_19_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_1_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_1_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_20_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_20_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_21_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_21_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_22_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_22_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_23_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_23_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_24_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_24_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_25_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_25_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_26_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_26_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_27_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_27_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_28_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_28_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_29_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_29_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_2_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_2_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_30_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_30_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_31_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_31_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_32_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_32_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_33_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_33_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_34_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_34_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_35_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_35_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_36_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_36_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_37_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_37_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_38_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_38_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_39_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_39_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_3_float : libkonst_float
  generic map(
    op_wd => 32
    , val => ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'))
  port map(
    op => cst_3_float_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_40_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_40_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_41_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_41_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_42_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_42_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_43_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_43_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_44_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_44_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_45_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_45_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_46_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_46_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_47_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_47_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_48_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_48_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_49_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_49_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_4_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_4_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_50_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 2)
  port map(
    op => cst_50_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_51_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_51_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_52_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_52_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_53_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_53_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_54_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_54_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_55_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_55_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_56_float : libkonst_float
  generic map(
    op_wd => 32
    , val => ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'))
  port map(
    op => cst_56_float_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_57_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_57_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_58_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_58_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_59_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_59_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_5_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_5_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_60_float : libkonst_float
  generic map(
    op_wd => 32
    , val => ('0','0','1','1','1','1','1','1','1','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'))
  port map(
    op => cst_60_float_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_61_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_61_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_62_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_62_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_63_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_63_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_64_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_64_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_65_float : libkonst_float
  generic map(
    op_wd => 32
    , val => ('0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0','0'))
  port map(
    op => cst_65_float_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_66_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_66_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_67_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_67_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_68_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_68_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_69_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_69_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_6_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_6_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_70_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_70_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_71_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_71_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_72_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_72_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_73_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_73_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_74_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 2147483647)
  port map(
    op => cst_74_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_75_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_75_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_76_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_76_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_77_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_77_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_78_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_78_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_79_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_79_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_7_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_7_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_80_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_80_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_81_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_81_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_82_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_82_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_83_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_83_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_84_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_84_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_85_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_85_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_86_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_86_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_87_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_87_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_88_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_88_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_89_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_89_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_8_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_8_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_90_int : libkonst_int
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_90_int_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_91_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => cst_91_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_92_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => cst_92_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  cst_9_uint : libkonst_uint
  generic map(
    op_wd => 32
    , val => 0)
  port map(
    op => cst_9_uint_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_B : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 10)
  port map(
    op => location_start_B_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_L : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 19)
  port map(
    op => location_start_L_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_U : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 28)
  port map(
    op => location_start_U_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_call_divide_0_actual_0 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 1)
  port map(
    op => location_start_call_divide_0_actual_0_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_call_divide_0_actual_1 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 2)
  port map(
    op => location_start_call_divide_0_actual_1_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_call_divide_0_return : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 3)
  port map(
    op => location_start_call_divide_0_return_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_0 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 4)
  port map(
    op => location_start_formal_0_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_1 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 5)
  port map(
    op => location_start_formal_1_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_2 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 6)
  port map(
    op => location_start_formal_2_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_3 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 7)
  port map(
    op => location_start_formal_3_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_4 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 8)
  port map(
    op => location_start_formal_4_d_wire -- out
    , reset => reset
    , clk => clk);

  location_start_formal_5 : libkonst_uint -- actually an address
  generic map(
    op_wd => 32
    , val => 9)
  port map(
    op => location_start_formal_5_d_wire -- out
    , reset => reset
    , clk => clk);
end Behavioral;
