library work;
use work.cpath_components.all;

entity divide_cp is
  port (

    ip    : in bit_vector(45 downto 1);
    op    : out bit_vector(51 downto 1) := (others => '0');
    reset : in bit;
    clk   : in bit);
end divide_cp;

architecture behavioral of divide_cp is

  signal place_1_tip : bit_vector(0 downto 0);
  signal place_1_rst : bit_vector(0 downto 0);
  signal place_1_top : bit;
  signal place_10_tip : bit_vector(0 downto 0);
  signal place_10_rst : bit_vector(0 downto 0);
  signal place_10_top : bit;
  signal place_101_tip : bit_vector(0 downto 0);
  signal place_101_rst : bit_vector(0 downto 0);
  signal place_101_top : bit;
  signal place_102_tip : bit_vector(1 downto 0);
  signal place_102_rst : bit_vector(0 downto 0);
  signal place_102_top : bit;
  signal place_103_tip : bit_vector(0 downto 0);
  signal place_103_rst : bit_vector(0 downto 0);
  signal place_103_top : bit;
  signal place_104_tip : bit_vector(0 downto 0);
  signal place_104_rst : bit_vector(0 downto 0);
  signal place_104_top : bit;
  signal place_105_tip : bit_vector(0 downto 0);
  signal place_105_rst : bit_vector(0 downto 0);
  signal place_105_top : bit;
  signal place_106_tip : bit_vector(1 downto 0);
  signal place_106_rst : bit_vector(0 downto 0);
  signal place_106_top : bit;
  signal place_107_tip : bit_vector(0 downto 0);
  signal place_107_rst : bit_vector(0 downto 0);
  signal place_107_top : bit;
  signal place_108_tip : bit_vector(0 downto 0);
  signal place_108_rst : bit_vector(0 downto 0);
  signal place_108_top : bit;
  signal place_109_tip : bit_vector(0 downto 0);
  signal place_109_rst : bit_vector(0 downto 0);
  signal place_109_top : bit;
  signal place_11_tip : bit_vector(0 downto 0);
  signal place_11_rst : bit_vector(0 downto 0);
  signal place_11_top : bit;
  signal place_110_tip : bit_vector(1 downto 0);
  signal place_110_rst : bit_vector(0 downto 0);
  signal place_110_top : bit;
  signal place_111_tip : bit_vector(0 downto 0);
  signal place_111_rst : bit_vector(0 downto 0);
  signal place_111_top : bit;
  signal place_112_tip : bit_vector(0 downto 0);
  signal place_112_rst : bit_vector(0 downto 0);
  signal place_112_top : bit;
  signal place_113_tip : bit_vector(0 downto 0);
  signal place_113_rst : bit_vector(0 downto 0);
  signal place_113_top : bit;
  signal place_114_tip : bit_vector(0 downto 0);
  signal place_114_rst : bit_vector(0 downto 0);
  signal place_114_top : bit;
  signal place_115_tip : bit_vector(0 downto 0);
  signal place_115_rst : bit_vector(0 downto 0);
  signal place_115_top : bit;
  signal place_116_tip : bit_vector(0 downto 0);
  signal place_116_rst : bit_vector(0 downto 0);
  signal place_116_top : bit;
  signal place_117_tip : bit_vector(0 downto 0);
  signal place_117_rst : bit_vector(0 downto 0);
  signal place_117_top : bit;
  signal place_118_tip : bit_vector(0 downto 0);
  signal place_118_rst : bit_vector(0 downto 0);
  signal place_118_top : bit;
  signal place_119_tip : bit_vector(0 downto 0);
  signal place_119_rst : bit_vector(0 downto 0);
  signal place_119_top : bit;
  signal place_120_tip : bit_vector(0 downto 0);
  signal place_120_rst : bit_vector(0 downto 0);
  signal place_120_top : bit;
  signal place_121_tip : bit_vector(0 downto 0);
  signal place_121_rst : bit_vector(0 downto 0);
  signal place_121_top : bit;
  signal place_122_tip : bit_vector(0 downto 0);
  signal place_122_rst : bit_vector(0 downto 0);
  signal place_122_top : bit;
  signal place_123_tip : bit_vector(0 downto 0);
  signal place_123_rst : bit_vector(0 downto 0);
  signal place_123_top : bit;
  signal place_124_tip : bit_vector(0 downto 0);
  signal place_124_rst : bit_vector(0 downto 0);
  signal place_124_top : bit;
  signal place_125_tip : bit_vector(0 downto 0);
  signal place_125_rst : bit_vector(1 downto 0);
  signal place_125_top : bit;
  signal place_128_tip : bit_vector(1 downto 0);
  signal place_128_rst : bit_vector(0 downto 0);
  signal place_128_top : bit;
  signal place_129_tip : bit_vector(0 downto 0);
  signal place_129_rst : bit_vector(0 downto 0);
  signal place_129_top : bit;
  signal place_13_tip : bit_vector(0 downto 0);
  signal place_13_rst : bit_vector(0 downto 0);
  signal place_13_top : bit;
  signal place_130_tip : bit_vector(0 downto 0);
  signal place_130_rst : bit_vector(0 downto 0);
  signal place_130_top : bit;
  signal place_131_tip : bit_vector(0 downto 0);
  signal place_131_rst : bit_vector(0 downto 0);
  signal place_131_top : bit;
  signal place_15_tip : bit_vector(0 downto 0);
  signal place_15_rst : bit_vector(0 downto 0);
  signal place_15_top : bit;
  signal place_17_tip : bit_vector(0 downto 0);
  signal place_17_rst : bit_vector(0 downto 0);
  signal place_17_top : bit;
  signal place_19_tip : bit_vector(0 downto 0);
  signal place_19_rst : bit_vector(0 downto 0);
  signal place_19_top : bit;
  signal place_2_tip : bit_vector(0 downto 0);
  signal place_2_rst : bit_vector(0 downto 0);
  signal place_2_top : bit;
  signal place_20_tip : bit_vector(0 downto 0);
  signal place_20_rst : bit_vector(0 downto 0);
  signal place_20_top : bit;
  signal place_21_tip : bit_vector(0 downto 0);
  signal place_21_rst : bit_vector(0 downto 0);
  signal place_21_top : bit;
  signal place_22_tip : bit_vector(0 downto 0);
  signal place_22_rst : bit_vector(0 downto 0);
  signal place_22_top : bit;
  signal place_23_tip : bit_vector(0 downto 0);
  signal place_23_rst : bit_vector(0 downto 0);
  signal place_23_top : bit;
  signal place_24_tip : bit_vector(0 downto 0);
  signal place_24_rst : bit_vector(0 downto 0);
  signal place_24_top : bit;
  signal place_25_tip : bit_vector(0 downto 0);
  signal place_25_rst : bit_vector(0 downto 0);
  signal place_25_top : bit;
  signal place_26_tip : bit_vector(0 downto 0);
  signal place_26_rst : bit_vector(0 downto 0);
  signal place_26_top : bit;
  signal place_28_tip : bit_vector(0 downto 0);
  signal place_28_rst : bit_vector(0 downto 0);
  signal place_28_top : bit;
  signal place_29_tip : bit_vector(0 downto 0);
  signal place_29_rst : bit_vector(1 downto 0);
  signal place_29_top : bit;
  signal place_31_tip : bit_vector(0 downto 0);
  signal place_31_rst : bit_vector(0 downto 0);
  signal place_31_top : bit;
  signal place_32_tip : bit_vector(1 downto 0);
  signal place_32_rst : bit_vector(0 downto 0);
  signal place_32_top : bit;
  signal place_33_tip : bit_vector(0 downto 0);
  signal place_33_rst : bit_vector(0 downto 0);
  signal place_33_top : bit;
  signal place_34_tip : bit_vector(0 downto 0);
  signal place_34_rst : bit_vector(0 downto 0);
  signal place_34_top : bit;
  signal place_35_tip : bit_vector(0 downto 0);
  signal place_35_rst : bit_vector(0 downto 0);
  signal place_35_top : bit;
  signal place_36_tip : bit_vector(1 downto 0);
  signal place_36_rst : bit_vector(0 downto 0);
  signal place_36_top : bit;
  signal place_37_tip : bit_vector(0 downto 0);
  signal place_37_rst : bit_vector(0 downto 0);
  signal place_37_top : bit;
  signal place_38_tip : bit_vector(0 downto 0);
  signal place_38_rst : bit_vector(0 downto 0);
  signal place_38_top : bit;
  signal place_39_tip : bit_vector(0 downto 0);
  signal place_39_rst : bit_vector(0 downto 0);
  signal place_39_top : bit;
  signal place_4_tip : bit_vector(0 downto 0);
  signal place_4_rst : bit_vector(0 downto 0);
  signal place_4_top : bit;
  signal place_40_tip : bit_vector(0 downto 0);
  signal place_40_rst : bit_vector(0 downto 0);
  signal place_40_top : bit;
  signal place_41_tip : bit_vector(0 downto 0);
  signal place_41_rst : bit_vector(0 downto 0);
  signal place_41_top : bit;
  signal place_42_tip : bit_vector(0 downto 0);
  signal place_42_rst : bit_vector(0 downto 0);
  signal place_42_top : bit;
  signal place_43_tip : bit_vector(0 downto 0);
  signal place_43_rst : bit_vector(0 downto 0);
  signal place_43_top : bit;
  signal place_44_tip : bit_vector(0 downto 0);
  signal place_44_rst : bit_vector(0 downto 0);
  signal place_44_top : bit;
  signal place_45_tip : bit_vector(0 downto 0);
  signal place_45_rst : bit_vector(0 downto 0);
  signal place_45_top : bit;
  signal place_46_tip : bit_vector(0 downto 0);
  signal place_46_rst : bit_vector(0 downto 0);
  signal place_46_top : bit;
  signal place_47_tip : bit_vector(0 downto 0);
  signal place_47_rst : bit_vector(1 downto 0);
  signal place_47_top : bit;
  signal place_49_tip : bit_vector(0 downto 0);
  signal place_49_rst : bit_vector(0 downto 0);
  signal place_49_top : bit;
  signal place_5_tip : bit_vector(0 downto 0);
  signal place_5_rst : bit_vector(0 downto 0);
  signal place_5_top : bit;
  signal place_50_tip : bit_vector(1 downto 0);
  signal place_50_rst : bit_vector(0 downto 0);
  signal place_50_top : bit;
  signal place_51_tip : bit_vector(0 downto 0);
  signal place_51_rst : bit_vector(0 downto 0);
  signal place_51_top : bit;
  signal place_52_tip : bit_vector(0 downto 0);
  signal place_52_rst : bit_vector(0 downto 0);
  signal place_52_top : bit;
  signal place_53_tip : bit_vector(0 downto 0);
  signal place_53_rst : bit_vector(0 downto 0);
  signal place_53_top : bit;
  signal place_54_tip : bit_vector(1 downto 0);
  signal place_54_rst : bit_vector(0 downto 0);
  signal place_54_top : bit;
  signal place_55_tip : bit_vector(0 downto 0);
  signal place_55_rst : bit_vector(0 downto 0);
  signal place_55_top : bit;
  signal place_56_tip : bit_vector(0 downto 0);
  signal place_56_rst : bit_vector(0 downto 0);
  signal place_56_top : bit;
  signal place_57_tip : bit_vector(0 downto 0);
  signal place_57_rst : bit_vector(0 downto 0);
  signal place_57_top : bit;
  signal place_58_tip : bit_vector(0 downto 0);
  signal place_58_rst : bit_vector(0 downto 0);
  signal place_58_top : bit;
  signal place_59_tip : bit_vector(0 downto 0);
  signal place_59_rst : bit_vector(0 downto 0);
  signal place_59_top : bit;
  signal place_60_tip : bit_vector(0 downto 0);
  signal place_60_rst : bit_vector(0 downto 0);
  signal place_60_top : bit;
  signal place_61_tip : bit_vector(0 downto 0);
  signal place_61_rst : bit_vector(1 downto 0);
  signal place_61_top : bit;
  signal place_63_tip : bit_vector(0 downto 0);
  signal place_63_rst : bit_vector(0 downto 0);
  signal place_63_top : bit;
  signal place_64_tip : bit_vector(1 downto 0);
  signal place_64_rst : bit_vector(0 downto 0);
  signal place_64_top : bit;
  signal place_65_tip : bit_vector(0 downto 0);
  signal place_65_rst : bit_vector(0 downto 0);
  signal place_65_top : bit;
  signal place_66_tip : bit_vector(0 downto 0);
  signal place_66_rst : bit_vector(0 downto 0);
  signal place_66_top : bit;
  signal place_67_tip : bit_vector(0 downto 0);
  signal place_67_rst : bit_vector(0 downto 0);
  signal place_67_top : bit;
  signal place_68_tip : bit_vector(1 downto 0);
  signal place_68_rst : bit_vector(0 downto 0);
  signal place_68_top : bit;
  signal place_69_tip : bit_vector(0 downto 0);
  signal place_69_rst : bit_vector(0 downto 0);
  signal place_69_top : bit;
  signal place_7_tip : bit_vector(0 downto 0);
  signal place_7_rst : bit_vector(0 downto 0);
  signal place_7_top : bit;
  signal place_70_tip : bit_vector(0 downto 0);
  signal place_70_rst : bit_vector(0 downto 0);
  signal place_70_top : bit;
  signal place_71_tip : bit_vector(0 downto 0);
  signal place_71_rst : bit_vector(0 downto 0);
  signal place_71_top : bit;
  signal place_72_tip : bit_vector(0 downto 0);
  signal place_72_rst : bit_vector(0 downto 0);
  signal place_72_top : bit;
  signal place_73_tip : bit_vector(0 downto 0);
  signal place_73_rst : bit_vector(0 downto 0);
  signal place_73_top : bit;
  signal place_74_tip : bit_vector(0 downto 0);
  signal place_74_rst : bit_vector(0 downto 0);
  signal place_74_top : bit;
  signal place_75_tip : bit_vector(0 downto 0);
  signal place_75_rst : bit_vector(0 downto 0);
  signal place_75_top : bit;
  signal place_76_tip : bit_vector(0 downto 0);
  signal place_76_rst : bit_vector(0 downto 0);
  signal place_76_top : bit;
  signal place_77_tip : bit_vector(0 downto 0);
  signal place_77_rst : bit_vector(0 downto 0);
  signal place_77_top : bit;
  signal place_78_tip : bit_vector(0 downto 0);
  signal place_78_rst : bit_vector(0 downto 0);
  signal place_78_top : bit;
  signal place_79_tip : bit_vector(0 downto 0);
  signal place_79_rst : bit_vector(1 downto 0);
  signal place_79_top : bit;
  signal place_81_tip : bit_vector(0 downto 0);
  signal place_81_rst : bit_vector(0 downto 0);
  signal place_81_top : bit;
  signal place_82_tip : bit_vector(1 downto 0);
  signal place_82_rst : bit_vector(0 downto 0);
  signal place_82_top : bit;
  signal place_83_tip : bit_vector(0 downto 0);
  signal place_83_rst : bit_vector(0 downto 0);
  signal place_83_top : bit;
  signal place_84_tip : bit_vector(0 downto 0);
  signal place_84_rst : bit_vector(0 downto 0);
  signal place_84_top : bit;
  signal place_85_tip : bit_vector(0 downto 0);
  signal place_85_rst : bit_vector(0 downto 0);
  signal place_85_top : bit;
  signal place_86_tip : bit_vector(1 downto 0);
  signal place_86_rst : bit_vector(0 downto 0);
  signal place_86_top : bit;
  signal place_87_tip : bit_vector(0 downto 0);
  signal place_87_rst : bit_vector(0 downto 0);
  signal place_87_top : bit;
  signal place_88_tip : bit_vector(0 downto 0);
  signal place_88_rst : bit_vector(0 downto 0);
  signal place_88_top : bit;
  signal place_89_tip : bit_vector(0 downto 0);
  signal place_89_rst : bit_vector(0 downto 0);
  signal place_89_top : bit;
  signal place_9_tip : bit_vector(0 downto 0);
  signal place_9_rst : bit_vector(0 downto 0);
  signal place_9_top : bit;
  signal place_90_tip : bit_vector(0 downto 0);
  signal place_90_rst : bit_vector(0 downto 0);
  signal place_90_top : bit;
  signal place_91_tip : bit_vector(0 downto 0);
  signal place_91_rst : bit_vector(0 downto 0);
  signal place_91_top : bit;
  signal place_92_tip : bit_vector(0 downto 0);
  signal place_92_rst : bit_vector(0 downto 0);
  signal place_92_top : bit;
  signal place_93_tip : bit_vector(0 downto 0);
  signal place_93_rst : bit_vector(0 downto 0);
  signal place_93_top : bit;
  signal place_94_tip : bit_vector(0 downto 0);
  signal place_94_rst : bit_vector(0 downto 0);
  signal place_94_top : bit;
  signal place_95_tip : bit_vector(0 downto 0);
  signal place_95_rst : bit_vector(0 downto 0);
  signal place_95_top : bit;
  signal place_96_tip : bit_vector(0 downto 0);
  signal place_96_rst : bit_vector(0 downto 0);
  signal place_96_top : bit;
  signal place_97_tip : bit_vector(0 downto 0);
  signal place_97_rst : bit_vector(0 downto 0);
  signal place_97_top : bit;
  signal place_98_tip : bit_vector(0 downto 0);
  signal place_98_rst : bit_vector(0 downto 0);
  signal place_98_top : bit;
  signal place_99_tip : bit_vector(0 downto 0);
  signal place_99_rst : bit_vector(1 downto 0);
  signal place_99_top : bit;

  signal cbr_0_oper_tmp_d_35_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_0_oper_tmp_d_35_bool_d_req_ge : bit;
  signal cbr_0_oper_tmp_d_35_bool_d_req_top : bit;
  signal cbr_1_oper_tmp_d_3_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_1_oper_tmp_d_3_bool_d_req_ge : bit;
  signal cbr_1_oper_tmp_d_3_bool_d_req_top : bit;
  signal cbr_2_oper_tmp_d_11_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_2_oper_tmp_d_11_bool_d_req_ge : bit;
  signal cbr_2_oper_tmp_d_11_bool_d_req_top : bit;
  signal cbr_3_oper_tmp_d_1114_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_3_oper_tmp_d_1114_bool_d_req_ge : bit;
  signal cbr_3_oper_tmp_d_1114_bool_d_req_top : bit;
  signal cbr_4_oper_tmp_d_2621_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_4_oper_tmp_d_2621_bool_d_req_ge : bit;
  signal cbr_4_oper_tmp_d_2621_bool_d_req_top : bit;
  signal cbr_5_oper_tmp_d_26_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_5_oper_tmp_d_26_bool_d_req_ge : bit;
  signal cbr_5_oper_tmp_d_26_bool_d_req_top : bit;
  signal di_d_0_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal di_d_0_d_0_mux_1_d_ack_ge : bit;
  signal di_d_0_d_0_mux_1_d_ack_top : bit;
  signal di_d_0_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal di_d_0_d_0_mux_1_d_req0_ge : bit;
  signal di_d_0_d_0_mux_1_d_req0_top : bit;
  signal di_d_0_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal di_d_0_d_0_mux_1_d_req1_ge : bit;
  signal di_d_0_d_0_mux_1_d_req1_top : bit;
  signal di_d_1_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal di_d_1_d_0_mux_1_d_ack_ge : bit;
  signal di_d_1_d_0_mux_1_d_ack_top : bit;
  signal di_d_1_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal di_d_1_d_0_mux_1_d_req0_ge : bit;
  signal di_d_1_d_0_mux_1_d_req0_top : bit;
  signal di_d_1_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal di_d_1_d_0_mux_1_d_req1_ge : bit;
  signal di_d_1_d_0_mux_1_d_req1_top : bit;
  signal di_d_1_d_1_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal di_d_1_d_1_mux_1_d_ack_ge : bit;
  signal di_d_1_d_1_mux_1_d_ack_top : bit;
  signal di_d_1_d_1_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal di_d_1_d_1_mux_1_d_req0_ge : bit;
  signal di_d_1_d_1_mux_1_d_req0_top : bit;
  signal di_d_1_d_1_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal di_d_1_d_1_mux_1_d_req1_ge : bit;
  signal di_d_1_d_1_mux_1_d_req1_top : bit;
  signal di_d_1_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal di_d_1_mux_1_d_ack_ge : bit;
  signal di_d_1_mux_1_d_ack_top : bit;
  signal di_d_1_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal di_d_1_mux_1_d_req0_ge : bit;
  signal di_d_1_mux_1_d_req0_top : bit;
  signal di_d_1_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal di_d_1_mux_1_d_req1_ge : bit;
  signal di_d_1_mux_1_d_req1_top : bit;
  signal di_d_2_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal di_d_2_d_0_mux_1_d_ack_ge : bit;
  signal di_d_2_d_0_mux_1_d_ack_top : bit;
  signal di_d_2_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal di_d_2_d_0_mux_1_d_req0_ge : bit;
  signal di_d_2_d_0_mux_1_d_req0_top : bit;
  signal di_d_2_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal di_d_2_d_0_mux_1_d_req1_ge : bit;
  signal di_d_2_d_0_mux_1_d_req1_top : bit;
  signal entry_to_loopentry_d_1_src_tip : bit_vector(0 downto 0);
  signal entry_to_loopentry_d_1_src_ge : bit;
  signal entry_to_loopentry_d_1_src_top : bit;
  signal entry_to_no_exit_d_0_d_preheader_src_tip : bit_vector(0 downto 0);
  signal entry_to_no_exit_d_0_d_preheader_src_ge : bit;
  signal entry_to_no_exit_d_0_d_preheader_src_top : bit;
  signal fin_tip : bit_vector(0 downto 0);
  signal fin_ge : bit;
  signal fin_top : bit;
  signal init_tip : bit_vector(0 downto 0);
  signal init_ge : bit;
  signal init_top : bit;
  signal load_dividend_d_ack_tip : bit_vector(0 downto 0);
  signal load_dividend_d_ack_ge : bit;
  signal load_dividend_d_ack_top : bit;
  signal load_dividend_d_req_tip : bit_vector(0 downto 0);
  signal load_dividend_d_req_ge : bit;
  signal load_dividend_d_req_top : bit;
  signal load_divisor_d_ack_tip : bit_vector(0 downto 0);
  signal load_divisor_d_ack_ge : bit;
  signal load_divisor_d_ack_top : bit;
  signal load_divisor_d_req_tip : bit_vector(0 downto 0);
  signal load_divisor_d_req_ge : bit;
  signal load_divisor_d_req_top : bit;
  signal loopentry_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_1_d_entry_ge : bit;
  signal loopentry_d_1_d_entry_top : bit;
  signal loopentry_d_1_d_loopexit_to_loopentry_d_1_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_1_d_loopexit_to_loopentry_d_1_src_ge : bit;
  signal loopentry_d_1_d_loopexit_to_loopentry_d_1_src_top : bit;
  signal loopentry_d_1_d_pre_tip : bit_vector(1 downto 0);
  signal loopentry_d_1_d_pre_ge : bit;
  signal loopentry_d_1_d_pre_top : bit;
  signal loopentry_d_1_to_loopexit_d_1_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_1_to_loopexit_d_1_src_ge : bit;
  signal loopentry_d_1_to_loopexit_d_1_src_top : bit;
  signal loopentry_d_1_to_no_exit_d_1_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_1_to_no_exit_d_1_d_preheader_src_ge : bit;
  signal loopentry_d_1_to_no_exit_d_1_d_preheader_src_top : bit;
  signal loopexit_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_d_entry_ge : bit;
  signal loopexit_d_1_d_entry_top : bit;
  signal loopexit_d_1_d_loopexit_to_loopexit_d_1_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_d_loopexit_to_loopexit_d_1_src_ge : bit;
  signal loopexit_d_1_d_loopexit_to_loopexit_d_1_src_top : bit;
  signal loopexit_d_1_d_pre_tip : bit_vector(1 downto 0);
  signal loopexit_d_1_d_pre_ge : bit;
  signal loopexit_d_1_d_pre_top : bit;
  signal loopexit_d_1_to_loopexit_d_2_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_to_loopexit_d_2_src_ge : bit;
  signal loopexit_d_1_to_loopexit_d_2_src_top : bit;
  signal loopexit_d_1_to_no_exit_d_2_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_to_no_exit_d_2_d_preheader_src_ge : bit;
  signal loopexit_d_1_to_no_exit_d_2_d_preheader_src_top : bit;
  signal ni_d_0_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_0_d_0_mux_1_d_ack_ge : bit;
  signal ni_d_0_d_0_mux_1_d_ack_top : bit;
  signal ni_d_0_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_0_d_0_mux_1_d_req0_ge : bit;
  signal ni_d_0_d_0_mux_1_d_req0_top : bit;
  signal ni_d_0_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_0_d_0_mux_1_d_req1_ge : bit;
  signal ni_d_0_d_0_mux_1_d_req1_top : bit;
  signal ni_d_1_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_0_mux_1_d_ack_ge : bit;
  signal ni_d_1_d_0_mux_1_d_ack_top : bit;
  signal ni_d_1_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_0_mux_1_d_req0_ge : bit;
  signal ni_d_1_d_0_mux_1_d_req0_top : bit;
  signal ni_d_1_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_0_mux_1_d_req1_ge : bit;
  signal ni_d_1_d_0_mux_1_d_req1_top : bit;
  signal ni_d_1_d_1_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_1_mux_1_d_ack_ge : bit;
  signal ni_d_1_d_1_mux_1_d_ack_top : bit;
  signal ni_d_1_d_1_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_1_mux_1_d_req0_ge : bit;
  signal ni_d_1_d_1_mux_1_d_req0_top : bit;
  signal ni_d_1_d_1_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_1_d_1_mux_1_d_req1_ge : bit;
  signal ni_d_1_d_1_mux_1_d_req1_top : bit;
  signal ni_d_1_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_1_mux_1_d_ack_ge : bit;
  signal ni_d_1_mux_1_d_ack_top : bit;
  signal ni_d_1_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_1_mux_1_d_req0_ge : bit;
  signal ni_d_1_mux_1_d_req0_top : bit;
  signal ni_d_1_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_1_mux_1_d_req1_ge : bit;
  signal ni_d_1_mux_1_d_req1_top : bit;
  signal ni_d_2_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_0_mux_1_d_ack_ge : bit;
  signal ni_d_2_d_0_mux_1_d_ack_top : bit;
  signal ni_d_2_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_0_mux_1_d_req0_ge : bit;
  signal ni_d_2_d_0_mux_1_d_req0_top : bit;
  signal ni_d_2_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_0_mux_1_d_req1_ge : bit;
  signal ni_d_2_d_0_mux_1_d_req1_top : bit;
  signal ni_d_2_d_1_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_1_mux_1_d_ack_ge : bit;
  signal ni_d_2_d_1_mux_1_d_ack_top : bit;
  signal ni_d_2_d_1_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_1_mux_1_d_req0_ge : bit;
  signal ni_d_2_d_1_mux_1_d_req0_top : bit;
  signal ni_d_2_d_1_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ni_d_2_d_1_mux_1_d_req1_ge : bit;
  signal ni_d_2_d_1_mux_1_d_req1_top : bit;
  signal no_exit_d_0_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_0_d_entry_ge : bit;
  signal no_exit_d_0_d_entry_top : bit;
  signal no_exit_d_0_d_pre_tip : bit_vector(1 downto 0);
  signal no_exit_d_0_d_pre_ge : bit;
  signal no_exit_d_0_d_pre_top : bit;
  signal no_exit_d_0_d_preheader_to_no_exit_d_0_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_0_d_preheader_to_no_exit_d_0_src_ge : bit;
  signal no_exit_d_0_d_preheader_to_no_exit_d_0_src_top : bit;
  signal no_exit_d_0_to_loopentry_d_1_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_0_to_loopentry_d_1_d_loopexit_src_ge : bit;
  signal no_exit_d_0_to_loopentry_d_1_d_loopexit_src_top : bit;
  signal no_exit_d_0_to_no_exit_d_0_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_0_to_no_exit_d_0_src_ge : bit;
  signal no_exit_d_0_to_no_exit_d_0_src_top : bit;
  signal no_exit_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_d_entry_ge : bit;
  signal no_exit_d_1_d_entry_top : bit;
  signal no_exit_d_1_d_pre_tip : bit_vector(1 downto 0);
  signal no_exit_d_1_d_pre_ge : bit;
  signal no_exit_d_1_d_pre_top : bit;
  signal no_exit_d_1_d_preheader_to_no_exit_d_1_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_d_preheader_to_no_exit_d_1_src_ge : bit;
  signal no_exit_d_1_d_preheader_to_no_exit_d_1_src_top : bit;
  signal no_exit_d_1_to_loopexit_d_1_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_to_loopexit_d_1_d_loopexit_src_ge : bit;
  signal no_exit_d_1_to_loopexit_d_1_d_loopexit_src_top : bit;
  signal no_exit_d_1_to_no_exit_d_1_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_to_no_exit_d_1_src_ge : bit;
  signal no_exit_d_1_to_no_exit_d_1_src_top : bit;
  signal no_exit_d_2_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_d_entry_ge : bit;
  signal no_exit_d_2_d_entry_top : bit;
  signal no_exit_d_2_d_pre_tip : bit_vector(2 downto 0);
  signal no_exit_d_2_d_pre_ge : bit;
  signal no_exit_d_2_d_pre_top : bit;
  signal no_exit_d_2_d_preheader_to_no_exit_d_2_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_d_preheader_to_no_exit_d_2_src_ge : bit;
  signal no_exit_d_2_d_preheader_to_no_exit_d_2_src_top : bit;
  signal no_exit_d_2_to_loopexit_d_2_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_to_loopexit_d_2_d_loopexit_src_ge : bit;
  signal no_exit_d_2_to_loopexit_d_2_d_loopexit_src_top : bit;
  signal no_exit_d_2_to_no_exit_d_2_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_to_no_exit_d_2_src_ge : bit;
  signal no_exit_d_2_to_no_exit_d_2_src_top : bit;
  signal oper_tmp_d_1114_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1114_bool_d_ack_ge : bit;
  signal oper_tmp_d_1114_bool_d_ack_top : bit;
  signal oper_tmp_d_1114_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1114_bool_d_req_ge : bit;
  signal oper_tmp_d_1114_bool_d_req_top : bit;
  signal oper_tmp_d_11_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_bool_d_ack_ge : bit;
  signal oper_tmp_d_11_bool_d_ack_top : bit;
  signal oper_tmp_d_11_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_bool_d_req_ge : bit;
  signal oper_tmp_d_11_bool_d_req_top : bit;
  signal oper_tmp_d_14_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14_float_d_ack_ge : bit;
  signal oper_tmp_d_14_float_d_ack_top : bit;
  signal oper_tmp_d_14_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14_float_d_req_ge : bit;
  signal oper_tmp_d_14_float_d_req_top : bit;
  signal oper_tmp_d_16_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_16_float_d_ack_ge : bit;
  signal oper_tmp_d_16_float_d_ack_top : bit;
  signal oper_tmp_d_16_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_16_float_d_req_ge : bit;
  signal oper_tmp_d_16_float_d_req_top : bit;
  signal oper_tmp_d_19_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_19_float_d_ack_ge : bit;
  signal oper_tmp_d_19_float_d_ack_top : bit;
  signal oper_tmp_d_19_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_19_float_d_req_ge : bit;
  signal oper_tmp_d_19_float_d_req_top : bit;
  signal oper_tmp_d_21_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_21_float_d_ack_ge : bit;
  signal oper_tmp_d_21_float_d_ack_top : bit;
  signal oper_tmp_d_21_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_21_float_d_req_ge : bit;
  signal oper_tmp_d_21_float_d_req_top : bit;
  signal oper_tmp_d_2420_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_2420_float_d_ack_ge : bit;
  signal oper_tmp_d_2420_float_d_ack_top : bit;
  signal oper_tmp_d_2420_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_2420_float_d_req_ge : bit;
  signal oper_tmp_d_2420_float_d_req_top : bit;
  signal oper_tmp_d_24_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_24_float_d_ack_ge : bit;
  signal oper_tmp_d_24_float_d_ack_top : bit;
  signal oper_tmp_d_24_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_24_float_d_req_ge : bit;
  signal oper_tmp_d_24_float_d_req_top : bit;
  signal oper_tmp_d_2621_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_2621_bool_d_ack_ge : bit;
  signal oper_tmp_d_2621_bool_d_ack_top : bit;
  signal oper_tmp_d_2621_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_2621_bool_d_req_ge : bit;
  signal oper_tmp_d_2621_bool_d_req_top : bit;
  signal oper_tmp_d_26_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_26_bool_d_ack_ge : bit;
  signal oper_tmp_d_26_bool_d_ack_top : bit;
  signal oper_tmp_d_26_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_26_bool_d_req_ge : bit;
  signal oper_tmp_d_26_bool_d_req_top : bit;
  signal oper_tmp_d_31_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_31_float_d_ack_ge : bit;
  signal oper_tmp_d_31_float_d_ack_top : bit;
  signal oper_tmp_d_31_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_31_float_d_req_ge : bit;
  signal oper_tmp_d_31_float_d_req_top : bit;
  signal oper_tmp_d_34_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_34_float_d_ack_ge : bit;
  signal oper_tmp_d_34_float_d_ack_top : bit;
  signal oper_tmp_d_34_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_34_float_d_req_ge : bit;
  signal oper_tmp_d_34_float_d_req_top : bit;
  signal oper_tmp_d_35_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_35_bool_d_ack_ge : bit;
  signal oper_tmp_d_35_bool_d_ack_top : bit;
  signal oper_tmp_d_35_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_35_bool_d_req_ge : bit;
  signal oper_tmp_d_35_bool_d_req_top : bit;
  signal oper_tmp_d_36_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_36_float_d_ack_ge : bit;
  signal oper_tmp_d_36_float_d_ack_top : bit;
  signal oper_tmp_d_36_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_36_float_d_req_ge : bit;
  signal oper_tmp_d_36_float_d_req_top : bit;
  signal oper_tmp_d_3_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_3_bool_d_ack_ge : bit;
  signal oper_tmp_d_3_bool_d_ack_top : bit;
  signal oper_tmp_d_3_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_3_bool_d_req_ge : bit;
  signal oper_tmp_d_3_bool_d_req_top : bit;
  signal oper_tmp_d_6_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_6_float_d_ack_ge : bit;
  signal oper_tmp_d_6_float_d_ack_top : bit;
  signal oper_tmp_d_6_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_6_float_d_req_ge : bit;
  signal oper_tmp_d_6_float_d_req_top : bit;
  signal oper_tmp_d_8_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_8_float_d_ack_ge : bit;
  signal oper_tmp_d_8_float_d_ack_top : bit;
  signal oper_tmp_d_8_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_8_float_d_req_ge : bit;
  signal oper_tmp_d_8_float_d_req_top : bit;
  signal ri_d_0_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ri_d_0_d_0_mux_1_d_ack_ge : bit;
  signal ri_d_0_d_0_mux_1_d_ack_top : bit;
  signal ri_d_0_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ri_d_0_d_0_mux_1_d_req0_ge : bit;
  signal ri_d_0_d_0_mux_1_d_req0_top : bit;
  signal ri_d_0_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ri_d_0_d_0_mux_1_d_req1_ge : bit;
  signal ri_d_0_d_0_mux_1_d_req1_top : bit;
  signal store_location_divide_return_d_ack_tip : bit_vector(0 downto 0);
  signal store_location_divide_return_d_ack_ge : bit;
  signal store_location_divide_return_d_ack_top : bit;
  signal store_location_divide_return_d_req_tip : bit_vector(0 downto 0);
  signal store_location_divide_return_d_req_ge : bit;
  signal store_location_divide_return_d_req_top : bit;

begin


  place_1 : place
  generic map(1, 1, '0')
  port map(place_1_tip, place_1_rst, place_1_top, reset, clk);

  place_10 : place
  generic map(1, 1, '0')
  port map(place_10_tip, place_10_rst, place_10_top, reset, clk);

  place_101 : place
  generic map(1, 1, '0')
  port map(place_101_tip, place_101_rst, place_101_top, reset, clk);

  place_102 : place
  generic map(2, 1, '0')
  port map(place_102_tip, place_102_rst, place_102_top, reset, clk);

  place_103 : place
  generic map(1, 1, '0')
  port map(place_103_tip, place_103_rst, place_103_top, reset, clk);

  place_104 : place
  generic map(1, 1, '0')
  port map(place_104_tip, place_104_rst, place_104_top, reset, clk);

  place_105 : place
  generic map(1, 1, '0')
  port map(place_105_tip, place_105_rst, place_105_top, reset, clk);

  place_106 : place
  generic map(2, 1, '0')
  port map(place_106_tip, place_106_rst, place_106_top, reset, clk);

  place_107 : place
  generic map(1, 1, '0')
  port map(place_107_tip, place_107_rst, place_107_top, reset, clk);

  place_108 : place
  generic map(1, 1, '0')
  port map(place_108_tip, place_108_rst, place_108_top, reset, clk);

  place_109 : place
  generic map(1, 1, '0')
  port map(place_109_tip, place_109_rst, place_109_top, reset, clk);

  place_11 : place
  generic map(1, 1, '0')
  port map(place_11_tip, place_11_rst, place_11_top, reset, clk);

  place_110 : place
  generic map(2, 1, '0')
  port map(place_110_tip, place_110_rst, place_110_top, reset, clk);

  place_111 : place
  generic map(1, 1, '0')
  port map(place_111_tip, place_111_rst, place_111_top, reset, clk);

  place_112 : place
  generic map(1, 1, '0')
  port map(place_112_tip, place_112_rst, place_112_top, reset, clk);

  place_113 : place
  generic map(1, 1, '0')
  port map(place_113_tip, place_113_rst, place_113_top, reset, clk);

  place_114 : place
  generic map(1, 1, '0')
  port map(place_114_tip, place_114_rst, place_114_top, reset, clk);

  place_115 : place
  generic map(1, 1, '0')
  port map(place_115_tip, place_115_rst, place_115_top, reset, clk);

  place_116 : place
  generic map(1, 1, '0')
  port map(place_116_tip, place_116_rst, place_116_top, reset, clk);

  place_117 : place
  generic map(1, 1, '0')
  port map(place_117_tip, place_117_rst, place_117_top, reset, clk);

  place_118 : place
  generic map(1, 1, '0')
  port map(place_118_tip, place_118_rst, place_118_top, reset, clk);

  place_119 : place
  generic map(1, 1, '0')
  port map(place_119_tip, place_119_rst, place_119_top, reset, clk);

  place_120 : place
  generic map(1, 1, '0')
  port map(place_120_tip, place_120_rst, place_120_top, reset, clk);

  place_121 : place
  generic map(1, 1, '0')
  port map(place_121_tip, place_121_rst, place_121_top, reset, clk);

  place_122 : place
  generic map(1, 1, '0')
  port map(place_122_tip, place_122_rst, place_122_top, reset, clk);

  place_123 : place
  generic map(1, 1, '0')
  port map(place_123_tip, place_123_rst, place_123_top, reset, clk);

  place_124 : place
  generic map(1, 1, '0')
  port map(place_124_tip, place_124_rst, place_124_top, reset, clk);

  place_125 : place
  generic map(1, 2, '0')
  port map(place_125_tip, place_125_rst, place_125_top, reset, clk);

  place_128 : place
  generic map(2, 1, '0')
  port map(place_128_tip, place_128_rst, place_128_top, reset, clk);

  place_129 : place
  generic map(1, 1, '0')
  port map(place_129_tip, place_129_rst, place_129_top, reset, clk);

  place_13 : place
  generic map(1, 1, '0')
  port map(place_13_tip, place_13_rst, place_13_top, reset, clk);

  place_130 : place
  generic map(1, 1, '0')
  port map(place_130_tip, place_130_rst, place_130_top, reset, clk);

  place_131 : place
  generic map(1, 1, '0')
  port map(place_131_tip, place_131_rst, place_131_top, reset, clk);

  place_15 : place
  generic map(1, 1, '0')
  port map(place_15_tip, place_15_rst, place_15_top, reset, clk);

  place_17 : place
  generic map(1, 1, '0')
  port map(place_17_tip, place_17_rst, place_17_top, reset, clk);

  place_19 : place
  generic map(1, 1, '0')
  port map(place_19_tip, place_19_rst, place_19_top, reset, clk);

  place_2 : place
  generic map(1, 1, '0')
  port map(place_2_tip, place_2_rst, place_2_top, reset, clk);

  place_20 : place
  generic map(1, 1, '1')
  port map(place_20_tip, place_20_rst, place_20_top, reset, clk);

  place_21 : place
  generic map(1, 1, '0')
  port map(place_21_tip, place_21_rst, place_21_top, reset, clk);

  place_22 : place
  generic map(1, 1, '0')
  port map(place_22_tip, place_22_rst, place_22_top, reset, clk);

  place_23 : place
  generic map(1, 1, '0')
  port map(place_23_tip, place_23_rst, place_23_top, reset, clk);

  place_24 : place
  generic map(1, 1, '0')
  port map(place_24_tip, place_24_rst, place_24_top, reset, clk);

  place_25 : place
  generic map(1, 1, '0')
  port map(place_25_tip, place_25_rst, place_25_top, reset, clk);

  place_26 : place
  generic map(1, 1, '0')
  port map(place_26_tip, place_26_rst, place_26_top, reset, clk);

  place_28 : place
  generic map(1, 1, '0')
  port map(place_28_tip, place_28_rst, place_28_top, reset, clk);

  place_29 : place
  generic map(1, 2, '0')
  port map(place_29_tip, place_29_rst, place_29_top, reset, clk);

  place_31 : place
  generic map(1, 1, '0')
  port map(place_31_tip, place_31_rst, place_31_top, reset, clk);

  place_32 : place
  generic map(2, 1, '0')
  port map(place_32_tip, place_32_rst, place_32_top, reset, clk);

  place_33 : place
  generic map(1, 1, '0')
  port map(place_33_tip, place_33_rst, place_33_top, reset, clk);

  place_34 : place
  generic map(1, 1, '0')
  port map(place_34_tip, place_34_rst, place_34_top, reset, clk);

  place_35 : place
  generic map(1, 1, '0')
  port map(place_35_tip, place_35_rst, place_35_top, reset, clk);

  place_36 : place
  generic map(2, 1, '0')
  port map(place_36_tip, place_36_rst, place_36_top, reset, clk);

  place_37 : place
  generic map(1, 1, '0')
  port map(place_37_tip, place_37_rst, place_37_top, reset, clk);

  place_38 : place
  generic map(1, 1, '0')
  port map(place_38_tip, place_38_rst, place_38_top, reset, clk);

  place_39 : place
  generic map(1, 1, '0')
  port map(place_39_tip, place_39_rst, place_39_top, reset, clk);

  place_4 : place
  generic map(1, 1, '0')
  port map(place_4_tip, place_4_rst, place_4_top, reset, clk);

  place_40 : place
  generic map(1, 1, '0')
  port map(place_40_tip, place_40_rst, place_40_top, reset, clk);

  place_41 : place
  generic map(1, 1, '0')
  port map(place_41_tip, place_41_rst, place_41_top, reset, clk);

  place_42 : place
  generic map(1, 1, '0')
  port map(place_42_tip, place_42_rst, place_42_top, reset, clk);

  place_43 : place
  generic map(1, 1, '0')
  port map(place_43_tip, place_43_rst, place_43_top, reset, clk);

  place_44 : place
  generic map(1, 1, '0')
  port map(place_44_tip, place_44_rst, place_44_top, reset, clk);

  place_45 : place
  generic map(1, 1, '0')
  port map(place_45_tip, place_45_rst, place_45_top, reset, clk);

  place_46 : place
  generic map(1, 1, '0')
  port map(place_46_tip, place_46_rst, place_46_top, reset, clk);

  place_47 : place
  generic map(1, 2, '0')
  port map(place_47_tip, place_47_rst, place_47_top, reset, clk);

  place_49 : place
  generic map(1, 1, '0')
  port map(place_49_tip, place_49_rst, place_49_top, reset, clk);

  place_5 : place
  generic map(1, 1, '0')
  port map(place_5_tip, place_5_rst, place_5_top, reset, clk);

  place_50 : place
  generic map(2, 1, '0')
  port map(place_50_tip, place_50_rst, place_50_top, reset, clk);

  place_51 : place
  generic map(1, 1, '0')
  port map(place_51_tip, place_51_rst, place_51_top, reset, clk);

  place_52 : place
  generic map(1, 1, '0')
  port map(place_52_tip, place_52_rst, place_52_top, reset, clk);

  place_53 : place
  generic map(1, 1, '0')
  port map(place_53_tip, place_53_rst, place_53_top, reset, clk);

  place_54 : place
  generic map(2, 1, '0')
  port map(place_54_tip, place_54_rst, place_54_top, reset, clk);

  place_55 : place
  generic map(1, 1, '0')
  port map(place_55_tip, place_55_rst, place_55_top, reset, clk);

  place_56 : place
  generic map(1, 1, '0')
  port map(place_56_tip, place_56_rst, place_56_top, reset, clk);

  place_57 : place
  generic map(1, 1, '0')
  port map(place_57_tip, place_57_rst, place_57_top, reset, clk);

  place_58 : place
  generic map(1, 1, '0')
  port map(place_58_tip, place_58_rst, place_58_top, reset, clk);

  place_59 : place
  generic map(1, 1, '0')
  port map(place_59_tip, place_59_rst, place_59_top, reset, clk);

  place_60 : place
  generic map(1, 1, '0')
  port map(place_60_tip, place_60_rst, place_60_top, reset, clk);

  place_61 : place
  generic map(1, 2, '0')
  port map(place_61_tip, place_61_rst, place_61_top, reset, clk);

  place_63 : place
  generic map(1, 1, '0')
  port map(place_63_tip, place_63_rst, place_63_top, reset, clk);

  place_64 : place
  generic map(2, 1, '0')
  port map(place_64_tip, place_64_rst, place_64_top, reset, clk);

  place_65 : place
  generic map(1, 1, '0')
  port map(place_65_tip, place_65_rst, place_65_top, reset, clk);

  place_66 : place
  generic map(1, 1, '0')
  port map(place_66_tip, place_66_rst, place_66_top, reset, clk);

  place_67 : place
  generic map(1, 1, '0')
  port map(place_67_tip, place_67_rst, place_67_top, reset, clk);

  place_68 : place
  generic map(2, 1, '0')
  port map(place_68_tip, place_68_rst, place_68_top, reset, clk);

  place_69 : place
  generic map(1, 1, '0')
  port map(place_69_tip, place_69_rst, place_69_top, reset, clk);

  place_7 : place
  generic map(1, 1, '0')
  port map(place_7_tip, place_7_rst, place_7_top, reset, clk);

  place_70 : place
  generic map(1, 1, '0')
  port map(place_70_tip, place_70_rst, place_70_top, reset, clk);

  place_71 : place
  generic map(1, 1, '0')
  port map(place_71_tip, place_71_rst, place_71_top, reset, clk);

  place_72 : place
  generic map(1, 1, '0')
  port map(place_72_tip, place_72_rst, place_72_top, reset, clk);

  place_73 : place
  generic map(1, 1, '0')
  port map(place_73_tip, place_73_rst, place_73_top, reset, clk);

  place_74 : place
  generic map(1, 1, '0')
  port map(place_74_tip, place_74_rst, place_74_top, reset, clk);

  place_75 : place
  generic map(1, 1, '0')
  port map(place_75_tip, place_75_rst, place_75_top, reset, clk);

  place_76 : place
  generic map(1, 1, '0')
  port map(place_76_tip, place_76_rst, place_76_top, reset, clk);

  place_77 : place
  generic map(1, 1, '0')
  port map(place_77_tip, place_77_rst, place_77_top, reset, clk);

  place_78 : place
  generic map(1, 1, '0')
  port map(place_78_tip, place_78_rst, place_78_top, reset, clk);

  place_79 : place
  generic map(1, 2, '0')
  port map(place_79_tip, place_79_rst, place_79_top, reset, clk);

  place_81 : place
  generic map(1, 1, '0')
  port map(place_81_tip, place_81_rst, place_81_top, reset, clk);

  place_82 : place
  generic map(2, 1, '0')
  port map(place_82_tip, place_82_rst, place_82_top, reset, clk);

  place_83 : place
  generic map(1, 1, '0')
  port map(place_83_tip, place_83_rst, place_83_top, reset, clk);

  place_84 : place
  generic map(1, 1, '0')
  port map(place_84_tip, place_84_rst, place_84_top, reset, clk);

  place_85 : place
  generic map(1, 1, '0')
  port map(place_85_tip, place_85_rst, place_85_top, reset, clk);

  place_86 : place
  generic map(2, 1, '0')
  port map(place_86_tip, place_86_rst, place_86_top, reset, clk);

  place_87 : place
  generic map(1, 1, '0')
  port map(place_87_tip, place_87_rst, place_87_top, reset, clk);

  place_88 : place
  generic map(1, 1, '0')
  port map(place_88_tip, place_88_rst, place_88_top, reset, clk);

  place_89 : place
  generic map(1, 1, '0')
  port map(place_89_tip, place_89_rst, place_89_top, reset, clk);

  place_9 : place
  generic map(1, 1, '0')
  port map(place_9_tip, place_9_rst, place_9_top, reset, clk);

  place_90 : place
  generic map(1, 1, '0')
  port map(place_90_tip, place_90_rst, place_90_top, reset, clk);

  place_91 : place
  generic map(1, 1, '0')
  port map(place_91_tip, place_91_rst, place_91_top, reset, clk);

  place_92 : place
  generic map(1, 1, '0')
  port map(place_92_tip, place_92_rst, place_92_top, reset, clk);

  place_93 : place
  generic map(1, 1, '0')
  port map(place_93_tip, place_93_rst, place_93_top, reset, clk);

  place_94 : place
  generic map(1, 1, '0')
  port map(place_94_tip, place_94_rst, place_94_top, reset, clk);

  place_95 : place
  generic map(1, 1, '0')
  port map(place_95_tip, place_95_rst, place_95_top, reset, clk);

  place_96 : place
  generic map(1, 1, '0')
  port map(place_96_tip, place_96_rst, place_96_top, reset, clk);

  place_97 : place
  generic map(1, 1, '0')
  port map(place_97_tip, place_97_rst, place_97_top, reset, clk);

  place_98 : place
  generic map(1, 1, '0')
  port map(place_98_tip, place_98_rst, place_98_top, reset, clk);

  place_99 : place
  generic map(1, 2, '0')
  port map(place_99_tip, place_99_rst, place_99_top, reset, clk);


  cbr_0_oper_tmp_d_35_bool_d_req : transition
  generic map(1)
  port map(cbr_0_oper_tmp_d_35_bool_d_req_tip, cbr_0_oper_tmp_d_35_bool_d_req_ge, cbr_0_oper_tmp_d_35_bool_d_req_top);

  cbr_1_oper_tmp_d_3_bool_d_req : transition
  generic map(2)
  port map(cbr_1_oper_tmp_d_3_bool_d_req_tip, cbr_1_oper_tmp_d_3_bool_d_req_ge, cbr_1_oper_tmp_d_3_bool_d_req_top);

  cbr_2_oper_tmp_d_11_bool_d_req : transition
  generic map(2)
  port map(cbr_2_oper_tmp_d_11_bool_d_req_tip, cbr_2_oper_tmp_d_11_bool_d_req_ge, cbr_2_oper_tmp_d_11_bool_d_req_top);

  cbr_3_oper_tmp_d_1114_bool_d_req : transition
  generic map(2)
  port map(cbr_3_oper_tmp_d_1114_bool_d_req_tip, cbr_3_oper_tmp_d_1114_bool_d_req_ge, cbr_3_oper_tmp_d_1114_bool_d_req_top);

  cbr_4_oper_tmp_d_2621_bool_d_req : transition
  generic map(2)
  port map(cbr_4_oper_tmp_d_2621_bool_d_req_tip, cbr_4_oper_tmp_d_2621_bool_d_req_ge, cbr_4_oper_tmp_d_2621_bool_d_req_top);

  cbr_5_oper_tmp_d_26_bool_d_req : transition
  generic map(2)
  port map(cbr_5_oper_tmp_d_26_bool_d_req_tip, cbr_5_oper_tmp_d_26_bool_d_req_ge, cbr_5_oper_tmp_d_26_bool_d_req_top);

  di_d_0_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(di_d_0_d_0_mux_1_d_ack_tip, di_d_0_d_0_mux_1_d_ack_ge, di_d_0_d_0_mux_1_d_ack_top);

  di_d_0_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(di_d_0_d_0_mux_1_d_req0_tip, di_d_0_d_0_mux_1_d_req0_ge, di_d_0_d_0_mux_1_d_req0_top);

  di_d_0_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(di_d_0_d_0_mux_1_d_req1_tip, di_d_0_d_0_mux_1_d_req1_ge, di_d_0_d_0_mux_1_d_req1_top);

  di_d_1_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(di_d_1_d_0_mux_1_d_ack_tip, di_d_1_d_0_mux_1_d_ack_ge, di_d_1_d_0_mux_1_d_ack_top);

  di_d_1_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(di_d_1_d_0_mux_1_d_req0_tip, di_d_1_d_0_mux_1_d_req0_ge, di_d_1_d_0_mux_1_d_req0_top);

  di_d_1_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(di_d_1_d_0_mux_1_d_req1_tip, di_d_1_d_0_mux_1_d_req1_ge, di_d_1_d_0_mux_1_d_req1_top);

  di_d_1_d_1_mux_1_d_ack : transition
  generic map(1)
  port map(di_d_1_d_1_mux_1_d_ack_tip, di_d_1_d_1_mux_1_d_ack_ge, di_d_1_d_1_mux_1_d_ack_top);

  di_d_1_d_1_mux_1_d_req0 : transition
  generic map(1)
  port map(di_d_1_d_1_mux_1_d_req0_tip, di_d_1_d_1_mux_1_d_req0_ge, di_d_1_d_1_mux_1_d_req0_top);

  di_d_1_d_1_mux_1_d_req1 : transition
  generic map(1)
  port map(di_d_1_d_1_mux_1_d_req1_tip, di_d_1_d_1_mux_1_d_req1_ge, di_d_1_d_1_mux_1_d_req1_top);

  di_d_1_mux_1_d_ack : transition
  generic map(1)
  port map(di_d_1_mux_1_d_ack_tip, di_d_1_mux_1_d_ack_ge, di_d_1_mux_1_d_ack_top);

  di_d_1_mux_1_d_req0 : transition
  generic map(1)
  port map(di_d_1_mux_1_d_req0_tip, di_d_1_mux_1_d_req0_ge, di_d_1_mux_1_d_req0_top);

  di_d_1_mux_1_d_req1 : transition
  generic map(1)
  port map(di_d_1_mux_1_d_req1_tip, di_d_1_mux_1_d_req1_ge, di_d_1_mux_1_d_req1_top);

  di_d_2_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(di_d_2_d_0_mux_1_d_ack_tip, di_d_2_d_0_mux_1_d_ack_ge, di_d_2_d_0_mux_1_d_ack_top);

  di_d_2_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(di_d_2_d_0_mux_1_d_req0_tip, di_d_2_d_0_mux_1_d_req0_ge, di_d_2_d_0_mux_1_d_req0_top);

  di_d_2_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(di_d_2_d_0_mux_1_d_req1_tip, di_d_2_d_0_mux_1_d_req1_ge, di_d_2_d_0_mux_1_d_req1_top);

  entry_to_loopentry_d_1_src : transition
  generic map(1)
  port map(entry_to_loopentry_d_1_src_tip, entry_to_loopentry_d_1_src_ge, entry_to_loopentry_d_1_src_top);

  entry_to_no_exit_d_0_d_preheader_src : transition
  generic map(1)
  port map(entry_to_no_exit_d_0_d_preheader_src_tip, entry_to_no_exit_d_0_d_preheader_src_ge, entry_to_no_exit_d_0_d_preheader_src_top);

  fin : transition
  generic map(1)
  port map(fin_tip, fin_ge, fin_top);

  init : transition
  generic map(1)
  port map(init_tip, init_ge, init_top);

  load_dividend_d_ack : transition
  generic map(1)
  port map(load_dividend_d_ack_tip, load_dividend_d_ack_ge, load_dividend_d_ack_top);

  load_dividend_d_req : transition
  generic map(1)
  port map(load_dividend_d_req_tip, load_dividend_d_req_ge, load_dividend_d_req_top);

  load_divisor_d_ack : transition
  generic map(1)
  port map(load_divisor_d_ack_tip, load_divisor_d_ack_ge, load_divisor_d_ack_top);

  load_divisor_d_req : transition
  generic map(1)
  port map(load_divisor_d_req_tip, load_divisor_d_req_ge, load_divisor_d_req_top);

  loopentry_d_1_d_entry : transition
  generic map(1)
  port map(loopentry_d_1_d_entry_tip, loopentry_d_1_d_entry_ge, loopentry_d_1_d_entry_top);

  loopentry_d_1_d_loopexit_to_loopentry_d_1_src : transition
  generic map(1)
  port map(loopentry_d_1_d_loopexit_to_loopentry_d_1_src_tip, loopentry_d_1_d_loopexit_to_loopentry_d_1_src_ge, loopentry_d_1_d_loopexit_to_loopentry_d_1_src_top);

  loopentry_d_1_d_pre : transition
  generic map(2)
  port map(loopentry_d_1_d_pre_tip, loopentry_d_1_d_pre_ge, loopentry_d_1_d_pre_top);

  loopentry_d_1_to_loopexit_d_1_src : transition
  generic map(1)
  port map(loopentry_d_1_to_loopexit_d_1_src_tip, loopentry_d_1_to_loopexit_d_1_src_ge, loopentry_d_1_to_loopexit_d_1_src_top);

  loopentry_d_1_to_no_exit_d_1_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_1_to_no_exit_d_1_d_preheader_src_tip, loopentry_d_1_to_no_exit_d_1_d_preheader_src_ge, loopentry_d_1_to_no_exit_d_1_d_preheader_src_top);

  loopexit_d_1_d_entry : transition
  generic map(1)
  port map(loopexit_d_1_d_entry_tip, loopexit_d_1_d_entry_ge, loopexit_d_1_d_entry_top);

  loopexit_d_1_d_loopexit_to_loopexit_d_1_src : transition
  generic map(1)
  port map(loopexit_d_1_d_loopexit_to_loopexit_d_1_src_tip, loopexit_d_1_d_loopexit_to_loopexit_d_1_src_ge, loopexit_d_1_d_loopexit_to_loopexit_d_1_src_top);

  loopexit_d_1_d_pre : transition
  generic map(2)
  port map(loopexit_d_1_d_pre_tip, loopexit_d_1_d_pre_ge, loopexit_d_1_d_pre_top);

  loopexit_d_1_to_loopexit_d_2_src : transition
  generic map(1)
  port map(loopexit_d_1_to_loopexit_d_2_src_tip, loopexit_d_1_to_loopexit_d_2_src_ge, loopexit_d_1_to_loopexit_d_2_src_top);

  loopexit_d_1_to_no_exit_d_2_d_preheader_src : transition
  generic map(1)
  port map(loopexit_d_1_to_no_exit_d_2_d_preheader_src_tip, loopexit_d_1_to_no_exit_d_2_d_preheader_src_ge, loopexit_d_1_to_no_exit_d_2_d_preheader_src_top);

  ni_d_0_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_0_d_0_mux_1_d_ack_tip, ni_d_0_d_0_mux_1_d_ack_ge, ni_d_0_d_0_mux_1_d_ack_top);

  ni_d_0_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_0_d_0_mux_1_d_req0_tip, ni_d_0_d_0_mux_1_d_req0_ge, ni_d_0_d_0_mux_1_d_req0_top);

  ni_d_0_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_0_d_0_mux_1_d_req1_tip, ni_d_0_d_0_mux_1_d_req1_ge, ni_d_0_d_0_mux_1_d_req1_top);

  ni_d_1_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_1_d_0_mux_1_d_ack_tip, ni_d_1_d_0_mux_1_d_ack_ge, ni_d_1_d_0_mux_1_d_ack_top);

  ni_d_1_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_1_d_0_mux_1_d_req0_tip, ni_d_1_d_0_mux_1_d_req0_ge, ni_d_1_d_0_mux_1_d_req0_top);

  ni_d_1_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_1_d_0_mux_1_d_req1_tip, ni_d_1_d_0_mux_1_d_req1_ge, ni_d_1_d_0_mux_1_d_req1_top);

  ni_d_1_d_1_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_1_d_1_mux_1_d_ack_tip, ni_d_1_d_1_mux_1_d_ack_ge, ni_d_1_d_1_mux_1_d_ack_top);

  ni_d_1_d_1_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_1_d_1_mux_1_d_req0_tip, ni_d_1_d_1_mux_1_d_req0_ge, ni_d_1_d_1_mux_1_d_req0_top);

  ni_d_1_d_1_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_1_d_1_mux_1_d_req1_tip, ni_d_1_d_1_mux_1_d_req1_ge, ni_d_1_d_1_mux_1_d_req1_top);

  ni_d_1_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_1_mux_1_d_ack_tip, ni_d_1_mux_1_d_ack_ge, ni_d_1_mux_1_d_ack_top);

  ni_d_1_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_1_mux_1_d_req0_tip, ni_d_1_mux_1_d_req0_ge, ni_d_1_mux_1_d_req0_top);

  ni_d_1_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_1_mux_1_d_req1_tip, ni_d_1_mux_1_d_req1_ge, ni_d_1_mux_1_d_req1_top);

  ni_d_2_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_2_d_0_mux_1_d_ack_tip, ni_d_2_d_0_mux_1_d_ack_ge, ni_d_2_d_0_mux_1_d_ack_top);

  ni_d_2_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_2_d_0_mux_1_d_req0_tip, ni_d_2_d_0_mux_1_d_req0_ge, ni_d_2_d_0_mux_1_d_req0_top);

  ni_d_2_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_2_d_0_mux_1_d_req1_tip, ni_d_2_d_0_mux_1_d_req1_ge, ni_d_2_d_0_mux_1_d_req1_top);

  ni_d_2_d_1_mux_1_d_ack : transition
  generic map(1)
  port map(ni_d_2_d_1_mux_1_d_ack_tip, ni_d_2_d_1_mux_1_d_ack_ge, ni_d_2_d_1_mux_1_d_ack_top);

  ni_d_2_d_1_mux_1_d_req0 : transition
  generic map(1)
  port map(ni_d_2_d_1_mux_1_d_req0_tip, ni_d_2_d_1_mux_1_d_req0_ge, ni_d_2_d_1_mux_1_d_req0_top);

  ni_d_2_d_1_mux_1_d_req1 : transition
  generic map(1)
  port map(ni_d_2_d_1_mux_1_d_req1_tip, ni_d_2_d_1_mux_1_d_req1_ge, ni_d_2_d_1_mux_1_d_req1_top);

  no_exit_d_0_d_entry : transition
  generic map(1)
  port map(no_exit_d_0_d_entry_tip, no_exit_d_0_d_entry_ge, no_exit_d_0_d_entry_top);

  no_exit_d_0_d_pre : transition
  generic map(2)
  port map(no_exit_d_0_d_pre_tip, no_exit_d_0_d_pre_ge, no_exit_d_0_d_pre_top);

  no_exit_d_0_d_preheader_to_no_exit_d_0_src : transition
  generic map(1)
  port map(no_exit_d_0_d_preheader_to_no_exit_d_0_src_tip, no_exit_d_0_d_preheader_to_no_exit_d_0_src_ge, no_exit_d_0_d_preheader_to_no_exit_d_0_src_top);

  no_exit_d_0_to_loopentry_d_1_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_0_to_loopentry_d_1_d_loopexit_src_tip, no_exit_d_0_to_loopentry_d_1_d_loopexit_src_ge, no_exit_d_0_to_loopentry_d_1_d_loopexit_src_top);

  no_exit_d_0_to_no_exit_d_0_src : transition
  generic map(1)
  port map(no_exit_d_0_to_no_exit_d_0_src_tip, no_exit_d_0_to_no_exit_d_0_src_ge, no_exit_d_0_to_no_exit_d_0_src_top);

  no_exit_d_1_d_entry : transition
  generic map(1)
  port map(no_exit_d_1_d_entry_tip, no_exit_d_1_d_entry_ge, no_exit_d_1_d_entry_top);

  no_exit_d_1_d_pre : transition
  generic map(2)
  port map(no_exit_d_1_d_pre_tip, no_exit_d_1_d_pre_ge, no_exit_d_1_d_pre_top);

  no_exit_d_1_d_preheader_to_no_exit_d_1_src : transition
  generic map(1)
  port map(no_exit_d_1_d_preheader_to_no_exit_d_1_src_tip, no_exit_d_1_d_preheader_to_no_exit_d_1_src_ge, no_exit_d_1_d_preheader_to_no_exit_d_1_src_top);

  no_exit_d_1_to_loopexit_d_1_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_1_to_loopexit_d_1_d_loopexit_src_tip, no_exit_d_1_to_loopexit_d_1_d_loopexit_src_ge, no_exit_d_1_to_loopexit_d_1_d_loopexit_src_top);

  no_exit_d_1_to_no_exit_d_1_src : transition
  generic map(1)
  port map(no_exit_d_1_to_no_exit_d_1_src_tip, no_exit_d_1_to_no_exit_d_1_src_ge, no_exit_d_1_to_no_exit_d_1_src_top);

  no_exit_d_2_d_entry : transition
  generic map(1)
  port map(no_exit_d_2_d_entry_tip, no_exit_d_2_d_entry_ge, no_exit_d_2_d_entry_top);

  no_exit_d_2_d_pre : transition
  generic map(3)
  port map(no_exit_d_2_d_pre_tip, no_exit_d_2_d_pre_ge, no_exit_d_2_d_pre_top);

  no_exit_d_2_d_preheader_to_no_exit_d_2_src : transition
  generic map(1)
  port map(no_exit_d_2_d_preheader_to_no_exit_d_2_src_tip, no_exit_d_2_d_preheader_to_no_exit_d_2_src_ge, no_exit_d_2_d_preheader_to_no_exit_d_2_src_top);

  no_exit_d_2_to_loopexit_d_2_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_2_to_loopexit_d_2_d_loopexit_src_tip, no_exit_d_2_to_loopexit_d_2_d_loopexit_src_ge, no_exit_d_2_to_loopexit_d_2_d_loopexit_src_top);

  no_exit_d_2_to_no_exit_d_2_src : transition
  generic map(1)
  port map(no_exit_d_2_to_no_exit_d_2_src_tip, no_exit_d_2_to_no_exit_d_2_src_ge, no_exit_d_2_to_no_exit_d_2_src_top);

  oper_tmp_d_1114_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_1114_bool_d_ack_tip, oper_tmp_d_1114_bool_d_ack_ge, oper_tmp_d_1114_bool_d_ack_top);

  oper_tmp_d_1114_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_1114_bool_d_req_tip, oper_tmp_d_1114_bool_d_req_ge, oper_tmp_d_1114_bool_d_req_top);

  oper_tmp_d_11_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11_bool_d_ack_tip, oper_tmp_d_11_bool_d_ack_ge, oper_tmp_d_11_bool_d_ack_top);

  oper_tmp_d_11_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11_bool_d_req_tip, oper_tmp_d_11_bool_d_req_ge, oper_tmp_d_11_bool_d_req_top);

  oper_tmp_d_14_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_14_float_d_ack_tip, oper_tmp_d_14_float_d_ack_ge, oper_tmp_d_14_float_d_ack_top);

  oper_tmp_d_14_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_14_float_d_req_tip, oper_tmp_d_14_float_d_req_ge, oper_tmp_d_14_float_d_req_top);

  oper_tmp_d_16_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_16_float_d_ack_tip, oper_tmp_d_16_float_d_ack_ge, oper_tmp_d_16_float_d_ack_top);

  oper_tmp_d_16_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_16_float_d_req_tip, oper_tmp_d_16_float_d_req_ge, oper_tmp_d_16_float_d_req_top);

  oper_tmp_d_19_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_19_float_d_ack_tip, oper_tmp_d_19_float_d_ack_ge, oper_tmp_d_19_float_d_ack_top);

  oper_tmp_d_19_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_19_float_d_req_tip, oper_tmp_d_19_float_d_req_ge, oper_tmp_d_19_float_d_req_top);

  oper_tmp_d_21_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_21_float_d_ack_tip, oper_tmp_d_21_float_d_ack_ge, oper_tmp_d_21_float_d_ack_top);

  oper_tmp_d_21_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_21_float_d_req_tip, oper_tmp_d_21_float_d_req_ge, oper_tmp_d_21_float_d_req_top);

  oper_tmp_d_2420_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_2420_float_d_ack_tip, oper_tmp_d_2420_float_d_ack_ge, oper_tmp_d_2420_float_d_ack_top);

  oper_tmp_d_2420_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_2420_float_d_req_tip, oper_tmp_d_2420_float_d_req_ge, oper_tmp_d_2420_float_d_req_top);

  oper_tmp_d_24_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_24_float_d_ack_tip, oper_tmp_d_24_float_d_ack_ge, oper_tmp_d_24_float_d_ack_top);

  oper_tmp_d_24_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_24_float_d_req_tip, oper_tmp_d_24_float_d_req_ge, oper_tmp_d_24_float_d_req_top);

  oper_tmp_d_2621_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_2621_bool_d_ack_tip, oper_tmp_d_2621_bool_d_ack_ge, oper_tmp_d_2621_bool_d_ack_top);

  oper_tmp_d_2621_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_2621_bool_d_req_tip, oper_tmp_d_2621_bool_d_req_ge, oper_tmp_d_2621_bool_d_req_top);

  oper_tmp_d_26_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_26_bool_d_ack_tip, oper_tmp_d_26_bool_d_ack_ge, oper_tmp_d_26_bool_d_ack_top);

  oper_tmp_d_26_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_26_bool_d_req_tip, oper_tmp_d_26_bool_d_req_ge, oper_tmp_d_26_bool_d_req_top);

  oper_tmp_d_31_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_31_float_d_ack_tip, oper_tmp_d_31_float_d_ack_ge, oper_tmp_d_31_float_d_ack_top);

  oper_tmp_d_31_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_31_float_d_req_tip, oper_tmp_d_31_float_d_req_ge, oper_tmp_d_31_float_d_req_top);

  oper_tmp_d_34_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_34_float_d_ack_tip, oper_tmp_d_34_float_d_ack_ge, oper_tmp_d_34_float_d_ack_top);

  oper_tmp_d_34_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_34_float_d_req_tip, oper_tmp_d_34_float_d_req_ge, oper_tmp_d_34_float_d_req_top);

  oper_tmp_d_35_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_35_bool_d_ack_tip, oper_tmp_d_35_bool_d_ack_ge, oper_tmp_d_35_bool_d_ack_top);

  oper_tmp_d_35_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_35_bool_d_req_tip, oper_tmp_d_35_bool_d_req_ge, oper_tmp_d_35_bool_d_req_top);

  oper_tmp_d_36_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_36_float_d_ack_tip, oper_tmp_d_36_float_d_ack_ge, oper_tmp_d_36_float_d_ack_top);

  oper_tmp_d_36_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_36_float_d_req_tip, oper_tmp_d_36_float_d_req_ge, oper_tmp_d_36_float_d_req_top);

  oper_tmp_d_3_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_3_bool_d_ack_tip, oper_tmp_d_3_bool_d_ack_ge, oper_tmp_d_3_bool_d_ack_top);

  oper_tmp_d_3_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_3_bool_d_req_tip, oper_tmp_d_3_bool_d_req_ge, oper_tmp_d_3_bool_d_req_top);

  oper_tmp_d_6_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_6_float_d_ack_tip, oper_tmp_d_6_float_d_ack_ge, oper_tmp_d_6_float_d_ack_top);

  oper_tmp_d_6_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_6_float_d_req_tip, oper_tmp_d_6_float_d_req_ge, oper_tmp_d_6_float_d_req_top);

  oper_tmp_d_8_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_8_float_d_ack_tip, oper_tmp_d_8_float_d_ack_ge, oper_tmp_d_8_float_d_ack_top);

  oper_tmp_d_8_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_8_float_d_req_tip, oper_tmp_d_8_float_d_req_ge, oper_tmp_d_8_float_d_req_top);

  ri_d_0_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(ri_d_0_d_0_mux_1_d_ack_tip, ri_d_0_d_0_mux_1_d_ack_ge, ri_d_0_d_0_mux_1_d_ack_top);

  ri_d_0_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(ri_d_0_d_0_mux_1_d_req0_tip, ri_d_0_d_0_mux_1_d_req0_ge, ri_d_0_d_0_mux_1_d_req0_top);

  ri_d_0_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(ri_d_0_d_0_mux_1_d_req1_tip, ri_d_0_d_0_mux_1_d_req1_ge, ri_d_0_d_0_mux_1_d_req1_top);

  store_location_divide_return_d_ack : transition
  generic map(1)
  port map(store_location_divide_return_d_ack_tip, store_location_divide_return_d_ack_ge, store_location_divide_return_d_ack_top);

  store_location_divide_return_d_req : transition
  generic map(1)
  port map(store_location_divide_return_d_req_tip, store_location_divide_return_d_req_ge, store_location_divide_return_d_req_top);

  place_1_tip(0) <= load_divisor_d_ack_top;
  place_1_rst(0) <= oper_tmp_d_35_bool_d_req_top;
  place_10_tip(0) <= loopexit_d_1_d_pre_top;
  place_10_rst(0) <= loopexit_d_1_d_entry_top;
  place_101_tip(0) <= no_exit_d_2_d_preheader_to_no_exit_d_2_src_top;
  place_101_rst(0) <= di_d_2_d_0_mux_1_d_req1_top;
  place_102_tip(0) <= di_d_2_d_0_mux_1_d_req0_top;
  place_102_tip(1) <= di_d_2_d_0_mux_1_d_req1_top;
  place_102_rst(0) <= di_d_2_d_0_mux_1_d_ack_top;
  place_103_tip(0) <= di_d_2_d_0_mux_1_d_ack_top;
  place_103_rst(0) <= no_exit_d_2_d_pre_top;
  place_104_tip(0) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_104_rst(0) <= di_d_2_d_0_mux_1_d_req0_top;
  place_105_tip(0) <= no_exit_d_2_d_preheader_to_no_exit_d_2_src_top;
  place_105_rst(0) <= ni_d_2_d_0_mux_1_d_req1_top;
  place_106_tip(0) <= ni_d_2_d_0_mux_1_d_req0_top;
  place_106_tip(1) <= ni_d_2_d_0_mux_1_d_req1_top;
  place_106_rst(0) <= ni_d_2_d_0_mux_1_d_ack_top;
  place_107_tip(0) <= ni_d_2_d_0_mux_1_d_ack_top;
  place_107_rst(0) <= no_exit_d_2_d_pre_top;
  place_108_tip(0) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_108_rst(0) <= ni_d_2_d_0_mux_1_d_req0_top;
  place_109_tip(0) <= no_exit_d_2_d_preheader_to_no_exit_d_2_src_top;
  place_109_rst(0) <= ri_d_0_d_0_mux_1_d_req1_top;
  place_11_tip(0) <= no_exit_d_1_d_pre_top;
  place_11_rst(0) <= no_exit_d_1_d_entry_top;
  place_110_tip(0) <= ri_d_0_d_0_mux_1_d_req0_top;
  place_110_tip(1) <= ri_d_0_d_0_mux_1_d_req1_top;
  place_110_rst(0) <= ri_d_0_d_0_mux_1_d_ack_top;
  place_111_tip(0) <= ri_d_0_d_0_mux_1_d_ack_top;
  place_111_rst(0) <= no_exit_d_2_d_pre_top;
  place_112_tip(0) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_112_rst(0) <= ri_d_0_d_0_mux_1_d_req0_top;
  place_113_tip(0) <= oper_tmp_d_31_float_d_req_top;
  place_113_rst(0) <= oper_tmp_d_31_float_d_ack_top;
  place_114_tip(0) <= no_exit_d_2_d_entry_top;
  place_114_rst(0) <= oper_tmp_d_31_float_d_req_top;
  place_115_tip(0) <= oper_tmp_d_34_float_d_req_top;
  place_115_rst(0) <= oper_tmp_d_34_float_d_ack_top;
  place_116_tip(0) <= no_exit_d_2_d_entry_top;
  place_116_rst(0) <= oper_tmp_d_34_float_d_req_top;
  place_117_tip(0) <= oper_tmp_d_36_float_d_req_top;
  place_117_rst(0) <= oper_tmp_d_36_float_d_ack_top;
  place_118_tip(0) <= oper_tmp_d_31_float_d_ack_top;
  place_118_rst(0) <= oper_tmp_d_36_float_d_req_top;
  place_119_tip(0) <= oper_tmp_d_36_float_d_ack_top;
  place_119_rst(0) <= cbr_5_oper_tmp_d_26_bool_d_req_top;
  place_120_tip(0) <= oper_tmp_d_24_float_d_req_top;
  place_120_rst(0) <= oper_tmp_d_24_float_d_ack_top;
  place_121_tip(0) <= oper_tmp_d_34_float_d_ack_top;
  place_121_rst(0) <= oper_tmp_d_24_float_d_req_top;
  place_122_tip(0) <= oper_tmp_d_26_bool_d_req_top;
  place_122_rst(0) <= oper_tmp_d_26_bool_d_ack_top;
  place_123_tip(0) <= oper_tmp_d_24_float_d_ack_top;
  place_123_rst(0) <= oper_tmp_d_26_bool_d_req_top;
  place_124_tip(0) <= oper_tmp_d_26_bool_d_ack_top;
  place_124_rst(0) <= cbr_5_oper_tmp_d_26_bool_d_req_top;
  place_125_tip(0) <= cbr_5_oper_tmp_d_26_bool_d_req_top;
  place_125_rst(0) <= no_exit_d_2_to_loopexit_d_2_d_loopexit_src_top;
  place_125_rst(1) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_128_tip(0) <= ni_d_2_d_1_mux_1_d_req0_top;
  place_128_tip(1) <= ni_d_2_d_1_mux_1_d_req1_top;
  place_128_rst(0) <= ni_d_2_d_1_mux_1_d_ack_top;
  place_129_tip(0) <= ni_d_2_d_1_mux_1_d_ack_top;
  place_129_rst(0) <= store_location_divide_return_d_req_top;
  place_13_tip(0) <= no_exit_d_1_to_loopexit_d_1_d_loopexit_src_top;
  place_13_rst(0) <= loopexit_d_1_d_loopexit_to_loopexit_d_1_src_top;
  place_130_tip(0) <= loopexit_d_1_to_loopexit_d_2_src_top;
  place_130_rst(0) <= ni_d_2_d_1_mux_1_d_req0_top;
  place_131_tip(0) <= store_location_divide_return_d_req_top;
  place_131_rst(0) <= store_location_divide_return_d_ack_top;
  place_15_tip(0) <= loopexit_d_1_to_no_exit_d_2_d_preheader_src_top;
  place_15_rst(0) <= no_exit_d_2_d_preheader_to_no_exit_d_2_src_top;
  place_17_tip(0) <= no_exit_d_2_d_pre_top;
  place_17_rst(0) <= no_exit_d_2_d_entry_top;
  place_19_tip(0) <= no_exit_d_2_to_loopexit_d_2_d_loopexit_src_top;
  place_19_rst(0) <= ni_d_2_d_1_mux_1_d_req1_top;
  place_2_tip(0) <= loopentry_d_1_d_pre_top;
  place_2_rst(0) <= loopentry_d_1_d_entry_top;
  place_20_tip(0) <= fin_top;
  place_20_rst(0) <= init_top;
  place_21_tip(0) <= store_location_divide_return_d_ack_top;
  place_21_rst(0) <= fin_top;
  place_22_tip(0) <= init_top;
  place_22_rst(0) <= load_dividend_d_req_top;
  place_23_tip(0) <= load_dividend_d_req_top;
  place_23_rst(0) <= load_dividend_d_ack_top;
  place_24_tip(0) <= load_dividend_d_ack_top;
  place_24_rst(0) <= load_divisor_d_req_top;
  place_25_tip(0) <= load_divisor_d_req_top;
  place_25_rst(0) <= load_divisor_d_ack_top;
  place_26_tip(0) <= oper_tmp_d_35_bool_d_req_top;
  place_26_rst(0) <= oper_tmp_d_35_bool_d_ack_top;
  place_28_tip(0) <= oper_tmp_d_35_bool_d_ack_top;
  place_28_rst(0) <= cbr_0_oper_tmp_d_35_bool_d_req_top;
  place_29_tip(0) <= cbr_0_oper_tmp_d_35_bool_d_req_top;
  place_29_rst(0) <= entry_to_loopentry_d_1_src_top;
  place_29_rst(1) <= entry_to_no_exit_d_0_d_preheader_src_top;
  place_31_tip(0) <= no_exit_d_0_d_preheader_to_no_exit_d_0_src_top;
  place_31_rst(0) <= di_d_0_d_0_mux_1_d_req1_top;
  place_32_tip(0) <= di_d_0_d_0_mux_1_d_req0_top;
  place_32_tip(1) <= di_d_0_d_0_mux_1_d_req1_top;
  place_32_rst(0) <= di_d_0_d_0_mux_1_d_ack_top;
  place_33_tip(0) <= di_d_0_d_0_mux_1_d_ack_top;
  place_33_rst(0) <= no_exit_d_0_d_pre_top;
  place_34_tip(0) <= no_exit_d_0_to_no_exit_d_0_src_top;
  place_34_rst(0) <= di_d_0_d_0_mux_1_d_req0_top;
  place_35_tip(0) <= no_exit_d_0_d_preheader_to_no_exit_d_0_src_top;
  place_35_rst(0) <= ni_d_0_d_0_mux_1_d_req1_top;
  place_36_tip(0) <= ni_d_0_d_0_mux_1_d_req0_top;
  place_36_tip(1) <= ni_d_0_d_0_mux_1_d_req1_top;
  place_36_rst(0) <= ni_d_0_d_0_mux_1_d_ack_top;
  place_37_tip(0) <= ni_d_0_d_0_mux_1_d_ack_top;
  place_37_rst(0) <= no_exit_d_0_d_pre_top;
  place_38_tip(0) <= no_exit_d_0_to_no_exit_d_0_src_top;
  place_38_rst(0) <= ni_d_0_d_0_mux_1_d_req0_top;
  place_39_tip(0) <= oper_tmp_d_6_float_d_req_top;
  place_39_rst(0) <= oper_tmp_d_6_float_d_ack_top;
  place_4_tip(0) <= entry_to_no_exit_d_0_d_preheader_src_top;
  place_4_rst(0) <= no_exit_d_0_d_preheader_to_no_exit_d_0_src_top;
  place_40_tip(0) <= no_exit_d_0_d_entry_top;
  place_40_rst(0) <= oper_tmp_d_6_float_d_req_top;
  place_41_tip(0) <= oper_tmp_d_8_float_d_req_top;
  place_41_rst(0) <= oper_tmp_d_8_float_d_ack_top;
  place_42_tip(0) <= no_exit_d_0_d_entry_top;
  place_42_rst(0) <= oper_tmp_d_8_float_d_req_top;
  place_43_tip(0) <= oper_tmp_d_8_float_d_ack_top;
  place_43_rst(0) <= cbr_1_oper_tmp_d_3_bool_d_req_top;
  place_44_tip(0) <= oper_tmp_d_3_bool_d_req_top;
  place_44_rst(0) <= oper_tmp_d_3_bool_d_ack_top;
  place_45_tip(0) <= oper_tmp_d_6_float_d_ack_top;
  place_45_rst(0) <= oper_tmp_d_3_bool_d_req_top;
  place_46_tip(0) <= oper_tmp_d_3_bool_d_ack_top;
  place_46_rst(0) <= cbr_1_oper_tmp_d_3_bool_d_req_top;
  place_47_tip(0) <= cbr_1_oper_tmp_d_3_bool_d_req_top;
  place_47_rst(0) <= no_exit_d_0_to_loopentry_d_1_d_loopexit_src_top;
  place_47_rst(1) <= no_exit_d_0_to_no_exit_d_0_src_top;
  place_49_tip(0) <= loopentry_d_1_d_loopexit_to_loopentry_d_1_src_top;
  place_49_rst(0) <= di_d_1_mux_1_d_req1_top;
  place_5_tip(0) <= no_exit_d_0_d_pre_top;
  place_5_rst(0) <= no_exit_d_0_d_entry_top;
  place_50_tip(0) <= di_d_1_mux_1_d_req0_top;
  place_50_tip(1) <= di_d_1_mux_1_d_req1_top;
  place_50_rst(0) <= di_d_1_mux_1_d_ack_top;
  place_51_tip(0) <= di_d_1_mux_1_d_ack_top;
  place_51_rst(0) <= loopentry_d_1_d_pre_top;
  place_52_tip(0) <= entry_to_loopentry_d_1_src_top;
  place_52_rst(0) <= di_d_1_mux_1_d_req0_top;
  place_53_tip(0) <= loopentry_d_1_d_loopexit_to_loopentry_d_1_src_top;
  place_53_rst(0) <= ni_d_1_mux_1_d_req1_top;
  place_54_tip(0) <= ni_d_1_mux_1_d_req0_top;
  place_54_tip(1) <= ni_d_1_mux_1_d_req1_top;
  place_54_rst(0) <= ni_d_1_mux_1_d_ack_top;
  place_55_tip(0) <= ni_d_1_mux_1_d_ack_top;
  place_55_rst(0) <= loopentry_d_1_d_pre_top;
  place_56_tip(0) <= entry_to_loopentry_d_1_src_top;
  place_56_rst(0) <= ni_d_1_mux_1_d_req0_top;
  place_57_tip(0) <= loopentry_d_1_d_entry_top;
  place_57_rst(0) <= cbr_2_oper_tmp_d_11_bool_d_req_top;
  place_58_tip(0) <= oper_tmp_d_11_bool_d_req_top;
  place_58_rst(0) <= oper_tmp_d_11_bool_d_ack_top;
  place_59_tip(0) <= loopentry_d_1_d_entry_top;
  place_59_rst(0) <= oper_tmp_d_11_bool_d_req_top;
  place_60_tip(0) <= oper_tmp_d_11_bool_d_ack_top;
  place_60_rst(0) <= cbr_2_oper_tmp_d_11_bool_d_req_top;
  place_61_tip(0) <= cbr_2_oper_tmp_d_11_bool_d_req_top;
  place_61_rst(0) <= loopentry_d_1_to_loopexit_d_1_src_top;
  place_61_rst(1) <= loopentry_d_1_to_no_exit_d_1_d_preheader_src_top;
  place_63_tip(0) <= no_exit_d_1_d_preheader_to_no_exit_d_1_src_top;
  place_63_rst(0) <= di_d_1_d_0_mux_1_d_req1_top;
  place_64_tip(0) <= di_d_1_d_0_mux_1_d_req0_top;
  place_64_tip(1) <= di_d_1_d_0_mux_1_d_req1_top;
  place_64_rst(0) <= di_d_1_d_0_mux_1_d_ack_top;
  place_65_tip(0) <= di_d_1_d_0_mux_1_d_ack_top;
  place_65_rst(0) <= no_exit_d_1_d_pre_top;
  place_66_tip(0) <= no_exit_d_1_to_no_exit_d_1_src_top;
  place_66_rst(0) <= di_d_1_d_0_mux_1_d_req0_top;
  place_67_tip(0) <= no_exit_d_1_d_preheader_to_no_exit_d_1_src_top;
  place_67_rst(0) <= ni_d_1_d_0_mux_1_d_req1_top;
  place_68_tip(0) <= ni_d_1_d_0_mux_1_d_req0_top;
  place_68_tip(1) <= ni_d_1_d_0_mux_1_d_req1_top;
  place_68_rst(0) <= ni_d_1_d_0_mux_1_d_ack_top;
  place_69_tip(0) <= ni_d_1_d_0_mux_1_d_ack_top;
  place_69_rst(0) <= no_exit_d_1_d_pre_top;
  place_7_tip(0) <= no_exit_d_0_to_loopentry_d_1_d_loopexit_src_top;
  place_7_rst(0) <= loopentry_d_1_d_loopexit_to_loopentry_d_1_src_top;
  place_70_tip(0) <= no_exit_d_1_to_no_exit_d_1_src_top;
  place_70_rst(0) <= ni_d_1_d_0_mux_1_d_req0_top;
  place_71_tip(0) <= oper_tmp_d_14_float_d_req_top;
  place_71_rst(0) <= oper_tmp_d_14_float_d_ack_top;
  place_72_tip(0) <= no_exit_d_1_d_entry_top;
  place_72_rst(0) <= oper_tmp_d_14_float_d_req_top;
  place_73_tip(0) <= oper_tmp_d_16_float_d_req_top;
  place_73_rst(0) <= oper_tmp_d_16_float_d_ack_top;
  place_74_tip(0) <= no_exit_d_1_d_entry_top;
  place_74_rst(0) <= oper_tmp_d_16_float_d_req_top;
  place_75_tip(0) <= oper_tmp_d_16_float_d_ack_top;
  place_75_rst(0) <= cbr_3_oper_tmp_d_1114_bool_d_req_top;
  place_76_tip(0) <= oper_tmp_d_1114_bool_d_req_top;
  place_76_rst(0) <= oper_tmp_d_1114_bool_d_ack_top;
  place_77_tip(0) <= oper_tmp_d_14_float_d_ack_top;
  place_77_rst(0) <= oper_tmp_d_1114_bool_d_req_top;
  place_78_tip(0) <= oper_tmp_d_1114_bool_d_ack_top;
  place_78_rst(0) <= cbr_3_oper_tmp_d_1114_bool_d_req_top;
  place_79_tip(0) <= cbr_3_oper_tmp_d_1114_bool_d_req_top;
  place_79_rst(0) <= no_exit_d_1_to_loopexit_d_1_d_loopexit_src_top;
  place_79_rst(1) <= no_exit_d_1_to_no_exit_d_1_src_top;
  place_81_tip(0) <= loopexit_d_1_d_loopexit_to_loopexit_d_1_src_top;
  place_81_rst(0) <= di_d_1_d_1_mux_1_d_req1_top;
  place_82_tip(0) <= di_d_1_d_1_mux_1_d_req0_top;
  place_82_tip(1) <= di_d_1_d_1_mux_1_d_req1_top;
  place_82_rst(0) <= di_d_1_d_1_mux_1_d_ack_top;
  place_83_tip(0) <= di_d_1_d_1_mux_1_d_ack_top;
  place_83_rst(0) <= loopexit_d_1_d_pre_top;
  place_84_tip(0) <= loopentry_d_1_to_loopexit_d_1_src_top;
  place_84_rst(0) <= di_d_1_d_1_mux_1_d_req0_top;
  place_85_tip(0) <= loopexit_d_1_d_loopexit_to_loopexit_d_1_src_top;
  place_85_rst(0) <= ni_d_1_d_1_mux_1_d_req1_top;
  place_86_tip(0) <= ni_d_1_d_1_mux_1_d_req0_top;
  place_86_tip(1) <= ni_d_1_d_1_mux_1_d_req1_top;
  place_86_rst(0) <= ni_d_1_d_1_mux_1_d_ack_top;
  place_87_tip(0) <= ni_d_1_d_1_mux_1_d_ack_top;
  place_87_rst(0) <= loopexit_d_1_d_pre_top;
  place_88_tip(0) <= loopentry_d_1_to_loopexit_d_1_src_top;
  place_88_rst(0) <= ni_d_1_d_1_mux_1_d_req0_top;
  place_89_tip(0) <= oper_tmp_d_19_float_d_req_top;
  place_89_rst(0) <= oper_tmp_d_19_float_d_ack_top;
  place_9_tip(0) <= loopentry_d_1_to_no_exit_d_1_d_preheader_src_top;
  place_9_rst(0) <= no_exit_d_1_d_preheader_to_no_exit_d_1_src_top;
  place_90_tip(0) <= loopexit_d_1_d_entry_top;
  place_90_rst(0) <= oper_tmp_d_19_float_d_req_top;
  place_91_tip(0) <= oper_tmp_d_21_float_d_req_top;
  place_91_rst(0) <= oper_tmp_d_21_float_d_ack_top;
  place_92_tip(0) <= loopexit_d_1_d_entry_top;
  place_92_rst(0) <= oper_tmp_d_21_float_d_req_top;
  place_93_tip(0) <= oper_tmp_d_21_float_d_ack_top;
  place_93_rst(0) <= cbr_4_oper_tmp_d_2621_bool_d_req_top;
  place_94_tip(0) <= oper_tmp_d_2420_float_d_req_top;
  place_94_rst(0) <= oper_tmp_d_2420_float_d_ack_top;
  place_95_tip(0) <= oper_tmp_d_19_float_d_ack_top;
  place_95_rst(0) <= oper_tmp_d_2420_float_d_req_top;
  place_96_tip(0) <= oper_tmp_d_2621_bool_d_req_top;
  place_96_rst(0) <= oper_tmp_d_2621_bool_d_ack_top;
  place_97_tip(0) <= oper_tmp_d_2420_float_d_ack_top;
  place_97_rst(0) <= oper_tmp_d_2621_bool_d_req_top;
  place_98_tip(0) <= oper_tmp_d_2621_bool_d_ack_top;
  place_98_rst(0) <= cbr_4_oper_tmp_d_2621_bool_d_req_top;
  place_99_tip(0) <= cbr_4_oper_tmp_d_2621_bool_d_req_top;
  place_99_rst(0) <= loopexit_d_1_to_loopexit_d_2_src_top;
  place_99_rst(1) <= loopexit_d_1_to_no_exit_d_2_d_preheader_src_top;

  cbr_0_oper_tmp_d_35_bool_d_req_tip(0) <= place_28_top;
  cbr_1_oper_tmp_d_3_bool_d_req_tip(0) <= place_43_top;
  cbr_1_oper_tmp_d_3_bool_d_req_tip(1) <= place_46_top;
  cbr_2_oper_tmp_d_11_bool_d_req_tip(0) <= place_57_top;
  cbr_2_oper_tmp_d_11_bool_d_req_tip(1) <= place_60_top;
  cbr_3_oper_tmp_d_1114_bool_d_req_tip(0) <= place_75_top;
  cbr_3_oper_tmp_d_1114_bool_d_req_tip(1) <= place_78_top;
  cbr_4_oper_tmp_d_2621_bool_d_req_tip(0) <= place_93_top;
  cbr_4_oper_tmp_d_2621_bool_d_req_tip(1) <= place_98_top;
  cbr_5_oper_tmp_d_26_bool_d_req_tip(0) <= place_119_top;
  cbr_5_oper_tmp_d_26_bool_d_req_tip(1) <= place_124_top;
  di_d_0_d_0_mux_1_d_ack_tip(0) <= place_32_top;
  di_d_0_d_0_mux_1_d_req0_tip(0) <= place_34_top;
  di_d_0_d_0_mux_1_d_req1_tip(0) <= place_31_top;
  di_d_1_d_0_mux_1_d_ack_tip(0) <= place_64_top;
  di_d_1_d_0_mux_1_d_req0_tip(0) <= place_66_top;
  di_d_1_d_0_mux_1_d_req1_tip(0) <= place_63_top;
  di_d_1_d_1_mux_1_d_ack_tip(0) <= place_82_top;
  di_d_1_d_1_mux_1_d_req0_tip(0) <= place_84_top;
  di_d_1_d_1_mux_1_d_req1_tip(0) <= place_81_top;
  di_d_1_mux_1_d_ack_tip(0) <= place_50_top;
  di_d_1_mux_1_d_req0_tip(0) <= place_52_top;
  di_d_1_mux_1_d_req1_tip(0) <= place_49_top;
  di_d_2_d_0_mux_1_d_ack_tip(0) <= place_102_top;
  di_d_2_d_0_mux_1_d_req0_tip(0) <= place_104_top;
  di_d_2_d_0_mux_1_d_req1_tip(0) <= place_101_top;
  entry_to_loopentry_d_1_src_tip(0) <= place_29_top;
  entry_to_no_exit_d_0_d_preheader_src_tip(0) <= place_29_top;
  fin_tip(0) <= place_21_top;
  init_tip(0) <= place_20_top;
  load_dividend_d_ack_tip(0) <= place_23_top;
  load_dividend_d_req_tip(0) <= place_22_top;
  load_divisor_d_ack_tip(0) <= place_25_top;
  load_divisor_d_req_tip(0) <= place_24_top;
  loopentry_d_1_d_entry_tip(0) <= place_2_top;
  loopentry_d_1_d_loopexit_to_loopentry_d_1_src_tip(0) <= place_7_top;
  loopentry_d_1_d_pre_tip(0) <= place_51_top;
  loopentry_d_1_d_pre_tip(1) <= place_55_top;
  loopentry_d_1_to_loopexit_d_1_src_tip(0) <= place_61_top;
  loopentry_d_1_to_no_exit_d_1_d_preheader_src_tip(0) <= place_61_top;
  loopexit_d_1_d_entry_tip(0) <= place_10_top;
  loopexit_d_1_d_loopexit_to_loopexit_d_1_src_tip(0) <= place_13_top;
  loopexit_d_1_d_pre_tip(0) <= place_83_top;
  loopexit_d_1_d_pre_tip(1) <= place_87_top;
  loopexit_d_1_to_loopexit_d_2_src_tip(0) <= place_99_top;
  loopexit_d_1_to_no_exit_d_2_d_preheader_src_tip(0) <= place_99_top;
  ni_d_0_d_0_mux_1_d_ack_tip(0) <= place_36_top;
  ni_d_0_d_0_mux_1_d_req0_tip(0) <= place_38_top;
  ni_d_0_d_0_mux_1_d_req1_tip(0) <= place_35_top;
  ni_d_1_d_0_mux_1_d_ack_tip(0) <= place_68_top;
  ni_d_1_d_0_mux_1_d_req0_tip(0) <= place_70_top;
  ni_d_1_d_0_mux_1_d_req1_tip(0) <= place_67_top;
  ni_d_1_d_1_mux_1_d_ack_tip(0) <= place_86_top;
  ni_d_1_d_1_mux_1_d_req0_tip(0) <= place_88_top;
  ni_d_1_d_1_mux_1_d_req1_tip(0) <= place_85_top;
  ni_d_1_mux_1_d_ack_tip(0) <= place_54_top;
  ni_d_1_mux_1_d_req0_tip(0) <= place_56_top;
  ni_d_1_mux_1_d_req1_tip(0) <= place_53_top;
  ni_d_2_d_0_mux_1_d_ack_tip(0) <= place_106_top;
  ni_d_2_d_0_mux_1_d_req0_tip(0) <= place_108_top;
  ni_d_2_d_0_mux_1_d_req1_tip(0) <= place_105_top;
  ni_d_2_d_1_mux_1_d_ack_tip(0) <= place_128_top;
  ni_d_2_d_1_mux_1_d_req0_tip(0) <= place_130_top;
  ni_d_2_d_1_mux_1_d_req1_tip(0) <= place_19_top;
  no_exit_d_0_d_entry_tip(0) <= place_5_top;
  no_exit_d_0_d_pre_tip(0) <= place_33_top;
  no_exit_d_0_d_pre_tip(1) <= place_37_top;
  no_exit_d_0_d_preheader_to_no_exit_d_0_src_tip(0) <= place_4_top;
  no_exit_d_0_to_loopentry_d_1_d_loopexit_src_tip(0) <= place_47_top;
  no_exit_d_0_to_no_exit_d_0_src_tip(0) <= place_47_top;
  no_exit_d_1_d_entry_tip(0) <= place_11_top;
  no_exit_d_1_d_pre_tip(0) <= place_65_top;
  no_exit_d_1_d_pre_tip(1) <= place_69_top;
  no_exit_d_1_d_preheader_to_no_exit_d_1_src_tip(0) <= place_9_top;
  no_exit_d_1_to_loopexit_d_1_d_loopexit_src_tip(0) <= place_79_top;
  no_exit_d_1_to_no_exit_d_1_src_tip(0) <= place_79_top;
  no_exit_d_2_d_entry_tip(0) <= place_17_top;
  no_exit_d_2_d_pre_tip(0) <= place_103_top;
  no_exit_d_2_d_pre_tip(1) <= place_107_top;
  no_exit_d_2_d_pre_tip(2) <= place_111_top;
  no_exit_d_2_d_preheader_to_no_exit_d_2_src_tip(0) <= place_15_top;
  no_exit_d_2_to_loopexit_d_2_d_loopexit_src_tip(0) <= place_125_top;
  no_exit_d_2_to_no_exit_d_2_src_tip(0) <= place_125_top;
  oper_tmp_d_1114_bool_d_ack_tip(0) <= place_76_top;
  oper_tmp_d_1114_bool_d_req_tip(0) <= place_77_top;
  oper_tmp_d_11_bool_d_ack_tip(0) <= place_58_top;
  oper_tmp_d_11_bool_d_req_tip(0) <= place_59_top;
  oper_tmp_d_14_float_d_ack_tip(0) <= place_71_top;
  oper_tmp_d_14_float_d_req_tip(0) <= place_72_top;
  oper_tmp_d_16_float_d_ack_tip(0) <= place_73_top;
  oper_tmp_d_16_float_d_req_tip(0) <= place_74_top;
  oper_tmp_d_19_float_d_ack_tip(0) <= place_89_top;
  oper_tmp_d_19_float_d_req_tip(0) <= place_90_top;
  oper_tmp_d_21_float_d_ack_tip(0) <= place_91_top;
  oper_tmp_d_21_float_d_req_tip(0) <= place_92_top;
  oper_tmp_d_2420_float_d_ack_tip(0) <= place_94_top;
  oper_tmp_d_2420_float_d_req_tip(0) <= place_95_top;
  oper_tmp_d_24_float_d_ack_tip(0) <= place_120_top;
  oper_tmp_d_24_float_d_req_tip(0) <= place_121_top;
  oper_tmp_d_2621_bool_d_ack_tip(0) <= place_96_top;
  oper_tmp_d_2621_bool_d_req_tip(0) <= place_97_top;
  oper_tmp_d_26_bool_d_ack_tip(0) <= place_122_top;
  oper_tmp_d_26_bool_d_req_tip(0) <= place_123_top;
  oper_tmp_d_31_float_d_ack_tip(0) <= place_113_top;
  oper_tmp_d_31_float_d_req_tip(0) <= place_114_top;
  oper_tmp_d_34_float_d_ack_tip(0) <= place_115_top;
  oper_tmp_d_34_float_d_req_tip(0) <= place_116_top;
  oper_tmp_d_35_bool_d_ack_tip(0) <= place_26_top;
  oper_tmp_d_35_bool_d_req_tip(0) <= place_1_top;
  oper_tmp_d_36_float_d_ack_tip(0) <= place_117_top;
  oper_tmp_d_36_float_d_req_tip(0) <= place_118_top;
  oper_tmp_d_3_bool_d_ack_tip(0) <= place_44_top;
  oper_tmp_d_3_bool_d_req_tip(0) <= place_45_top;
  oper_tmp_d_6_float_d_ack_tip(0) <= place_39_top;
  oper_tmp_d_6_float_d_req_tip(0) <= place_40_top;
  oper_tmp_d_8_float_d_ack_tip(0) <= place_41_top;
  oper_tmp_d_8_float_d_req_tip(0) <= place_42_top;
  ri_d_0_d_0_mux_1_d_ack_tip(0) <= place_110_top;
  ri_d_0_d_0_mux_1_d_req0_tip(0) <= place_112_top;
  ri_d_0_d_0_mux_1_d_req1_tip(0) <= place_109_top;
  store_location_divide_return_d_ack_tip(0) <= place_131_top;
  store_location_divide_return_d_req_tip(0) <= place_129_top;

  cbr_0_oper_tmp_d_35_bool_d_req_ge <= '1';
  op(5) <= cbr_0_oper_tmp_d_35_bool_d_req_top;
  cbr_1_oper_tmp_d_3_bool_d_req_ge <= '1';
  op(13) <= cbr_1_oper_tmp_d_3_bool_d_req_top;
  cbr_2_oper_tmp_d_11_bool_d_req_ge <= '1';
  op(19) <= cbr_2_oper_tmp_d_11_bool_d_req_top;
  cbr_3_oper_tmp_d_1114_bool_d_req_ge <= '1';
  op(27) <= cbr_3_oper_tmp_d_1114_bool_d_req_top;
  cbr_4_oper_tmp_d_2621_bool_d_req_ge <= '1';
  op(36) <= cbr_4_oper_tmp_d_2621_bool_d_req_top;
  cbr_5_oper_tmp_d_26_bool_d_req_ge <= '1';
  op(48) <= cbr_5_oper_tmp_d_26_bool_d_req_top;
  di_d_0_d_0_mux_1_d_ack_ge <= ip(7);
  di_d_0_d_0_mux_1_d_req0_ge <= '1';
  op(7) <= di_d_0_d_0_mux_1_d_req0_top;
  di_d_0_d_0_mux_1_d_req1_ge <= '1';
  op(6) <= di_d_0_d_0_mux_1_d_req1_top;
  di_d_1_d_0_mux_1_d_ack_ge <= ip(19);
  di_d_1_d_0_mux_1_d_req0_ge <= '1';
  op(21) <= di_d_1_d_0_mux_1_d_req0_top;
  di_d_1_d_0_mux_1_d_req1_ge <= '1';
  op(20) <= di_d_1_d_0_mux_1_d_req1_top;
  di_d_1_d_1_mux_1_d_ack_ge <= ip(26);
  di_d_1_d_1_mux_1_d_req0_ge <= '1';
  op(29) <= di_d_1_d_1_mux_1_d_req0_top;
  di_d_1_d_1_mux_1_d_req1_ge <= '1';
  op(28) <= di_d_1_d_1_mux_1_d_req1_top;
  di_d_1_mux_1_d_ack_ge <= ip(14);
  di_d_1_mux_1_d_req0_ge <= '1';
  op(15) <= di_d_1_mux_1_d_req0_top;
  di_d_1_mux_1_d_req1_ge <= '1';
  op(14) <= di_d_1_mux_1_d_req1_top;
  di_d_2_d_0_mux_1_d_ack_ge <= ip(34);
  di_d_2_d_0_mux_1_d_req0_ge <= '1';
  op(38) <= di_d_2_d_0_mux_1_d_req0_top;
  di_d_2_d_0_mux_1_d_req1_ge <= '1';
  op(37) <= di_d_2_d_0_mux_1_d_req1_top;
  entry_to_loopentry_d_1_src_ge <= ip(5);
  entry_to_no_exit_d_0_d_preheader_src_ge <= ip(6);
  fin_ge <= '1';
  op(1) <= fin_top;
  init_ge <= ip(1);
  load_dividend_d_ack_ge <= ip(2);
  load_dividend_d_req_ge <= '1';
  op(2) <= load_dividend_d_req_top;
  load_divisor_d_ack_ge <= ip(3);
  load_divisor_d_req_ge <= '1';
  op(3) <= load_divisor_d_req_top;
  loopentry_d_1_d_entry_ge <= '1';
  loopentry_d_1_d_loopexit_to_loopentry_d_1_src_ge <= '1';
  loopentry_d_1_d_pre_ge <= '1';
  loopentry_d_1_to_loopexit_d_1_src_ge <= ip(18);
  loopentry_d_1_to_no_exit_d_1_d_preheader_src_ge <= ip(17);
  loopexit_d_1_d_entry_ge <= '1';
  loopexit_d_1_d_loopexit_to_loopexit_d_1_src_ge <= '1';
  loopexit_d_1_d_pre_ge <= '1';
  loopexit_d_1_to_loopexit_d_2_src_ge <= ip(33);
  loopexit_d_1_to_no_exit_d_2_d_preheader_src_ge <= ip(32);
  ni_d_0_d_0_mux_1_d_ack_ge <= ip(8);
  ni_d_0_d_0_mux_1_d_req0_ge <= '1';
  op(9) <= ni_d_0_d_0_mux_1_d_req0_top;
  ni_d_0_d_0_mux_1_d_req1_ge <= '1';
  op(8) <= ni_d_0_d_0_mux_1_d_req1_top;
  ni_d_1_d_0_mux_1_d_ack_ge <= ip(20);
  ni_d_1_d_0_mux_1_d_req0_ge <= '1';
  op(23) <= ni_d_1_d_0_mux_1_d_req0_top;
  ni_d_1_d_0_mux_1_d_req1_ge <= '1';
  op(22) <= ni_d_1_d_0_mux_1_d_req1_top;
  ni_d_1_d_1_mux_1_d_ack_ge <= ip(27);
  ni_d_1_d_1_mux_1_d_req0_ge <= '1';
  op(31) <= ni_d_1_d_1_mux_1_d_req0_top;
  ni_d_1_d_1_mux_1_d_req1_ge <= '1';
  op(30) <= ni_d_1_d_1_mux_1_d_req1_top;
  ni_d_1_mux_1_d_ack_ge <= ip(15);
  ni_d_1_mux_1_d_req0_ge <= '1';
  op(17) <= ni_d_1_mux_1_d_req0_top;
  ni_d_1_mux_1_d_req1_ge <= '1';
  op(16) <= ni_d_1_mux_1_d_req1_top;
  ni_d_2_d_0_mux_1_d_ack_ge <= ip(35);
  ni_d_2_d_0_mux_1_d_req0_ge <= '1';
  op(40) <= ni_d_2_d_0_mux_1_d_req0_top;
  ni_d_2_d_0_mux_1_d_req1_ge <= '1';
  op(39) <= ni_d_2_d_0_mux_1_d_req1_top;
  ni_d_2_d_1_mux_1_d_ack_ge <= ip(44);
  ni_d_2_d_1_mux_1_d_req0_ge <= '1';
  op(50) <= ni_d_2_d_1_mux_1_d_req0_top;
  ni_d_2_d_1_mux_1_d_req1_ge <= '1';
  op(49) <= ni_d_2_d_1_mux_1_d_req1_top;
  no_exit_d_0_d_entry_ge <= '1';
  no_exit_d_0_d_pre_ge <= '1';
  no_exit_d_0_d_preheader_to_no_exit_d_0_src_ge <= '1';
  no_exit_d_0_to_loopentry_d_1_d_loopexit_src_ge <= ip(12);
  no_exit_d_0_to_no_exit_d_0_src_ge <= ip(13);
  no_exit_d_1_d_entry_ge <= '1';
  no_exit_d_1_d_pre_ge <= '1';
  no_exit_d_1_d_preheader_to_no_exit_d_1_src_ge <= '1';
  no_exit_d_1_to_loopexit_d_1_d_loopexit_src_ge <= ip(25);
  no_exit_d_1_to_no_exit_d_1_src_ge <= ip(24);
  no_exit_d_2_d_entry_ge <= '1';
  no_exit_d_2_d_pre_ge <= '1';
  no_exit_d_2_d_preheader_to_no_exit_d_2_src_ge <= '1';
  no_exit_d_2_to_loopexit_d_2_d_loopexit_src_ge <= ip(43);
  no_exit_d_2_to_no_exit_d_2_src_ge <= ip(42);
  oper_tmp_d_1114_bool_d_ack_ge <= ip(23);
  oper_tmp_d_1114_bool_d_req_ge <= '1';
  op(26) <= oper_tmp_d_1114_bool_d_req_top;
  oper_tmp_d_11_bool_d_ack_ge <= ip(16);
  oper_tmp_d_11_bool_d_req_ge <= '1';
  op(18) <= oper_tmp_d_11_bool_d_req_top;
  oper_tmp_d_14_float_d_ack_ge <= ip(21);
  oper_tmp_d_14_float_d_req_ge <= '1';
  op(24) <= oper_tmp_d_14_float_d_req_top;
  oper_tmp_d_16_float_d_ack_ge <= ip(22);
  oper_tmp_d_16_float_d_req_ge <= '1';
  op(25) <= oper_tmp_d_16_float_d_req_top;
  oper_tmp_d_19_float_d_ack_ge <= ip(28);
  oper_tmp_d_19_float_d_req_ge <= '1';
  op(32) <= oper_tmp_d_19_float_d_req_top;
  oper_tmp_d_21_float_d_ack_ge <= ip(29);
  oper_tmp_d_21_float_d_req_ge <= '1';
  op(33) <= oper_tmp_d_21_float_d_req_top;
  oper_tmp_d_2420_float_d_ack_ge <= ip(30);
  oper_tmp_d_2420_float_d_req_ge <= '1';
  op(34) <= oper_tmp_d_2420_float_d_req_top;
  oper_tmp_d_24_float_d_ack_ge <= ip(40);
  oper_tmp_d_24_float_d_req_ge <= '1';
  op(46) <= oper_tmp_d_24_float_d_req_top;
  oper_tmp_d_2621_bool_d_ack_ge <= ip(31);
  oper_tmp_d_2621_bool_d_req_ge <= '1';
  op(35) <= oper_tmp_d_2621_bool_d_req_top;
  oper_tmp_d_26_bool_d_ack_ge <= ip(41);
  oper_tmp_d_26_bool_d_req_ge <= '1';
  op(47) <= oper_tmp_d_26_bool_d_req_top;
  oper_tmp_d_31_float_d_ack_ge <= ip(37);
  oper_tmp_d_31_float_d_req_ge <= '1';
  op(43) <= oper_tmp_d_31_float_d_req_top;
  oper_tmp_d_34_float_d_ack_ge <= ip(38);
  oper_tmp_d_34_float_d_req_ge <= '1';
  op(44) <= oper_tmp_d_34_float_d_req_top;
  oper_tmp_d_35_bool_d_ack_ge <= ip(4);
  oper_tmp_d_35_bool_d_req_ge <= '1';
  op(4) <= oper_tmp_d_35_bool_d_req_top;
  oper_tmp_d_36_float_d_ack_ge <= ip(39);
  oper_tmp_d_36_float_d_req_ge <= '1';
  op(45) <= oper_tmp_d_36_float_d_req_top;
  oper_tmp_d_3_bool_d_ack_ge <= ip(11);
  oper_tmp_d_3_bool_d_req_ge <= '1';
  op(12) <= oper_tmp_d_3_bool_d_req_top;
  oper_tmp_d_6_float_d_ack_ge <= ip(9);
  oper_tmp_d_6_float_d_req_ge <= '1';
  op(10) <= oper_tmp_d_6_float_d_req_top;
  oper_tmp_d_8_float_d_ack_ge <= ip(10);
  oper_tmp_d_8_float_d_req_ge <= '1';
  op(11) <= oper_tmp_d_8_float_d_req_top;
  ri_d_0_d_0_mux_1_d_ack_ge <= ip(36);
  ri_d_0_d_0_mux_1_d_req0_ge <= '1';
  op(42) <= ri_d_0_d_0_mux_1_d_req0_top;
  ri_d_0_d_0_mux_1_d_req1_ge <= '1';
  op(41) <= ri_d_0_d_0_mux_1_d_req1_top;
  store_location_divide_return_d_ack_ge <= ip(45);
  store_location_divide_return_d_req_ge <= '1';
  op(51) <= store_location_divide_return_d_req_top;

end behavioral;
