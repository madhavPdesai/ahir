package GlobalConstants is
    constant global_debug_flag: boolean := false;
end package GlobalConstants;
