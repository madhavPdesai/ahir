-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity getData is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(3 downto 0);
    in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity getData;
architecture Default of getData is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal getData_CP_660_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_213_root_address_inst_ack_0 : boolean;
  signal ptr_deref_235_base_resize_req_0 : boolean;
  signal ptr_deref_235_base_resize_ack_0 : boolean;
  signal ptr_deref_213_store_0_req_1 : boolean;
  signal ptr_deref_230_base_resize_ack_0 : boolean;
  signal ptr_deref_182_store_0_ack_0 : boolean;
  signal ptr_deref_182_store_0_req_0 : boolean;
  signal ptr_deref_218_load_0_ack_1 : boolean;
  signal ptr_deref_218_load_0_req_1 : boolean;
  signal ptr_deref_213_store_0_ack_0 : boolean;
  signal ptr_deref_230_store_0_ack_1 : boolean;
  signal ptr_deref_230_base_resize_req_0 : boolean;
  signal ptr_deref_213_root_address_inst_req_0 : boolean;
  signal ptr_deref_218_addr_0_req_0 : boolean;
  signal array_obj_ref_226_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_226_index_0_resize_req_0 : boolean;
  signal ptr_deref_222_gather_scatter_ack_0 : boolean;
  signal ptr_deref_222_gather_scatter_req_0 : boolean;
  signal ptr_deref_230_store_0_req_1 : boolean;
  signal ptr_deref_235_load_0_ack_1 : boolean;
  signal ptr_deref_235_gather_scatter_req_0 : boolean;
  signal ptr_deref_235_gather_scatter_ack_0 : boolean;
  signal ptr_deref_222_load_0_req_0 : boolean;
  signal ptr_deref_182_addr_0_req_0 : boolean;
  signal ptr_deref_182_gather_scatter_ack_0 : boolean;
  signal ptr_deref_222_load_0_ack_1 : boolean;
  signal ptr_deref_222_load_0_req_1 : boolean;
  signal ptr_deref_218_load_0_ack_0 : boolean;
  signal ptr_deref_235_load_0_req_1 : boolean;
  signal ptr_deref_218_load_0_req_0 : boolean;
  signal ptr_deref_182_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_210_inst_ack_0 : boolean;
  signal ptr_deref_213_store_0_req_0 : boolean;
  signal ptr_deref_182_addr_0_ack_0 : boolean;
  signal array_obj_ref_226_index_0_rename_ack_0 : boolean;
  signal ptr_deref_222_load_0_ack_0 : boolean;
  signal array_obj_ref_226_root_address_inst_req_0 : boolean;
  signal ptr_deref_190_addr_0_ack_0 : boolean;
  signal ptr_deref_190_addr_0_req_0 : boolean;
  signal ptr_deref_182_store_0_ack_1 : boolean;
  signal ptr_deref_182_store_0_req_1 : boolean;
  signal simple_obj_ref_210_inst_req_0 : boolean;
  signal array_obj_ref_226_index_0_rename_req_0 : boolean;
  signal if_stmt_202_branch_ack_0 : boolean;
  signal ptr_deref_190_root_address_inst_ack_0 : boolean;
  signal ptr_deref_190_root_address_inst_req_0 : boolean;
  signal ptr_deref_182_root_address_inst_ack_0 : boolean;
  signal ptr_deref_222_addr_0_ack_0 : boolean;
  signal ptr_deref_182_root_address_inst_req_0 : boolean;
  signal ptr_deref_222_addr_0_req_0 : boolean;
  signal if_stmt_202_branch_ack_1 : boolean;
  signal ptr_deref_190_gather_scatter_ack_0 : boolean;
  signal ptr_deref_190_base_resize_ack_0 : boolean;
  signal addr_of_227_final_reg_ack_0 : boolean;
  signal addr_of_227_final_reg_req_0 : boolean;
  signal ptr_deref_213_addr_0_ack_0 : boolean;
  signal ptr_deref_190_base_resize_req_0 : boolean;
  signal ptr_deref_218_root_address_inst_ack_0 : boolean;
  signal ptr_deref_218_addr_0_ack_0 : boolean;
  signal ptr_deref_230_gather_scatter_req_0 : boolean;
  signal ptr_deref_230_addr_0_req_0 : boolean;
  signal ptr_deref_213_gather_scatter_req_0 : boolean;
  signal ptr_deref_230_store_0_ack_0 : boolean;
  signal ptr_deref_230_store_0_req_0 : boolean;
  signal ptr_deref_230_addr_0_ack_0 : boolean;
  signal ptr_deref_239_addr_0_req_0 : boolean;
  signal ptr_deref_239_addr_0_ack_0 : boolean;
  signal ptr_deref_239_base_resize_req_0 : boolean;
  signal ptr_deref_235_root_address_inst_ack_0 : boolean;
  signal ptr_deref_230_root_address_inst_ack_0 : boolean;
  signal ptr_deref_230_root_address_inst_req_0 : boolean;
  signal ptr_deref_239_base_resize_ack_0 : boolean;
  signal ptr_deref_235_root_address_inst_req_0 : boolean;
  signal ptr_deref_235_addr_0_req_0 : boolean;
  signal ptr_deref_235_load_0_req_0 : boolean;
  signal ptr_deref_235_load_0_ack_0 : boolean;
  signal ptr_deref_239_root_address_inst_req_0 : boolean;
  signal ptr_deref_239_root_address_inst_ack_0 : boolean;
  signal ptr_deref_190_gather_scatter_req_0 : boolean;
  signal ptr_deref_190_load_0_ack_1 : boolean;
  signal ptr_deref_190_load_0_req_1 : boolean;
  signal if_stmt_202_branch_req_0 : boolean;
  signal ptr_deref_190_load_0_ack_0 : boolean;
  signal ptr_deref_190_load_0_req_0 : boolean;
  signal ptr_deref_222_root_address_inst_ack_0 : boolean;
  signal ptr_deref_182_base_resize_ack_0 : boolean;
  signal ptr_deref_218_root_address_inst_req_0 : boolean;
  signal ptr_deref_222_root_address_inst_req_0 : boolean;
  signal ptr_deref_182_base_resize_req_0 : boolean;
  signal binary_199_inst_ack_1 : boolean;
  signal ptr_deref_213_gather_scatter_ack_0 : boolean;
  signal ptr_deref_218_base_resize_ack_0 : boolean;
  signal ptr_deref_222_base_resize_ack_0 : boolean;
  signal ptr_deref_218_gather_scatter_ack_0 : boolean;
  signal ptr_deref_222_base_resize_req_0 : boolean;
  signal binary_199_inst_req_1 : boolean;
  signal ptr_deref_218_base_resize_req_0 : boolean;
  signal ptr_deref_218_gather_scatter_req_0 : boolean;
  signal binary_199_inst_ack_0 : boolean;
  signal binary_199_inst_req_0 : boolean;
  signal array_obj_ref_226_offset_inst_ack_0 : boolean;
  signal ptr_deref_213_store_0_ack_1 : boolean;
  signal array_obj_ref_226_offset_inst_req_0 : boolean;
  signal type_cast_195_inst_ack_0 : boolean;
  signal type_cast_195_inst_req_0 : boolean;
  signal ptr_deref_213_base_resize_ack_0 : boolean;
  signal ptr_deref_213_addr_0_req_0 : boolean;
  signal ptr_deref_213_base_resize_req_0 : boolean;
  signal array_obj_ref_226_root_address_inst_ack_0 : boolean;
  signal ptr_deref_230_gather_scatter_ack_0 : boolean;
  signal ptr_deref_235_addr_0_ack_0 : boolean;
  signal ptr_deref_239_load_0_req_0 : boolean;
  signal ptr_deref_239_load_0_ack_0 : boolean;
  signal ptr_deref_239_load_0_req_1 : boolean;
  signal ptr_deref_239_load_0_ack_1 : boolean;
  signal ptr_deref_239_gather_scatter_req_0 : boolean;
  signal ptr_deref_239_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_243_index_0_resize_req_0 : boolean;
  signal array_obj_ref_243_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_243_index_0_rename_req_0 : boolean;
  signal array_obj_ref_243_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_243_offset_inst_req_0 : boolean;
  signal array_obj_ref_243_offset_inst_ack_0 : boolean;
  signal array_obj_ref_243_root_address_inst_req_0 : boolean;
  signal array_obj_ref_243_root_address_inst_ack_0 : boolean;
  signal addr_of_244_final_reg_req_0 : boolean;
  signal addr_of_244_final_reg_ack_0 : boolean;
  signal ptr_deref_247_base_resize_req_0 : boolean;
  signal ptr_deref_247_base_resize_ack_0 : boolean;
  signal ptr_deref_247_root_address_inst_req_0 : boolean;
  signal ptr_deref_247_root_address_inst_ack_0 : boolean;
  signal ptr_deref_247_addr_0_req_0 : boolean;
  signal ptr_deref_247_addr_0_ack_0 : boolean;
  signal ptr_deref_247_gather_scatter_req_0 : boolean;
  signal ptr_deref_247_gather_scatter_ack_0 : boolean;
  signal ptr_deref_247_store_0_req_0 : boolean;
  signal ptr_deref_247_store_0_ack_0 : boolean;
  signal ptr_deref_247_store_0_req_1 : boolean;
  signal ptr_deref_247_store_0_ack_1 : boolean;
  signal ptr_deref_254_base_resize_req_0 : boolean;
  signal ptr_deref_254_base_resize_ack_0 : boolean;
  signal ptr_deref_254_root_address_inst_req_0 : boolean;
  signal ptr_deref_254_root_address_inst_ack_0 : boolean;
  signal ptr_deref_254_addr_0_req_0 : boolean;
  signal ptr_deref_254_addr_0_ack_0 : boolean;
  signal ptr_deref_254_load_0_req_0 : boolean;
  signal ptr_deref_254_load_0_ack_0 : boolean;
  signal ptr_deref_254_load_0_req_1 : boolean;
  signal ptr_deref_254_load_0_ack_1 : boolean;
  signal ptr_deref_254_gather_scatter_req_0 : boolean;
  signal ptr_deref_254_gather_scatter_ack_0 : boolean;
  signal binary_260_inst_req_0 : boolean;
  signal binary_260_inst_ack_0 : boolean;
  signal binary_260_inst_req_1 : boolean;
  signal binary_260_inst_ack_1 : boolean;
  signal ptr_deref_263_base_resize_req_0 : boolean;
  signal ptr_deref_263_base_resize_ack_0 : boolean;
  signal ptr_deref_263_root_address_inst_req_0 : boolean;
  signal ptr_deref_263_root_address_inst_ack_0 : boolean;
  signal ptr_deref_263_addr_0_req_0 : boolean;
  signal ptr_deref_263_addr_0_ack_0 : boolean;
  signal ptr_deref_263_gather_scatter_req_0 : boolean;
  signal ptr_deref_263_gather_scatter_ack_0 : boolean;
  signal ptr_deref_263_store_0_req_0 : boolean;
  signal ptr_deref_263_store_0_ack_0 : boolean;
  signal ptr_deref_263_store_0_req_1 : boolean;
  signal ptr_deref_263_store_0_ack_1 : boolean;
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(1 downto 0);
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"getData start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"getData start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"getData fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"getData fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  getData_CP_660: Block -- control-path 
    signal cp_elements: BooleanArray(137 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(39);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(39), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 5 
    -- members (4) 
      -- 	branch_block_stmt_169/$entry
      -- 	$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185__entry__
      -- 	branch_block_stmt_169/branch_block_stmt_169__entry__
      -- 
    -- CP-element group 1 branch  place  bypass 
    -- predecessors 30 
    -- successors 34 31 
    -- members (2) 
      -- 	branch_block_stmt_169/if_stmt_202__entry__
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201__exit__
      -- 
    cp_elements(1) <= cp_elements(30);
    -- CP-element group 2 merge  transition  place  output  bypass 
    -- predecessors 37 137 
    -- successors 40 
    -- members (7) 
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_active_
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_trigger_
      -- 	branch_block_stmt_169/assign_stmt_211/$entry
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_complete/req
      -- 	branch_block_stmt_169/assign_stmt_211__entry__
      -- 	branch_block_stmt_169/merge_stmt_208__exit__
      -- 
    cp_elements(2) <= OrReduce(cp_elements(37) & cp_elements(137));
    req_862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => simple_obj_ref_210_inst_req_0); -- 
    -- CP-element group 3 transition  place  bypass 
    -- predecessors 110 
    -- successors 111 
    -- members (10) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265__entry__
      -- 	branch_block_stmt_169/merge_stmt_251__exit__
      -- 	branch_block_stmt_169/bb_2_bb_3
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249__exit__
      -- 	branch_block_stmt_169/bb_2_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_169/bb_2_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_169/merge_stmt_251_PhiReqMerge
      -- 	branch_block_stmt_169/merge_stmt_251_PhiAck/$entry
      -- 	branch_block_stmt_169/merge_stmt_251_PhiAck/$exit
      -- 	branch_block_stmt_169/merge_stmt_251_PhiAck/dummy
      -- 
    cp_elements(3) <= cp_elements(110);
    -- CP-element group 4 transition  place  bypass 
    -- predecessors 133 
    -- successors 134 
    -- members (4) 
      -- 	branch_block_stmt_169/bb_3_bb_1
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265__exit__
      -- 	branch_block_stmt_169/bb_3_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_169/bb_3_bb_1_PhiReq/$exit
      -- 
    cp_elements(4) <= cp_elements(133);
    -- CP-element group 5 fork  transition  bypass 
    -- predecessors 0 
    -- successors 8 6 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/$entry
      -- 
    cp_elements(5) <= cp_elements(0);
    -- CP-element group 6 transition  bypass 
    -- predecessors 5 
    -- successors 7 
    -- members (2) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/assign_stmt_185_active_
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/assign_stmt_185_trigger_
      -- 
    cp_elements(6) <= cp_elements(5);
    -- CP-element group 7 join  transition  output  no-bypass 
    -- predecessors 11 6 
    -- successors 12 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/split_req
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_trigger_
      -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(11);
      predecessors(1) <= cp_elements(6);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(7)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_182_gather_scatter_req_0); -- 
    -- CP-element group 8 transition  output  bypass 
    -- predecessors 5 
    -- successors 9 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/simple_obj_ref_181_trigger_
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/simple_obj_ref_181_completed_
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/simple_obj_ref_181_active_
      -- 
    cp_elements(8) <= cp_elements(5);
    base_resize_req_709_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => ptr_deref_182_base_resize_req_0); -- 
    -- CP-element group 9 transition  input  output  no-bypass 
    -- predecessors 8 
    -- successors 10 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_address_resized
      -- 
    base_resize_ack_710_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_base_resize_ack_0, ack => cp_elements(9)); -- 
    sum_rename_req_714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => ptr_deref_182_root_address_inst_req_0); -- 
    -- CP-element group 10 transition  input  output  no-bypass 
    -- predecessors 9 
    -- successors 11 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_root_address_calculated
      -- 
    sum_rename_ack_715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_root_address_inst_ack_0, ack => cp_elements(10)); -- 
    root_register_req_719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_182_addr_0_req_0); -- 
    -- CP-element group 11 transition  input  no-bypass 
    -- predecessors 10 
    -- successors 7 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_word_address_calculated
      -- 
    root_register_ack_720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_addr_0_ack_0, ack => cp_elements(11)); -- 
    -- CP-element group 12 transition  input  output  no-bypass 
    -- predecessors 7 
    -- successors 13 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/split_ack
      -- 
    split_ack_725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_gather_scatter_ack_0, ack => cp_elements(12)); -- 
    rr_732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => ptr_deref_182_store_0_req_0); -- 
    -- CP-element group 13 transition  input  output  no-bypass 
    -- predecessors 12 
    -- successors 14 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_active_
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/$entry
      -- 
    ra_733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_store_0_ack_0, ack => cp_elements(13)); -- 
    cr_743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_182_store_0_req_1); -- 
    -- CP-element group 14 transition  place  input  no-bypass 
    -- predecessors 13 
    -- successors 134 
    -- members (11) 
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_completed_
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/assign_stmt_185_completed_
      -- 	branch_block_stmt_169/bb_0_bb_1
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185__exit__
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_176_to_assign_stmt_185/ptr_deref_182_complete/$exit
      -- 	branch_block_stmt_169/bb_0_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_169/bb_0_bb_1_PhiReq/$exit
      -- 
    ca_744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_182_store_0_ack_1, ack => cp_elements(14)); -- 
    -- CP-element group 15 fork  transition  bypass 
    -- predecessors 135 
    -- successors 23 16 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/$entry
      -- 
    cp_elements(15) <= cp_elements(135);
    -- CP-element group 16 transition  output  bypass 
    -- predecessors 15 
    -- successors 17 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_189_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_189_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_189_trigger_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_address_calculated
      -- 
    cp_elements(16) <= cp_elements(15);
    base_resize_req_764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_190_base_resize_req_0); -- 
    -- CP-element group 17 transition  input  output  no-bypass 
    -- predecessors 16 
    -- successors 18 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_address_resized
      -- 
    base_resize_ack_765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_base_resize_ack_0, ack => cp_elements(17)); -- 
    sum_rename_req_769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_190_root_address_inst_req_0); -- 
    -- CP-element group 18 transition  input  output  no-bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_root_address_calculated
      -- 
    sum_rename_ack_770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_root_address_inst_ack_0, ack => cp_elements(18)); -- 
    root_register_req_774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_190_addr_0_req_0); -- 
    -- CP-element group 19 transition  input  output  no-bypass 
    -- predecessors 18 
    -- successors 20 
    -- members (8) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_trigger_
      -- 
    root_register_ack_775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_addr_0_ack_0, ack => cp_elements(19)); -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_190_load_0_req_0); -- 
    -- CP-element group 20 transition  input  output  no-bypass 
    -- predecessors 19 
    -- successors 21 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/$entry
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_load_0_ack_0, ack => cp_elements(20)); -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_190_load_0_req_1); -- 
    -- CP-element group 21 transition  input  output  no-bypass 
    -- predecessors 20 
    -- successors 22 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/merge_req
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/word_access/$exit
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_load_0_ack_1, ack => cp_elements(21)); -- 
    merge_req_798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_190_gather_scatter_req_0); -- 
    -- CP-element group 22 transition  input  output  no-bypass 
    -- predecessors 21 
    -- successors 27 
    -- members (12) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_194_trigger_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_trigger_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_194_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/simple_obj_ref_194_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_complete/merge_ack
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/ptr_deref_190_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_191_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_191_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_191_trigger_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_complete/req
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_complete/$entry
      -- 
    merge_ack_799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_190_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    req_819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => type_cast_195_inst_req_0); -- 
    -- CP-element group 23 transition  bypass 
    -- predecessors 15 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_active_
      -- 
    cp_elements(23) <= cp_elements(15);
    -- CP-element group 24 join  transition  bypass 
    -- predecessors 28 29 
    -- successors 30 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_201_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_201_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/assign_stmt_201_trigger_
      -- 
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(28);
      predecessors(1) <= cp_elements(29);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(24)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 25 transition  output  bypass 
    -- predecessors 27 
    -- successors 28 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_sample_start_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Sample/rr
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Sample/$entry
      -- 
    cp_elements(25) <= cp_elements(27);
    rr_824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => binary_199_inst_req_0); -- 
    -- CP-element group 26 transition  output  bypass 
    -- predecessors 27 
    -- successors 29 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_update_start_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Update/$entry
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Update/cr
      -- 
    cp_elements(26) <= cp_elements(27);
    cr_829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_199_inst_req_1); -- 
    -- CP-element group 27 fork  transition  input  no-bypass 
    -- predecessors 22 
    -- successors 26 25 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_active_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_trigger_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_complete/ack
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/type_cast_195_complete/$exit
      -- 
    ack_820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_195_inst_ack_0, ack => cp_elements(27)); -- 
    -- CP-element group 28 transition  input  no-bypass 
    -- predecessors 25 
    -- successors 24 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_sample_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Sample/ra
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Sample/$exit
      -- 
    ra_825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_199_inst_ack_0, ack => cp_elements(28)); -- 
    -- CP-element group 29 transition  input  no-bypass 
    -- predecessors 26 
    -- successors 24 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_update_completed_
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Update/$exit
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/binary_199_Update/ca
      -- 
    ca_830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_199_inst_ack_1, ack => cp_elements(29)); -- 
    -- CP-element group 30 join  transition  no-bypass 
    -- predecessors 23 24 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201/$exit
      -- 
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(23);
      predecessors(1) <= cp_elements(24);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(30)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 31 transition  bypass 
    -- predecessors 1 
    -- successors 32 
    -- members (1) 
      -- 	branch_block_stmt_169/if_stmt_202_dead_link/$entry
      -- 
    cp_elements(31) <= cp_elements(1);
    -- CP-element group 32 transition  dead  bypass 
    -- predecessors 31 
    -- successors 33 
    -- members (1) 
      -- 	branch_block_stmt_169/if_stmt_202_dead_link/dead_transition
      -- 
    cp_elements(32) <= false;
    -- CP-element group 33 transition  place  bypass 
    -- predecessors 32 
    -- successors 136 
    -- members (4) 
      -- 	branch_block_stmt_169/merge_stmt_208__entry__
      -- 	branch_block_stmt_169/if_stmt_202__exit__
      -- 	branch_block_stmt_169/if_stmt_202_dead_link/$exit
      -- 	branch_block_stmt_169/merge_stmt_208_dead_link/$entry
      -- 
    cp_elements(33) <= cp_elements(32);
    -- CP-element group 34 transition  output  bypass 
    -- predecessors 1 
    -- successors 35 
    -- members (3) 
      -- 	branch_block_stmt_169/if_stmt_202_eval_test/branch_req
      -- 	branch_block_stmt_169/if_stmt_202_eval_test/$exit
      -- 	branch_block_stmt_169/if_stmt_202_eval_test/$entry
      -- 
    cp_elements(34) <= cp_elements(1);
    branch_req_838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => if_stmt_202_branch_req_0); -- 
    -- CP-element group 35 branch  place  bypass 
    -- predecessors 34 
    -- successors 36 38 
    -- members (1) 
      -- 	branch_block_stmt_169/simple_obj_ref_203_place
      -- 
    cp_elements(35) <= cp_elements(34);
    -- CP-element group 36 transition  bypass 
    -- predecessors 35 
    -- successors 37 
    -- members (1) 
      -- 	branch_block_stmt_169/if_stmt_202_if_link/$entry
      -- 
    cp_elements(36) <= cp_elements(35);
    -- CP-element group 37 transition  place  input  no-bypass 
    -- predecessors 36 
    -- successors 2 
    -- members (9) 
      -- 	branch_block_stmt_169/bb_1_bb_2
      -- 	branch_block_stmt_169/if_stmt_202_if_link/if_choice_transition
      -- 	branch_block_stmt_169/if_stmt_202_if_link/$exit
      -- 	branch_block_stmt_169/bb_1_bb_2_PhiReq/$entry
      -- 	branch_block_stmt_169/bb_1_bb_2_PhiReq/$exit
      -- 	branch_block_stmt_169/merge_stmt_208_PhiReqMerge
      -- 	branch_block_stmt_169/merge_stmt_208_PhiAck/$entry
      -- 	branch_block_stmt_169/merge_stmt_208_PhiAck/$exit
      -- 	branch_block_stmt_169/merge_stmt_208_PhiAck/dummy
      -- 
    if_choice_transition_843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_202_branch_ack_1, ack => cp_elements(37)); -- 
    -- CP-element group 38 transition  bypass 
    -- predecessors 35 
    -- successors 39 
    -- members (1) 
      -- 	branch_block_stmt_169/if_stmt_202_else_link/$entry
      -- 
    cp_elements(38) <= cp_elements(35);
    -- CP-element group 39 transition  place  input  no-bypass 
    -- predecessors 38 
    -- successors 
    -- members (21) 
      -- 	branch_block_stmt_169/$exit
      -- 	branch_block_stmt_169/merge_stmt_269__exit__
      -- 	$exit
      -- 	branch_block_stmt_169/return__
      -- 	branch_block_stmt_169/merge_stmt_267__exit__
      -- 	branch_block_stmt_169/bb_1_bb_4
      -- 	branch_block_stmt_169/if_stmt_202_else_link/else_choice_transition
      -- 	branch_block_stmt_169/if_stmt_202_else_link/$exit
      -- 	branch_block_stmt_169/branch_block_stmt_169__exit__
      -- 	branch_block_stmt_169/bb_1_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_169/bb_1_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_169/merge_stmt_267_PhiReqMerge
      -- 	branch_block_stmt_169/merge_stmt_267_PhiAck/$entry
      -- 	branch_block_stmt_169/merge_stmt_267_PhiAck/$exit
      -- 	branch_block_stmt_169/merge_stmt_267_PhiAck/dummy
      -- 	branch_block_stmt_169/return___PhiReq/$entry
      -- 	branch_block_stmt_169/return___PhiReq/$exit
      -- 	branch_block_stmt_169/merge_stmt_269_PhiReqMerge
      -- 	branch_block_stmt_169/merge_stmt_269_PhiAck/$entry
      -- 	branch_block_stmt_169/merge_stmt_269_PhiAck/$exit
      -- 	branch_block_stmt_169/merge_stmt_269_PhiAck/dummy
      -- 
    else_choice_transition_847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_202_branch_ack_0, ack => cp_elements(39)); -- 
    -- CP-element group 40 transition  place  input  no-bypass 
    -- predecessors 2 
    -- successors 41 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_completed_
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_complete/ack
      -- 	branch_block_stmt_169/assign_stmt_211/assign_stmt_211_completed_
      -- 	branch_block_stmt_169/assign_stmt_211/assign_stmt_211_active_
      -- 	branch_block_stmt_169/assign_stmt_211/assign_stmt_211_trigger_
      -- 	branch_block_stmt_169/assign_stmt_211/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249__entry__
      -- 	branch_block_stmt_169/assign_stmt_211__exit__
      -- 	branch_block_stmt_169/assign_stmt_211/simple_obj_ref_210_complete/$exit
      -- 
    ack_863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_210_inst_ack_0, ack => cp_elements(40)); -- 
    -- CP-element group 41 fork  transition  bypass 
    -- predecessors 40 
    -- successors 82 89 96 42 53 60 44 67 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/$entry
      -- 
    cp_elements(41) <= cp_elements(40);
    -- CP-element group 42 transition  bypass 
    -- predecessors 41 
    -- successors 43 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_214_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_214_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_214_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_215_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_215_trigger_
      -- 
    cp_elements(42) <= cp_elements(41);
    -- CP-element group 43 join  transition  output  bypass 
    -- predecessors 42 47 
    -- successors 48 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/split_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/$entry
      -- 
    cpelement_group_43 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(42);
      predecessors(1) <= cp_elements(47);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(43)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(43),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_213_gather_scatter_req_0); -- 
    -- CP-element group 44 transition  output  bypass 
    -- predecessors 41 
    -- successors 45 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_212_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_212_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_212_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_addr_resize/base_resize_req
      -- 
    cp_elements(44) <= cp_elements(41);
    base_resize_req_886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_213_base_resize_req_0); -- 
    -- CP-element group 45 transition  input  output  no-bypass 
    -- predecessors 44 
    -- successors 46 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_base_resize_ack_0, ack => cp_elements(45)); -- 
    sum_rename_req_891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_213_root_address_inst_req_0); -- 
    -- CP-element group 46 transition  input  output  no-bypass 
    -- predecessors 45 
    -- successors 47 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_word_addrgen/root_register_req
      -- 
    sum_rename_ack_892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_root_address_inst_ack_0, ack => cp_elements(46)); -- 
    root_register_req_896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_213_addr_0_req_0); -- 
    -- CP-element group 47 transition  input  no-bypass 
    -- predecessors 46 
    -- successors 43 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_word_addrgen/$exit
      -- 
    root_register_ack_897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_addr_0_ack_0, ack => cp_elements(47)); -- 
    -- CP-element group 48 transition  input  output  no-bypass 
    -- predecessors 43 
    -- successors 49 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/split_ack
      -- 
    split_ack_902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_gather_scatter_ack_0, ack => cp_elements(48)); -- 
    rr_909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_213_store_0_req_0); -- 
    -- CP-element group 49 fork  transition  input  no-bypass 
    -- predecessors 48 
    -- successors 81 50 52 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_active_
      -- 
    ra_910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_store_0_ack_0, ack => cp_elements(49)); -- 
    -- CP-element group 50 transition  output  bypass 
    -- predecessors 49 
    -- successors 51 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/$entry
      -- 
    cp_elements(50) <= cp_elements(49);
    cr_920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => ptr_deref_213_store_0_req_1); -- 
    -- CP-element group 51 transition  input  no-bypass 
    -- predecessors 50 
    -- successors 110 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_215_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_213_complete/word_access/word_access_0/ca
      -- 
    ca_921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_213_store_0_ack_1, ack => cp_elements(51)); -- 
    -- CP-element group 52 join  transition  output  bypass 
    -- predecessors 49 56 
    -- successors 57 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/$entry
      -- 
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(49);
      predecessors(1) <= cp_elements(56);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(52)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_218_load_0_req_0); -- 
    -- CP-element group 53 transition  output  bypass 
    -- predecessors 41 
    -- successors 54 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_217_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_217_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_217_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_address_calculated
      -- 
    cp_elements(53) <= cp_elements(41);
    base_resize_req_938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => ptr_deref_218_base_resize_req_0); -- 
    -- CP-element group 54 transition  input  output  no-bypass 
    -- predecessors 53 
    -- successors 55 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_plus_offset/$entry
      -- 
    base_resize_ack_939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_base_resize_ack_0, ack => cp_elements(54)); -- 
    sum_rename_req_943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_218_root_address_inst_req_0); -- 
    -- CP-element group 55 transition  input  output  no-bypass 
    -- predecessors 54 
    -- successors 56 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_base_plus_offset/$exit
      -- 
    sum_rename_ack_944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_root_address_inst_ack_0, ack => cp_elements(55)); -- 
    root_register_req_948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_218_addr_0_req_0); -- 
    -- CP-element group 56 transition  input  no-bypass 
    -- predecessors 55 
    -- successors 52 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_word_addrgen/root_register_ack
      -- 
    root_register_ack_949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_addr_0_ack_0, ack => cp_elements(56)); -- 
    -- CP-element group 57 transition  input  output  no-bypass 
    -- predecessors 52 
    -- successors 58 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_request/$exit
      -- 
    ra_960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_load_0_ack_0, ack => cp_elements(57)); -- 
    cr_970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => ptr_deref_218_load_0_req_1); -- 
    -- CP-element group 58 transition  input  output  no-bypass 
    -- predecessors 57 
    -- successors 59 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/merge_req
      -- 
    ca_971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_load_0_ack_1, ack => cp_elements(58)); -- 
    merge_req_972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_218_gather_scatter_req_0); -- 
    -- CP-element group 59 transition  input  no-bypass 
    -- predecessors 58 
    -- successors 74 
    -- members (11) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_231_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_232_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_231_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_219_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_232_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_219_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_219_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_231_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_218_complete/merge_ack
      -- 
    merge_ack_973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_218_gather_scatter_ack_0, ack => cp_elements(59)); -- 
    -- CP-element group 60 transition  output  bypass 
    -- predecessors 41 
    -- successors 61 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_221_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_221_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_221_active_
      -- 
    cp_elements(60) <= cp_elements(41);
    base_resize_req_990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => ptr_deref_222_base_resize_req_0); -- 
    -- CP-element group 61 transition  input  output  no-bypass 
    -- predecessors 60 
    -- successors 62 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_base_resize_ack_0, ack => cp_elements(61)); -- 
    sum_rename_req_995_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_222_root_address_inst_req_0); -- 
    -- CP-element group 62 transition  input  output  no-bypass 
    -- predecessors 61 
    -- successors 63 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_base_plus_offset/$exit
      -- 
    sum_rename_ack_996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_root_address_inst_ack_0, ack => cp_elements(62)); -- 
    root_register_req_1000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_222_addr_0_req_0); -- 
    -- CP-element group 63 transition  input  output  no-bypass 
    -- predecessors 62 
    -- successors 64 
    -- members (8) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_word_address_calculated
      -- 
    root_register_ack_1001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_addr_0_ack_0, ack => cp_elements(63)); -- 
    rr_1011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_222_load_0_req_0); -- 
    -- CP-element group 64 transition  input  output  no-bypass 
    -- predecessors 63 
    -- successors 65 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_request/$exit
      -- 
    ra_1012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_load_0_ack_0, ack => cp_elements(64)); -- 
    cr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_222_load_0_req_1); -- 
    -- CP-element group 65 transition  input  output  no-bypass 
    -- predecessors 64 
    -- successors 66 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/merge_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/word_access/$exit
      -- 
    ca_1023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_load_0_ack_1, ack => cp_elements(65)); -- 
    merge_req_1024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_222_gather_scatter_req_0); -- 
    -- CP-element group 66 transition  input  output  no-bypass 
    -- predecessors 65 
    -- successors 69 
    -- members (12) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_223_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_resize_0/index_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/merge_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_223_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_223_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_resize_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_222_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_225_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_225_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_225_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_computed_0
      -- 
    merge_ack_1025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_222_gather_scatter_ack_0, ack => cp_elements(66)); -- 
    index_resize_req_1043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => array_obj_ref_226_index_0_resize_req_0); -- 
    -- CP-element group 67 transition  bypass 
    -- predecessors 41 
    -- successors 68 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_trigger_
      -- 
    cp_elements(67) <= cp_elements(41);
    -- CP-element group 68 join  transition  output  bypass 
    -- predecessors 72 67 
    -- successors 73 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_complete/final_reg_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_active_
      -- 
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(72);
      predecessors(1) <= cp_elements(67);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(68)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => addr_of_227_final_reg_req_0); -- 
    -- CP-element group 69 transition  input  output  no-bypass 
    -- predecessors 66 
    -- successors 70 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_scale_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_resize_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_resized_0
      -- 
    index_resize_ack_1044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_226_index_0_resize_ack_0, ack => cp_elements(69)); -- 
    scale_rename_req_1048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_226_index_0_rename_req_0); -- 
    -- CP-element group 70 transition  input  output  no-bypass 
    -- predecessors 69 
    -- successors 71 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_add_indices/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_index_scale_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_indices_scaled
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_add_indices/final_index_req
      -- 
    scale_rename_ack_1049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_226_index_0_rename_ack_0, ack => cp_elements(70)); -- 
    final_index_req_1053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_226_offset_inst_req_0); -- 
    -- CP-element group 71 transition  input  output  no-bypass 
    -- predecessors 70 
    -- successors 72 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_add_indices/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_offset_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_add_indices/final_index_ack
      -- 
    final_index_ack_1054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_226_offset_inst_ack_0, ack => cp_elements(71)); -- 
    sum_rename_req_1058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_226_root_address_inst_req_0); -- 
    -- CP-element group 72 transition  input  no-bypass 
    -- predecessors 71 
    -- successors 68 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_226_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_226_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    -- CP-element group 73 transition  input  output  no-bypass 
    -- predecessors 68 
    -- successors 75 
    -- members (12) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_228_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_229_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_229_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_228_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_229_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_228_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_complete/final_reg_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_227_completed_
      -- 
    final_reg_ack_1064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_227_final_reg_ack_0, ack => cp_elements(73)); -- 
    base_resize_req_1084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => ptr_deref_230_base_resize_req_0); -- 
    -- CP-element group 74 join  transition  output  bypass 
    -- predecessors 77 59 
    -- successors 78 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/split_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_trigger_
      -- 
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(77);
      predecessors(1) <= cp_elements(59);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(74)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_1099_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_230_gather_scatter_req_0); -- 
    -- CP-element group 75 transition  input  output  no-bypass 
    -- predecessors 73 
    -- successors 76 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_base_resize_ack_0, ack => cp_elements(75)); -- 
    sum_rename_req_1089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => ptr_deref_230_root_address_inst_req_0); -- 
    -- CP-element group 76 transition  input  output  no-bypass 
    -- predecessors 75 
    -- successors 77 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_root_address_calculated
      -- 
    sum_rename_ack_1090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_root_address_inst_ack_0, ack => cp_elements(76)); -- 
    root_register_req_1094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_230_addr_0_req_0); -- 
    -- CP-element group 77 transition  input  no-bypass 
    -- predecessors 76 
    -- successors 74 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_word_addrgen/$exit
      -- 
    root_register_ack_1095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_addr_0_ack_0, ack => cp_elements(77)); -- 
    -- CP-element group 78 transition  input  output  no-bypass 
    -- predecessors 74 
    -- successors 79 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/split_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/word_access_0/$entry
      -- 
    split_ack_1100_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_gather_scatter_ack_0, ack => cp_elements(78)); -- 
    rr_1107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => ptr_deref_230_store_0_req_0); -- 
    -- CP-element group 79 transition  input  output  no-bypass 
    -- predecessors 78 
    -- successors 80 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_request/word_access/word_access_0/$exit
      -- 
    ra_1108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_store_0_ack_0, ack => cp_elements(79)); -- 
    cr_1118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_230_store_0_req_1); -- 
    -- CP-element group 80 transition  input  no-bypass 
    -- predecessors 79 
    -- successors 110 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_232_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_230_completed_
      -- 
    ca_1119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_230_store_0_ack_1, ack => cp_elements(80)); -- 
    -- CP-element group 81 join  transition  output  bypass 
    -- predecessors 85 49 
    -- successors 86 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_trigger_
      -- 
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(85);
      predecessors(1) <= cp_elements(49);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(81)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_235_load_0_req_0); -- 
    -- CP-element group 82 transition  output  bypass 
    -- predecessors 41 
    -- successors 83 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_234_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_234_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_234_active_
      -- 
    cp_elements(82) <= cp_elements(41);
    base_resize_req_1136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_235_base_resize_req_0); -- 
    -- CP-element group 83 transition  input  output  no-bypass 
    -- predecessors 82 
    -- successors 84 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_address_resized
      -- 
    base_resize_ack_1137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_base_resize_ack_0, ack => cp_elements(83)); -- 
    sum_rename_req_1141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_235_root_address_inst_req_0); -- 
    -- CP-element group 84 transition  input  output  no-bypass 
    -- predecessors 83 
    -- successors 85 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_root_address_inst_ack_0, ack => cp_elements(84)); -- 
    root_register_req_1146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_235_addr_0_req_0); -- 
    -- CP-element group 85 transition  input  no-bypass 
    -- predecessors 84 
    -- successors 81 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_word_addrgen/root_register_ack
      -- 
    root_register_ack_1147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_addr_0_ack_0, ack => cp_elements(85)); -- 
    -- CP-element group 86 transition  input  output  no-bypass 
    -- predecessors 81 
    -- successors 87 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_active_
      -- 
    ra_1158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_load_0_ack_0, ack => cp_elements(86)); -- 
    cr_1168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_235_load_0_req_1); -- 
    -- CP-element group 87 transition  input  output  no-bypass 
    -- predecessors 86 
    -- successors 88 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/merge_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/word_access/$exit
      -- 
    ca_1169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_load_0_ack_1, ack => cp_elements(87)); -- 
    merge_req_1170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => ptr_deref_235_gather_scatter_req_0); -- 
    -- CP-element group 88 transition  input  no-bypass 
    -- predecessors 87 
    -- successors 103 
    -- members (11) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/merge_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_236_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_236_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_236_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_235_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_249_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_249_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_248_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_248_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_248_completed_
      -- 
    merge_ack_1171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_235_gather_scatter_ack_0, ack => cp_elements(88)); -- 
    -- CP-element group 89 transition  output  bypass 
    -- predecessors 41 
    -- successors 90 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_238_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_238_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_238_completed_
      -- 
    cp_elements(89) <= cp_elements(41);
    base_resize_req_1188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_239_base_resize_req_0); -- 
    -- CP-element group 90 transition  input  output  no-bypass 
    -- predecessors 89 
    -- successors 91 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_base_resize_ack_0, ack => cp_elements(90)); -- 
    sum_rename_req_1193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => ptr_deref_239_root_address_inst_req_0); -- 
    -- CP-element group 91 transition  input  output  no-bypass 
    -- predecessors 90 
    -- successors 92 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_word_addrgen/root_register_req
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_word_addrgen/$entry
      -- 
    sum_rename_ack_1194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_root_address_inst_ack_0, ack => cp_elements(91)); -- 
    root_register_req_1198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => ptr_deref_239_addr_0_req_0); -- 
    -- CP-element group 92 transition  input  output  no-bypass 
    -- predecessors 91 
    -- successors 93 
    -- members (8) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/word_access_0/rr
      -- 
    root_register_ack_1199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_addr_0_ack_0, ack => cp_elements(92)); -- 
    rr_1209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_239_load_0_req_0); -- 
    -- CP-element group 93 transition  input  output  no-bypass 
    -- predecessors 92 
    -- successors 94 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/word_access_0/cr
      -- 
    ra_1210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_0, ack => cp_elements(93)); -- 
    cr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_239_load_0_req_1); -- 
    -- CP-element group 94 transition  input  output  no-bypass 
    -- predecessors 93 
    -- successors 95 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/merge_req
      -- 
    ca_1221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_load_0_ack_1, ack => cp_elements(94)); -- 
    merge_req_1222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_239_gather_scatter_req_0); -- 
    -- CP-element group 95 transition  input  output  no-bypass 
    -- predecessors 94 
    -- successors 98 
    -- members (12) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_240_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_240_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_240_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_239_complete/merge_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_computed_0
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_242_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_242_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_242_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_resize_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_resize_0/index_resize_req
      -- 
    merge_ack_1223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_239_gather_scatter_ack_0, ack => cp_elements(95)); -- 
    index_resize_req_1241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_243_index_0_resize_req_0); -- 
    -- CP-element group 96 transition  bypass 
    -- predecessors 41 
    -- successors 97 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_trigger_
      -- 
    cp_elements(96) <= cp_elements(41);
    -- CP-element group 97 join  transition  output  bypass 
    -- predecessors 96 101 
    -- successors 102 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_complete/final_reg_req
      -- 
    cpelement_group_97 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(96);
      predecessors(1) <= cp_elements(101);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(97)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(97),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => addr_of_244_final_reg_req_0); -- 
    -- CP-element group 98 transition  input  output  no-bypass 
    -- predecessors 95 
    -- successors 99 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_resized_0
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_resize_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_scale_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_1242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_index_0_resize_ack_0, ack => cp_elements(98)); -- 
    scale_rename_req_1246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_243_index_0_rename_req_0); -- 
    -- CP-element group 99 transition  input  output  no-bypass 
    -- predecessors 98 
    -- successors 100 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_indices_scaled
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_scale_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_add_indices/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_add_indices/final_index_req
      -- 
    scale_rename_ack_1247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_index_0_rename_ack_0, ack => cp_elements(99)); -- 
    final_index_req_1251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => array_obj_ref_243_offset_inst_req_0); -- 
    -- CP-element group 100 transition  input  output  no-bypass 
    -- predecessors 99 
    -- successors 101 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_offset_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_add_indices/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_add_indices/final_index_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_offset_inst_ack_0, ack => cp_elements(100)); -- 
    sum_rename_req_1256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => array_obj_ref_243_root_address_inst_req_0); -- 
    -- CP-element group 101 transition  input  no-bypass 
    -- predecessors 100 
    -- successors 97 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/array_obj_ref_243_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_243_root_address_inst_ack_0, ack => cp_elements(101)); -- 
    -- CP-element group 102 transition  input  output  no-bypass 
    -- predecessors 97 
    -- successors 104 
    -- members (12) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_245_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_245_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_245_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/addr_of_244_complete/final_reg_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_246_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_246_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/simple_obj_ref_246_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_1262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_244_final_reg_ack_0, ack => cp_elements(102)); -- 
    base_resize_req_1282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => ptr_deref_247_base_resize_req_0); -- 
    -- CP-element group 103 join  transition  output  bypass 
    -- predecessors 106 88 
    -- successors 107 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_trigger_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/split_req
      -- 
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(106);
      predecessors(1) <= cp_elements(88);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(103)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_1297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_247_gather_scatter_req_0); -- 
    -- CP-element group 104 transition  input  output  no-bypass 
    -- predecessors 102 
    -- successors 105 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_base_resize_ack_0, ack => cp_elements(104)); -- 
    sum_rename_req_1287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_247_root_address_inst_req_0); -- 
    -- CP-element group 105 transition  input  output  no-bypass 
    -- predecessors 104 
    -- successors 106 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_root_address_inst_ack_0, ack => cp_elements(105)); -- 
    root_register_req_1292_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_247_addr_0_req_0); -- 
    -- CP-element group 106 transition  input  no-bypass 
    -- predecessors 105 
    -- successors 103 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_word_addrgen/root_register_ack
      -- 
    root_register_ack_1293_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_addr_0_ack_0, ack => cp_elements(106)); -- 
    -- CP-element group 107 transition  input  output  no-bypass 
    -- predecessors 103 
    -- successors 108 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/split_ack
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/word_access_0/rr
      -- 
    split_ack_1298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_gather_scatter_ack_0, ack => cp_elements(107)); -- 
    rr_1305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_247_store_0_req_0); -- 
    -- CP-element group 108 transition  input  output  no-bypass 
    -- predecessors 107 
    -- successors 109 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_active_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/word_access_0/cr
      -- 
    ra_1306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_store_0_ack_0, ack => cp_elements(108)); -- 
    cr_1316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => ptr_deref_247_store_0_req_1); -- 
    -- CP-element group 109 transition  input  no-bypass 
    -- predecessors 108 
    -- successors 110 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/assign_stmt_249_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_completed_
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/ptr_deref_247_complete/word_access/word_access_0/ca
      -- 
    ca_1317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_247_store_0_ack_1, ack => cp_elements(109)); -- 
    -- CP-element group 110 join  transition  bypass 
    -- predecessors 80 109 51 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_215_to_assign_stmt_249/$exit
      -- 
    cpelement_group_110 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(80);
      predecessors(1) <= cp_elements(109);
      predecessors(2) <= cp_elements(51);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(110)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(110),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 111 fork  transition  bypass 
    -- predecessors 3 
    -- successors 112 119 126 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/$entry
      -- 
    cp_elements(111) <= cp_elements(3);
    -- CP-element group 112 transition  output  bypass 
    -- predecessors 111 
    -- successors 113 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_253_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_253_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_253_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_addr_resize/base_resize_req
      -- 
    cp_elements(112) <= cp_elements(111);
    base_resize_req_1337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => ptr_deref_254_base_resize_req_0); -- 
    -- CP-element group 113 transition  input  output  no-bypass 
    -- predecessors 112 
    -- successors 114 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_base_resize_ack_0, ack => cp_elements(113)); -- 
    sum_rename_req_1342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_254_root_address_inst_req_0); -- 
    -- CP-element group 114 transition  input  output  no-bypass 
    -- predecessors 113 
    -- successors 115 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_root_address_inst_ack_0, ack => cp_elements(114)); -- 
    root_register_req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_254_addr_0_req_0); -- 
    -- CP-element group 115 transition  input  output  no-bypass 
    -- predecessors 114 
    -- successors 116 
    -- members (8) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_word_addrgen/root_register_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/word_access_0/rr
      -- 
    root_register_ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_addr_0_ack_0, ack => cp_elements(115)); -- 
    rr_1358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_254_load_0_req_0); -- 
    -- CP-element group 116 transition  input  output  no-bypass 
    -- predecessors 115 
    -- successors 117 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/word_access_0/cr
      -- 
    ra_1359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_load_0_ack_0, ack => cp_elements(116)); -- 
    cr_1369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => ptr_deref_254_load_0_req_1); -- 
    -- CP-element group 117 transition  input  output  no-bypass 
    -- predecessors 116 
    -- successors 118 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/merge_req
      -- 
    ca_1370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_load_0_ack_1, ack => cp_elements(117)); -- 
    merge_req_1371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_254_gather_scatter_req_0); -- 
    -- CP-element group 118 fork  transition  input  no-bypass 
    -- predecessors 117 
    -- successors 121 122 
    -- members (10) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_255_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_255_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_255_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_254_complete/merge_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_257_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_257_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_257_completed_
      -- 
    merge_ack_1372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_254_gather_scatter_ack_0, ack => cp_elements(118)); -- 
    -- CP-element group 119 transition  bypass 
    -- predecessors 111 
    -- successors 133 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_active_
      -- 
    cp_elements(119) <= cp_elements(111);
    -- CP-element group 120 join  transition  bypass 
    -- predecessors 123 124 
    -- successors 125 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_261_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_261_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_261_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_265_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_265_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_264_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_264_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_264_completed_
      -- 
    cpelement_group_120 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(123);
      predecessors(1) <= cp_elements(124);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(120)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(120),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 121 transition  output  bypass 
    -- predecessors 118 
    -- successors 123 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_sample_start_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Sample/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Sample/rr
      -- 
    cp_elements(121) <= cp_elements(118);
    rr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => binary_260_inst_req_0); -- 
    -- CP-element group 122 transition  output  bypass 
    -- predecessors 118 
    -- successors 124 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_update_start_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Update/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Update/cr
      -- 
    cp_elements(122) <= cp_elements(118);
    cr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => binary_260_inst_req_1); -- 
    -- CP-element group 123 transition  input  no-bypass 
    -- predecessors 121 
    -- successors 120 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_sample_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Sample/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Sample/ra
      -- 
    ra_1390_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_260_inst_ack_0, ack => cp_elements(123)); -- 
    -- CP-element group 124 transition  input  no-bypass 
    -- predecessors 122 
    -- successors 120 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_update_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Update/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/binary_260_Update/ca
      -- 
    ca_1395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_260_inst_ack_1, ack => cp_elements(124)); -- 
    -- CP-element group 125 join  transition  output  bypass 
    -- predecessors 120 129 
    -- successors 130 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/split_req
      -- 
    cpelement_group_125 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(120);
      predecessors(1) <= cp_elements(129);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(125)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(125),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_1430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_263_gather_scatter_req_0); -- 
    -- CP-element group 126 transition  output  bypass 
    -- predecessors 111 
    -- successors 127 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_262_trigger_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_262_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/simple_obj_ref_262_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_addr_resize/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_addr_resize/base_resize_req
      -- 
    cp_elements(126) <= cp_elements(111);
    base_resize_req_1415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_263_base_resize_req_0); -- 
    -- CP-element group 127 transition  input  output  no-bypass 
    -- predecessors 126 
    -- successors 128 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_address_resized
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_addr_resize/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_plus_offset/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_base_resize_ack_0, ack => cp_elements(127)); -- 
    sum_rename_req_1420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(127), ack => ptr_deref_263_root_address_inst_req_0); -- 
    -- CP-element group 128 transition  input  output  no-bypass 
    -- predecessors 127 
    -- successors 129 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_root_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_plus_offset/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_word_addrgen/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_root_address_inst_ack_0, ack => cp_elements(128)); -- 
    root_register_req_1425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_263_addr_0_req_0); -- 
    -- CP-element group 129 transition  input  no-bypass 
    -- predecessors 128 
    -- successors 125 
    -- members (3) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_word_address_calculated
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_word_addrgen/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_word_addrgen/root_register_ack
      -- 
    root_register_ack_1426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_addr_0_ack_0, ack => cp_elements(129)); -- 
    -- CP-element group 130 transition  input  output  no-bypass 
    -- predecessors 125 
    -- successors 131 
    -- members (4) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/split_ack
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/word_access_0/rr
      -- 
    split_ack_1431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_gather_scatter_ack_0, ack => cp_elements(130)); -- 
    rr_1438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => ptr_deref_263_store_0_req_0); -- 
    -- CP-element group 131 transition  input  output  no-bypass 
    -- predecessors 130 
    -- successors 132 
    -- members (9) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_active_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/word_access_0/cr
      -- 
    ra_1439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_store_0_ack_0, ack => cp_elements(131)); -- 
    cr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_263_store_0_req_1); -- 
    -- CP-element group 132 transition  input  no-bypass 
    -- predecessors 131 
    -- successors 133 
    -- members (6) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/assign_stmt_265_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_completed_
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/ptr_deref_263_complete/word_access/word_access_0/ca
      -- 
    ca_1450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_263_store_0_ack_1, ack => cp_elements(132)); -- 
    -- CP-element group 133 join  transition  no-bypass 
    -- predecessors 119 132 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_169/assign_stmt_255_to_assign_stmt_265/$exit
      -- 
    cpelement_group_133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(119);
      predecessors(1) <= cp_elements(132);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(133)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 134 merge  place  bypass 
    -- predecessors 4 14 
    -- successors 135 
    -- members (1) 
      -- 	branch_block_stmt_169/merge_stmt_187_PhiReqMerge
      -- 
    cp_elements(134) <= OrReduce(cp_elements(4) & cp_elements(14));
    -- CP-element group 135 transition  place  bypass 
    -- predecessors 134 
    -- successors 15 
    -- members (5) 
      -- 	branch_block_stmt_169/assign_stmt_191_to_assign_stmt_201__entry__
      -- 	branch_block_stmt_169/merge_stmt_187__exit__
      -- 	branch_block_stmt_169/merge_stmt_187_PhiAck/$entry
      -- 	branch_block_stmt_169/merge_stmt_187_PhiAck/$exit
      -- 	branch_block_stmt_169/merge_stmt_187_PhiAck/dummy
      -- 
    cp_elements(135) <= cp_elements(134);
    -- CP-element group 136 transition  dead  bypass 
    -- predecessors 33 
    -- successors 137 
    -- members (1) 
      -- 	branch_block_stmt_169/merge_stmt_208_dead_link/dead_transition
      -- 
    cp_elements(136) <= false;
    -- CP-element group 137 transition  bypass 
    -- predecessors 136 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_169/merge_stmt_208_dead_link/$exit
      -- 
    cp_elements(137) <= cp_elements(136);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_226_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_226_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_226_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_226_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_243_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_243_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_243_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_243_root_address : std_logic_vector(6 downto 0);
    signal iNsTr_10_228 : std_logic_vector(31 downto 0);
    signal iNsTr_12_236 : std_logic_vector(31 downto 0);
    signal iNsTr_13_240 : std_logic_vector(31 downto 0);
    signal iNsTr_14_245 : std_logic_vector(31 downto 0);
    signal iNsTr_18_255 : std_logic_vector(31 downto 0);
    signal iNsTr_19_261 : std_logic_vector(31 downto 0);
    signal iNsTr_2_191 : std_logic_vector(31 downto 0);
    signal iNsTr_3_201 : std_logic_vector(0 downto 0);
    signal iNsTr_6_211 : std_logic_vector(31 downto 0);
    signal iNsTr_8_219 : std_logic_vector(31 downto 0);
    signal iNsTr_9_223 : std_logic_vector(31 downto 0);
    signal idx_176 : std_logic_vector(31 downto 0);
    signal ptr_deref_182_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_182_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_182_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_182_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_182_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_182_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_190_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_190_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_190_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_190_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_190_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_213_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_213_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_213_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_213_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_213_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_213_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_218_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_218_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_218_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_218_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_218_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_222_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_222_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_222_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_222_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_222_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_230_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_230_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_230_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_230_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_230_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_230_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_235_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_235_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_235_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_235_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_235_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_239_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_239_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_239_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_239_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_239_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_247_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_247_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_247_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_247_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_247_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_247_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_254_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_254_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_254_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_254_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_254_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_263_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_263_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_263_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_263_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_263_word_offset_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_225_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_225_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_242_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_242_scaled : std_logic_vector(6 downto 0);
    signal type_cast_184_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_195_wire : std_logic_vector(31 downto 0);
    signal type_cast_198_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_259_wire_constant : std_logic_vector(31 downto 0);
    signal val_180 : std_logic_vector(31 downto 0);
    signal xxgetDataxxbodyxxidx_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxgetDataxxbodyxxval_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_226_offset_scale_factor_0 <= "0000001";
    array_obj_ref_226_resized_base_address <= "0000000";
    array_obj_ref_243_offset_scale_factor_0 <= "0000001";
    array_obj_ref_243_resized_base_address <= "0000000";
    idx_176 <= "00000000000000000000000000000000";
    ptr_deref_182_word_offset_0 <= "0";
    ptr_deref_190_word_offset_0 <= "0";
    ptr_deref_213_word_offset_0 <= "0";
    ptr_deref_218_word_offset_0 <= "0";
    ptr_deref_222_word_offset_0 <= "0";
    ptr_deref_230_word_offset_0 <= "0000000";
    ptr_deref_235_word_offset_0 <= "0";
    ptr_deref_239_word_offset_0 <= "0";
    ptr_deref_247_word_offset_0 <= "0000000";
    ptr_deref_254_word_offset_0 <= "0";
    ptr_deref_263_word_offset_0 <= "0";
    type_cast_184_wire_constant <= "00000000000000000000000000000000";
    type_cast_198_wire_constant <= "00000000000000000000000001000000";
    type_cast_259_wire_constant <= "00000000000000000000000000000001";
    val_180 <= "00000000000000000000000000000000";
    xxgetDataxxbodyxxidx_alloc_base_address <= "0";
    xxgetDataxxbodyxxval_alloc_base_address <= "0";
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_227_final_reg_req_0,addr_of_227_final_reg_ack_0,sl_one,"addr_of_227_final_reg ",false,array_obj_ref_226_root_address,
    false,iNsTr_10_228);
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_227_final_reg_req_0;
      addr_of_227_final_reg_ack_0 <= ack; 
      addr_of_227_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_226_root_address, dout => iNsTr_10_228, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_244_final_reg_req_0,addr_of_244_final_reg_ack_0,sl_one,"addr_of_244_final_reg ",false,array_obj_ref_243_root_address,
    false,iNsTr_14_245);
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_244_final_reg_req_0;
      addr_of_244_final_reg_ack_0 <= ack; 
      addr_of_244_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_243_root_address, dout => iNsTr_14_245, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_195_inst_req_0,type_cast_195_inst_ack_0,sl_one,"type_cast_195_inst ",false,iNsTr_2_191,
    false,type_cast_195_wire);
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_195_inst_req_0;
      type_cast_195_inst_ack_0 <= ack; 
      type_cast_195_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_2_191, dout => type_cast_195_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_226_index_0_rename_req_0,array_obj_ref_226_index_0_rename_ack_0,sl_one,"array_obj_ref_226_index_0_rename ",false,simple_obj_ref_225_resized,
    false,simple_obj_ref_225_scaled);
    array_obj_ref_226_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_226_index_0_rename_ack_0 <= array_obj_ref_226_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_225_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_225_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_226_index_0_resize_req_0,array_obj_ref_226_index_0_resize_ack_0,sl_one,"array_obj_ref_226_index_0_resize ",false,iNsTr_9_223,
    false,simple_obj_ref_225_resized);
    array_obj_ref_226_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_226_index_0_resize_ack_0 <= array_obj_ref_226_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_9_223;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_225_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_226_offset_inst_req_0,array_obj_ref_226_offset_inst_ack_0,sl_one,"array_obj_ref_226_offset_inst ",false,simple_obj_ref_225_scaled,
    false,array_obj_ref_226_final_offset);
    array_obj_ref_226_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_226_offset_inst_ack_0 <= array_obj_ref_226_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_225_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_226_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_226_root_address_inst_req_0,array_obj_ref_226_root_address_inst_ack_0,sl_one,"array_obj_ref_226_root_address_inst ",false,array_obj_ref_226_final_offset,
    false,array_obj_ref_226_root_address);
    array_obj_ref_226_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_226_root_address_inst_ack_0 <= array_obj_ref_226_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_226_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_226_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_243_index_0_rename_req_0,array_obj_ref_243_index_0_rename_ack_0,sl_one,"array_obj_ref_243_index_0_rename ",false,simple_obj_ref_242_resized,
    false,simple_obj_ref_242_scaled);
    array_obj_ref_243_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_243_index_0_rename_ack_0 <= array_obj_ref_243_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_242_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_242_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_243_index_0_resize_req_0,array_obj_ref_243_index_0_resize_ack_0,sl_one,"array_obj_ref_243_index_0_resize ",false,iNsTr_13_240,
    false,simple_obj_ref_242_resized);
    array_obj_ref_243_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_243_index_0_resize_ack_0 <= array_obj_ref_243_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_13_240;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_242_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_243_offset_inst_req_0,array_obj_ref_243_offset_inst_ack_0,sl_one,"array_obj_ref_243_offset_inst ",false,simple_obj_ref_242_scaled,
    false,array_obj_ref_243_final_offset);
    array_obj_ref_243_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_243_offset_inst_ack_0 <= array_obj_ref_243_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_242_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_243_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_243_root_address_inst_req_0,array_obj_ref_243_root_address_inst_ack_0,sl_one,"array_obj_ref_243_root_address_inst ",false,array_obj_ref_243_final_offset,
    false,array_obj_ref_243_root_address);
    array_obj_ref_243_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_243_root_address_inst_ack_0 <= array_obj_ref_243_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_243_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_243_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_182_addr_0_req_0,ptr_deref_182_addr_0_ack_0,sl_one,"ptr_deref_182_addr_0 ",false,ptr_deref_182_root_address,
    false,ptr_deref_182_word_address_0);
    ptr_deref_182_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_182_addr_0_ack_0 <= ptr_deref_182_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_182_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_182_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_182_base_resize_req_0,ptr_deref_182_base_resize_ack_0,sl_one,"ptr_deref_182_base_resize ",false,idx_176,
    false,ptr_deref_182_resized_base_address);
    ptr_deref_182_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_182_base_resize_ack_0 <= ptr_deref_182_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_182_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_182_gather_scatter_req_0,ptr_deref_182_gather_scatter_ack_0,sl_one,"ptr_deref_182_gather_scatter ",false,type_cast_184_wire_constant,
    false,ptr_deref_182_data_0);
    ptr_deref_182_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_182_gather_scatter_ack_0 <= ptr_deref_182_gather_scatter_req_0;
      in_aggregated_sig <= type_cast_184_wire_constant;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_182_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_182_root_address_inst_req_0,ptr_deref_182_root_address_inst_ack_0,sl_one,"ptr_deref_182_root_address_inst ",false,ptr_deref_182_resized_base_address,
    false,ptr_deref_182_root_address);
    ptr_deref_182_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_182_root_address_inst_ack_0 <= ptr_deref_182_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_182_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_182_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_190_addr_0_req_0,ptr_deref_190_addr_0_ack_0,sl_one,"ptr_deref_190_addr_0 ",false,ptr_deref_190_root_address,
    false,ptr_deref_190_word_address_0);
    ptr_deref_190_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_190_addr_0_ack_0 <= ptr_deref_190_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_190_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_190_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_190_base_resize_req_0,ptr_deref_190_base_resize_ack_0,sl_one,"ptr_deref_190_base_resize ",false,idx_176,
    false,ptr_deref_190_resized_base_address);
    ptr_deref_190_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_190_base_resize_ack_0 <= ptr_deref_190_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_190_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_190_gather_scatter_req_0,ptr_deref_190_gather_scatter_ack_0,sl_one,"ptr_deref_190_gather_scatter ",false,ptr_deref_190_data_0,
    false,iNsTr_2_191);
    ptr_deref_190_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_190_gather_scatter_ack_0 <= ptr_deref_190_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_190_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_2_191 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_190_root_address_inst_req_0,ptr_deref_190_root_address_inst_ack_0,sl_one,"ptr_deref_190_root_address_inst ",false,ptr_deref_190_resized_base_address,
    false,ptr_deref_190_root_address);
    ptr_deref_190_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_190_root_address_inst_ack_0 <= ptr_deref_190_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_190_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_190_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_213_addr_0_req_0,ptr_deref_213_addr_0_ack_0,sl_one,"ptr_deref_213_addr_0 ",false,ptr_deref_213_root_address,
    false,ptr_deref_213_word_address_0);
    ptr_deref_213_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_213_addr_0_ack_0 <= ptr_deref_213_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_213_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_213_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_213_base_resize_req_0,ptr_deref_213_base_resize_ack_0,sl_one,"ptr_deref_213_base_resize ",false,val_180,
    false,ptr_deref_213_resized_base_address);
    ptr_deref_213_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_213_base_resize_ack_0 <= ptr_deref_213_base_resize_req_0;
      in_aggregated_sig <= val_180;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_213_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_213_gather_scatter_req_0,ptr_deref_213_gather_scatter_ack_0,sl_one,"ptr_deref_213_gather_scatter ",false,iNsTr_6_211,
    false,ptr_deref_213_data_0);
    ptr_deref_213_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_213_gather_scatter_ack_0 <= ptr_deref_213_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_6_211;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_213_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_213_root_address_inst_req_0,ptr_deref_213_root_address_inst_ack_0,sl_one,"ptr_deref_213_root_address_inst ",false,ptr_deref_213_resized_base_address,
    false,ptr_deref_213_root_address);
    ptr_deref_213_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_213_root_address_inst_ack_0 <= ptr_deref_213_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_213_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_213_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_218_addr_0_req_0,ptr_deref_218_addr_0_ack_0,sl_one,"ptr_deref_218_addr_0 ",false,ptr_deref_218_root_address,
    false,ptr_deref_218_word_address_0);
    ptr_deref_218_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_218_addr_0_ack_0 <= ptr_deref_218_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_218_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_218_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_218_base_resize_req_0,ptr_deref_218_base_resize_ack_0,sl_one,"ptr_deref_218_base_resize ",false,val_180,
    false,ptr_deref_218_resized_base_address);
    ptr_deref_218_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_218_base_resize_ack_0 <= ptr_deref_218_base_resize_req_0;
      in_aggregated_sig <= val_180;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_218_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_218_gather_scatter_req_0,ptr_deref_218_gather_scatter_ack_0,sl_one,"ptr_deref_218_gather_scatter ",false,ptr_deref_218_data_0,
    false,iNsTr_8_219);
    ptr_deref_218_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_218_gather_scatter_ack_0 <= ptr_deref_218_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_218_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_8_219 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_218_root_address_inst_req_0,ptr_deref_218_root_address_inst_ack_0,sl_one,"ptr_deref_218_root_address_inst ",false,ptr_deref_218_resized_base_address,
    false,ptr_deref_218_root_address);
    ptr_deref_218_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_218_root_address_inst_ack_0 <= ptr_deref_218_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_218_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_218_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_222_addr_0_req_0,ptr_deref_222_addr_0_ack_0,sl_one,"ptr_deref_222_addr_0 ",false,ptr_deref_222_root_address,
    false,ptr_deref_222_word_address_0);
    ptr_deref_222_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_222_addr_0_ack_0 <= ptr_deref_222_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_222_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_222_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_222_base_resize_req_0,ptr_deref_222_base_resize_ack_0,sl_one,"ptr_deref_222_base_resize ",false,idx_176,
    false,ptr_deref_222_resized_base_address);
    ptr_deref_222_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_222_base_resize_ack_0 <= ptr_deref_222_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_222_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_222_gather_scatter_req_0,ptr_deref_222_gather_scatter_ack_0,sl_one,"ptr_deref_222_gather_scatter ",false,ptr_deref_222_data_0,
    false,iNsTr_9_223);
    ptr_deref_222_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_222_gather_scatter_ack_0 <= ptr_deref_222_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_222_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_9_223 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_222_root_address_inst_req_0,ptr_deref_222_root_address_inst_ack_0,sl_one,"ptr_deref_222_root_address_inst ",false,ptr_deref_222_resized_base_address,
    false,ptr_deref_222_root_address);
    ptr_deref_222_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_222_root_address_inst_ack_0 <= ptr_deref_222_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_222_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_222_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_230_addr_0_req_0,ptr_deref_230_addr_0_ack_0,sl_one,"ptr_deref_230_addr_0 ",false,ptr_deref_230_root_address,
    false,ptr_deref_230_word_address_0);
    ptr_deref_230_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_230_addr_0_ack_0 <= ptr_deref_230_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_230_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_230_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_230_base_resize_req_0,ptr_deref_230_base_resize_ack_0,sl_one,"ptr_deref_230_base_resize ",false,iNsTr_10_228,
    false,ptr_deref_230_resized_base_address);
    ptr_deref_230_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_230_base_resize_ack_0 <= ptr_deref_230_base_resize_req_0;
      in_aggregated_sig <= iNsTr_10_228;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_230_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_230_gather_scatter_req_0,ptr_deref_230_gather_scatter_ack_0,sl_one,"ptr_deref_230_gather_scatter ",false,iNsTr_8_219,
    false,ptr_deref_230_data_0);
    ptr_deref_230_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_230_gather_scatter_ack_0 <= ptr_deref_230_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_8_219;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_230_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_230_root_address_inst_req_0,ptr_deref_230_root_address_inst_ack_0,sl_one,"ptr_deref_230_root_address_inst ",false,ptr_deref_230_resized_base_address,
    false,ptr_deref_230_root_address);
    ptr_deref_230_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_230_root_address_inst_ack_0 <= ptr_deref_230_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_230_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_230_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_235_addr_0_req_0,ptr_deref_235_addr_0_ack_0,sl_one,"ptr_deref_235_addr_0 ",false,ptr_deref_235_root_address,
    false,ptr_deref_235_word_address_0);
    ptr_deref_235_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_235_addr_0_ack_0 <= ptr_deref_235_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_235_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_235_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_235_base_resize_req_0,ptr_deref_235_base_resize_ack_0,sl_one,"ptr_deref_235_base_resize ",false,val_180,
    false,ptr_deref_235_resized_base_address);
    ptr_deref_235_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_235_base_resize_ack_0 <= ptr_deref_235_base_resize_req_0;
      in_aggregated_sig <= val_180;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_235_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_235_gather_scatter_req_0,ptr_deref_235_gather_scatter_ack_0,sl_one,"ptr_deref_235_gather_scatter ",false,ptr_deref_235_data_0,
    false,iNsTr_12_236);
    ptr_deref_235_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_235_gather_scatter_ack_0 <= ptr_deref_235_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_235_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_12_236 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_235_root_address_inst_req_0,ptr_deref_235_root_address_inst_ack_0,sl_one,"ptr_deref_235_root_address_inst ",false,ptr_deref_235_resized_base_address,
    false,ptr_deref_235_root_address);
    ptr_deref_235_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_235_root_address_inst_ack_0 <= ptr_deref_235_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_235_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_235_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_239_addr_0_req_0,ptr_deref_239_addr_0_ack_0,sl_one,"ptr_deref_239_addr_0 ",false,ptr_deref_239_root_address,
    false,ptr_deref_239_word_address_0);
    ptr_deref_239_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_239_addr_0_ack_0 <= ptr_deref_239_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_239_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_239_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_239_base_resize_req_0,ptr_deref_239_base_resize_ack_0,sl_one,"ptr_deref_239_base_resize ",false,idx_176,
    false,ptr_deref_239_resized_base_address);
    ptr_deref_239_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_239_base_resize_ack_0 <= ptr_deref_239_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_239_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_239_gather_scatter_req_0,ptr_deref_239_gather_scatter_ack_0,sl_one,"ptr_deref_239_gather_scatter ",false,ptr_deref_239_data_0,
    false,iNsTr_13_240);
    ptr_deref_239_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_239_gather_scatter_ack_0 <= ptr_deref_239_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_239_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_13_240 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_239_root_address_inst_req_0,ptr_deref_239_root_address_inst_ack_0,sl_one,"ptr_deref_239_root_address_inst ",false,ptr_deref_239_resized_base_address,
    false,ptr_deref_239_root_address);
    ptr_deref_239_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_239_root_address_inst_ack_0 <= ptr_deref_239_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_239_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_239_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_247_addr_0_req_0,ptr_deref_247_addr_0_ack_0,sl_one,"ptr_deref_247_addr_0 ",false,ptr_deref_247_root_address,
    false,ptr_deref_247_word_address_0);
    ptr_deref_247_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_247_addr_0_ack_0 <= ptr_deref_247_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_247_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_247_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_247_base_resize_req_0,ptr_deref_247_base_resize_ack_0,sl_one,"ptr_deref_247_base_resize ",false,iNsTr_14_245,
    false,ptr_deref_247_resized_base_address);
    ptr_deref_247_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_247_base_resize_ack_0 <= ptr_deref_247_base_resize_req_0;
      in_aggregated_sig <= iNsTr_14_245;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_247_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_247_gather_scatter_req_0,ptr_deref_247_gather_scatter_ack_0,sl_one,"ptr_deref_247_gather_scatter ",false,iNsTr_12_236,
    false,ptr_deref_247_data_0);
    ptr_deref_247_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_247_gather_scatter_ack_0 <= ptr_deref_247_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_12_236;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_247_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_247_root_address_inst_req_0,ptr_deref_247_root_address_inst_ack_0,sl_one,"ptr_deref_247_root_address_inst ",false,ptr_deref_247_resized_base_address,
    false,ptr_deref_247_root_address);
    ptr_deref_247_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_247_root_address_inst_ack_0 <= ptr_deref_247_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_247_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_247_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_254_addr_0_req_0,ptr_deref_254_addr_0_ack_0,sl_one,"ptr_deref_254_addr_0 ",false,ptr_deref_254_root_address,
    false,ptr_deref_254_word_address_0);
    ptr_deref_254_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_254_addr_0_ack_0 <= ptr_deref_254_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_254_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_254_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_254_base_resize_req_0,ptr_deref_254_base_resize_ack_0,sl_one,"ptr_deref_254_base_resize ",false,idx_176,
    false,ptr_deref_254_resized_base_address);
    ptr_deref_254_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_254_base_resize_ack_0 <= ptr_deref_254_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_254_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_254_gather_scatter_req_0,ptr_deref_254_gather_scatter_ack_0,sl_one,"ptr_deref_254_gather_scatter ",false,ptr_deref_254_data_0,
    false,iNsTr_18_255);
    ptr_deref_254_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_254_gather_scatter_ack_0 <= ptr_deref_254_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_254_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_18_255 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_254_root_address_inst_req_0,ptr_deref_254_root_address_inst_ack_0,sl_one,"ptr_deref_254_root_address_inst ",false,ptr_deref_254_resized_base_address,
    false,ptr_deref_254_root_address);
    ptr_deref_254_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_254_root_address_inst_ack_0 <= ptr_deref_254_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_254_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_254_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_263_addr_0_req_0,ptr_deref_263_addr_0_ack_0,sl_one,"ptr_deref_263_addr_0 ",false,ptr_deref_263_root_address,
    false,ptr_deref_263_word_address_0);
    ptr_deref_263_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_263_addr_0_ack_0 <= ptr_deref_263_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_263_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_263_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_263_base_resize_req_0,ptr_deref_263_base_resize_ack_0,sl_one,"ptr_deref_263_base_resize ",false,idx_176,
    false,ptr_deref_263_resized_base_address);
    ptr_deref_263_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_263_base_resize_ack_0 <= ptr_deref_263_base_resize_req_0;
      in_aggregated_sig <= idx_176;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_263_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_263_gather_scatter_req_0,ptr_deref_263_gather_scatter_ack_0,sl_one,"ptr_deref_263_gather_scatter ",false,iNsTr_19_261,
    false,ptr_deref_263_data_0);
    ptr_deref_263_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_263_gather_scatter_ack_0 <= ptr_deref_263_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_19_261;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_263_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_263_root_address_inst_req_0,ptr_deref_263_root_address_inst_ack_0,sl_one,"ptr_deref_263_root_address_inst ",false,ptr_deref_263_resized_base_address,
    false,ptr_deref_263_root_address);
    ptr_deref_263_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_263_root_address_inst_ack_0 <= ptr_deref_263_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_263_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_263_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_202_branch_req_0," req0 if_stmt_202_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_202_branch_ack_0," ack0 if_stmt_202_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_202_branch_ack_1," ack1 if_stmt_202_branch");
    if_stmt_202_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_201;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_202_branch_req_0,
          ack0 => if_stmt_202_branch_ack_0,
          ack1 => if_stmt_202_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_199_inst_req_0,binary_199_inst_ack_0,binary_199_inst_req_1,binary_199_inst_ack_1,sl_one,"binary_199_inst",false,type_cast_195_wire & type_cast_198_wire_constant,
    false,iNsTr_3_201);
    -- shared split operator group (0) : binary_199_inst 
    ApIntSlt_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_195_wire;
      iNsTr_3_201 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_199_inst_req_0;
      reqR(0) <= binary_199_inst_req_1;
      binary_199_inst_ack_0 <= ackL(0); 
      binary_199_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_260_inst_req_0,binary_260_inst_ack_0,binary_260_inst_req_1,binary_260_inst_ack_1,sl_one,"binary_260_inst",false,iNsTr_18_255 & type_cast_259_wire_constant,
    false,iNsTr_19_261);
    -- shared split operator group (1) : binary_260_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_18_255;
      iNsTr_19_261 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_260_inst_req_0;
      reqR(0) <= binary_260_inst_req_1;
      binary_260_inst_ack_0 <= ackL(0); 
      binary_260_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_190_load_0_req_0,ptr_deref_190_load_0_ack_0,ptr_deref_190_load_0_req_1,ptr_deref_190_load_0_ack_1,sl_one,"ptr_deref_190_load_0",false,ptr_deref_190_word_address_0,
    false,ptr_deref_190_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_222_load_0_req_0,ptr_deref_222_load_0_ack_0,ptr_deref_222_load_0_req_1,ptr_deref_222_load_0_ack_1,sl_one,"ptr_deref_222_load_0",false,ptr_deref_222_word_address_0,
    false,ptr_deref_222_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_254_load_0_req_0,ptr_deref_254_load_0_ack_0,ptr_deref_254_load_0_req_1,ptr_deref_254_load_0_ack_1,sl_one,"ptr_deref_254_load_0",false,ptr_deref_254_word_address_0,
    false,ptr_deref_254_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_239_load_0_req_0,ptr_deref_239_load_0_ack_0,ptr_deref_239_load_0_req_1,ptr_deref_239_load_0_ack_1,sl_one,"ptr_deref_239_load_0",false,ptr_deref_239_word_address_0,
    false,ptr_deref_239_data_0);
    -- shared load operator group (0) : ptr_deref_190_load_0 ptr_deref_222_load_0 ptr_deref_254_load_0 ptr_deref_239_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(3 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_190_load_0_req_0,
        ptr_deref_190_load_0_ack_0,
        ptr_deref_190_load_0_req_1,
        ptr_deref_190_load_0_ack_1,
        "ptr_deref_190_load_0",
        "memory_space_3" ,
        ptr_deref_190_data_0,
        ptr_deref_190_word_address_0,
        "ptr_deref_190_data_0",
        "ptr_deref_190_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_222_load_0_req_0,
        ptr_deref_222_load_0_ack_0,
        ptr_deref_222_load_0_req_1,
        ptr_deref_222_load_0_ack_1,
        "ptr_deref_222_load_0",
        "memory_space_3" ,
        ptr_deref_222_data_0,
        ptr_deref_222_word_address_0,
        "ptr_deref_222_data_0",
        "ptr_deref_222_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_254_load_0_req_0,
        ptr_deref_254_load_0_ack_0,
        ptr_deref_254_load_0_req_1,
        ptr_deref_254_load_0_ack_1,
        "ptr_deref_254_load_0",
        "memory_space_3" ,
        ptr_deref_254_data_0,
        ptr_deref_254_word_address_0,
        "ptr_deref_254_data_0",
        "ptr_deref_254_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_239_load_0_req_0,
        ptr_deref_239_load_0_ack_0,
        ptr_deref_239_load_0_req_1,
        ptr_deref_239_load_0_ack_1,
        "ptr_deref_239_load_0",
        "memory_space_3" ,
        ptr_deref_239_data_0,
        ptr_deref_239_word_address_0,
        "ptr_deref_239_data_0",
        "ptr_deref_239_word_address_0" -- 
      );
      reqL_unguarded(3) <= ptr_deref_190_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_222_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_254_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_239_load_0_req_0;
      ptr_deref_190_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_222_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_254_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_239_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= ptr_deref_190_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_222_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_254_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_239_load_0_req_1;
      ptr_deref_190_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_222_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_254_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_239_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 4) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 4) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_190_word_address_0 & ptr_deref_222_word_address_0 & ptr_deref_254_word_address_0 & ptr_deref_239_word_address_0;
      ptr_deref_190_data_0 <= data_out(127 downto 96);
      ptr_deref_222_data_0 <= data_out(95 downto 64);
      ptr_deref_254_data_0 <= data_out(63 downto 32);
      ptr_deref_239_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(0 downto 0),
          mtag => memory_space_3_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 4,  tag_length => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(31 downto 0),
          mtag => memory_space_3_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_235_load_0_req_0,ptr_deref_235_load_0_ack_0,ptr_deref_235_load_0_req_1,ptr_deref_235_load_0_ack_1,sl_one,"ptr_deref_235_load_0",false,ptr_deref_235_word_address_0,
    false,ptr_deref_235_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_218_load_0_req_0,ptr_deref_218_load_0_ack_0,ptr_deref_218_load_0_req_1,ptr_deref_218_load_0_ack_1,sl_one,"ptr_deref_218_load_0",false,ptr_deref_218_word_address_0,
    false,ptr_deref_218_data_0);
    -- shared load operator group (1) : ptr_deref_235_load_0 ptr_deref_218_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_235_load_0_req_0,
        ptr_deref_235_load_0_ack_0,
        ptr_deref_235_load_0_req_1,
        ptr_deref_235_load_0_ack_1,
        "ptr_deref_235_load_0",
        "memory_space_4" ,
        ptr_deref_235_data_0,
        ptr_deref_235_word_address_0,
        "ptr_deref_235_data_0",
        "ptr_deref_235_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_218_load_0_req_0,
        ptr_deref_218_load_0_ack_0,
        ptr_deref_218_load_0_req_1,
        ptr_deref_218_load_0_ack_1,
        "ptr_deref_218_load_0",
        "memory_space_4" ,
        ptr_deref_218_data_0,
        ptr_deref_218_word_address_0,
        "ptr_deref_218_data_0",
        "ptr_deref_218_word_address_0" -- 
      );
      reqL_unguarded(1) <= ptr_deref_235_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_218_load_0_req_0;
      ptr_deref_235_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_218_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_235_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_218_load_0_req_1;
      ptr_deref_235_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_218_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_235_word_address_0 & ptr_deref_218_word_address_0;
      ptr_deref_235_data_0 <= data_out(63 downto 32);
      ptr_deref_218_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 2,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_182_store_0_req_0,ptr_deref_182_store_0_ack_0,ptr_deref_182_store_0_req_1,ptr_deref_182_store_0_ack_1,sl_one,"ptr_deref_182_store_0",false,ptr_deref_182_word_address_0 & ptr_deref_182_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_263_store_0_req_0,ptr_deref_263_store_0_ack_0,ptr_deref_263_store_0_req_1,ptr_deref_263_store_0_ack_1,sl_one,"ptr_deref_263_store_0",false,ptr_deref_263_word_address_0 & ptr_deref_263_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_182_store_0_req_0,
      ptr_deref_182_store_0_ack_0,
      ptr_deref_182_store_0_req_1,
      ptr_deref_182_store_0_ack_1,
      "ptr_deref_182_store_0",
      "memory_space_3" ,
      ptr_deref_182_data_0,
      ptr_deref_182_word_address_0,
      "ptr_deref_182_data_0",
      "ptr_deref_182_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_263_store_0_req_0,
      ptr_deref_263_store_0_ack_0,
      ptr_deref_263_store_0_req_1,
      ptr_deref_263_store_0_ack_1,
      "ptr_deref_263_store_0",
      "memory_space_3" ,
      ptr_deref_263_data_0,
      ptr_deref_263_word_address_0,
      "ptr_deref_263_data_0",
      "ptr_deref_263_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_182_store_0 ptr_deref_263_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_182_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_263_store_0_req_0;
      ptr_deref_182_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_263_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_182_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_263_store_0_req_1;
      ptr_deref_182_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_263_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_182_word_address_0 & ptr_deref_263_word_address_0;
      data_in <= ptr_deref_182_data_0 & ptr_deref_263_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(0 downto 0),
          mdata => memory_space_3_sr_data(31 downto 0),
          mtag => memory_space_3_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_213_store_0_req_0,ptr_deref_213_store_0_ack_0,ptr_deref_213_store_0_req_1,ptr_deref_213_store_0_ack_1,sl_one,"ptr_deref_213_store_0",false,ptr_deref_213_word_address_0 & ptr_deref_213_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_213_store_0_req_0,
      ptr_deref_213_store_0_ack_0,
      ptr_deref_213_store_0_req_1,
      ptr_deref_213_store_0_ack_1,
      "ptr_deref_213_store_0",
      "memory_space_4" ,
      ptr_deref_213_data_0,
      ptr_deref_213_word_address_0,
      "ptr_deref_213_data_0",
      "ptr_deref_213_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_213_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_213_store_0_req_0;
      ptr_deref_213_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_213_store_0_req_1;
      ptr_deref_213_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_213_word_address_0;
      data_in <= ptr_deref_213_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_230_store_0_req_0,ptr_deref_230_store_0_ack_0,ptr_deref_230_store_0_req_1,ptr_deref_230_store_0_ack_1,sl_one,"ptr_deref_230_store_0",false,ptr_deref_230_word_address_0 & ptr_deref_230_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_230_store_0_req_0,
      ptr_deref_230_store_0_ack_0,
      ptr_deref_230_store_0_req_1,
      ptr_deref_230_store_0_ack_1,
      "ptr_deref_230_store_0",
      "memory_space_0" ,
      ptr_deref_230_data_0,
      ptr_deref_230_word_address_0,
      "ptr_deref_230_data_0",
      "ptr_deref_230_word_address_0" -- 
    );
    -- shared store operator group (2) : ptr_deref_230_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(6 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_230_store_0_req_0;
      ptr_deref_230_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_230_store_0_req_1;
      ptr_deref_230_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_230_word_address_0;
      data_in <= ptr_deref_230_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_247_store_0_req_0,ptr_deref_247_store_0_ack_0,ptr_deref_247_store_0_req_1,ptr_deref_247_store_0_ack_1,sl_one,"ptr_deref_247_store_0",false,ptr_deref_247_word_address_0 & ptr_deref_247_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_247_store_0_req_0,
      ptr_deref_247_store_0_ack_0,
      ptr_deref_247_store_0_req_1,
      ptr_deref_247_store_0_ack_1,
      "ptr_deref_247_store_0",
      "memory_space_1" ,
      ptr_deref_247_data_0,
      ptr_deref_247_word_address_0,
      "ptr_deref_247_data_0",
      "ptr_deref_247_word_address_0" -- 
    );
    -- shared store operator group (3) : ptr_deref_247_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(6 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_247_store_0_req_0;
      ptr_deref_247_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_247_store_0_req_1;
      ptr_deref_247_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_247_word_address_0;
      data_in <= ptr_deref_247_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_210_inst_req_0,simple_obj_ref_210_inst_ack_0,sl_one,"simple_obj_ref_210_inst  PipeRead from in_data_pipe",true, slv_zero,
    false,iNsTr_6_211);
    -- shared inport operator group (0) : simple_obj_ref_210_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_210_inst_ack_0 then -- 
            assert false report " ReadPipe in_data_pipe to wire iNsTr_6_211 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req_unguarded(0) <= simple_obj_ref_210_inst_req_0;
      simple_obj_ref_210_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      iNsTr_6_211 <= data_out(31 downto 0);
      in_data_pipe_read_0: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_pipe_read_req(0),
          oack => in_data_pipe_pipe_read_ack(0),
          odata => in_data_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity sendResult is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    out_data_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity sendResult;
architecture Default of sendResult is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal sendResult_CP_1524_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_293_store_0_req_0 : boolean;
  signal ptr_deref_293_store_0_ack_0 : boolean;
  signal ptr_deref_293_root_address_inst_req_0 : boolean;
  signal ptr_deref_301_root_address_inst_ack_0 : boolean;
  signal ptr_deref_301_addr_0_req_0 : boolean;
  signal ptr_deref_293_addr_0_req_0 : boolean;
  signal ptr_deref_301_load_0_req_0 : boolean;
  signal ptr_deref_301_load_0_ack_0 : boolean;
  signal ptr_deref_293_store_0_req_1 : boolean;
  signal ptr_deref_293_gather_scatter_ack_0 : boolean;
  signal ptr_deref_293_store_0_ack_1 : boolean;
  signal ptr_deref_293_gather_scatter_req_0 : boolean;
  signal ptr_deref_293_addr_0_ack_0 : boolean;
  signal ptr_deref_293_base_resize_ack_0 : boolean;
  signal ptr_deref_293_base_resize_req_0 : boolean;
  signal ptr_deref_301_base_resize_req_0 : boolean;
  signal ptr_deref_301_addr_0_ack_0 : boolean;
  signal ptr_deref_293_root_address_inst_ack_0 : boolean;
  signal ptr_deref_301_root_address_inst_req_0 : boolean;
  signal ptr_deref_301_base_resize_ack_0 : boolean;
  signal ptr_deref_301_load_0_req_1 : boolean;
  signal ptr_deref_301_load_0_ack_1 : boolean;
  signal ptr_deref_301_gather_scatter_req_0 : boolean;
  signal ptr_deref_301_gather_scatter_ack_0 : boolean;
  signal type_cast_305_inst_req_0 : boolean;
  signal type_cast_305_inst_ack_0 : boolean;
  signal binary_309_inst_req_0 : boolean;
  signal binary_309_inst_ack_0 : boolean;
  signal binary_309_inst_req_1 : boolean;
  signal binary_309_inst_ack_1 : boolean;
  signal if_stmt_311_branch_req_0 : boolean;
  signal if_stmt_311_branch_ack_1 : boolean;
  signal if_stmt_311_branch_ack_0 : boolean;
  signal ptr_deref_320_base_resize_req_0 : boolean;
  signal ptr_deref_320_base_resize_ack_0 : boolean;
  signal ptr_deref_320_root_address_inst_req_0 : boolean;
  signal ptr_deref_320_root_address_inst_ack_0 : boolean;
  signal ptr_deref_320_addr_0_req_0 : boolean;
  signal ptr_deref_320_addr_0_ack_0 : boolean;
  signal ptr_deref_320_load_0_req_0 : boolean;
  signal ptr_deref_320_load_0_ack_0 : boolean;
  signal ptr_deref_320_load_0_req_1 : boolean;
  signal ptr_deref_320_load_0_ack_1 : boolean;
  signal ptr_deref_320_gather_scatter_req_0 : boolean;
  signal ptr_deref_320_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_324_index_0_resize_req_0 : boolean;
  signal array_obj_ref_324_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_324_index_0_rename_req_0 : boolean;
  signal array_obj_ref_324_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_324_offset_inst_req_0 : boolean;
  signal array_obj_ref_324_offset_inst_ack_0 : boolean;
  signal array_obj_ref_324_root_address_inst_req_0 : boolean;
  signal array_obj_ref_324_root_address_inst_ack_0 : boolean;
  signal addr_of_325_final_reg_req_0 : boolean;
  signal addr_of_325_final_reg_ack_0 : boolean;
  signal ptr_deref_329_base_resize_req_0 : boolean;
  signal ptr_deref_329_base_resize_ack_0 : boolean;
  signal ptr_deref_329_root_address_inst_req_0 : boolean;
  signal ptr_deref_329_root_address_inst_ack_0 : boolean;
  signal ptr_deref_329_addr_0_req_0 : boolean;
  signal ptr_deref_329_addr_0_ack_0 : boolean;
  signal ptr_deref_329_load_0_req_0 : boolean;
  signal ptr_deref_329_load_0_ack_0 : boolean;
  signal ptr_deref_329_load_0_req_1 : boolean;
  signal ptr_deref_329_load_0_ack_1 : boolean;
  signal ptr_deref_329_gather_scatter_req_0 : boolean;
  signal ptr_deref_329_gather_scatter_ack_0 : boolean;
  signal ptr_deref_332_base_resize_req_0 : boolean;
  signal ptr_deref_332_base_resize_ack_0 : boolean;
  signal ptr_deref_332_root_address_inst_req_0 : boolean;
  signal ptr_deref_332_root_address_inst_ack_0 : boolean;
  signal ptr_deref_332_addr_0_req_0 : boolean;
  signal ptr_deref_332_addr_0_ack_0 : boolean;
  signal ptr_deref_332_gather_scatter_req_0 : boolean;
  signal ptr_deref_332_gather_scatter_ack_0 : boolean;
  signal ptr_deref_332_store_0_req_0 : boolean;
  signal ptr_deref_332_store_0_ack_0 : boolean;
  signal ptr_deref_332_store_0_req_1 : boolean;
  signal ptr_deref_332_store_0_ack_1 : boolean;
  signal ptr_deref_337_base_resize_req_0 : boolean;
  signal ptr_deref_337_base_resize_ack_0 : boolean;
  signal ptr_deref_337_root_address_inst_req_0 : boolean;
  signal ptr_deref_337_root_address_inst_ack_0 : boolean;
  signal ptr_deref_337_addr_0_req_0 : boolean;
  signal ptr_deref_337_addr_0_ack_0 : boolean;
  signal ptr_deref_337_load_0_req_0 : boolean;
  signal ptr_deref_337_load_0_ack_0 : boolean;
  signal ptr_deref_337_load_0_req_1 : boolean;
  signal ptr_deref_337_load_0_ack_1 : boolean;
  signal ptr_deref_337_gather_scatter_req_0 : boolean;
  signal ptr_deref_337_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_339_inst_req_0 : boolean;
  signal simple_obj_ref_339_inst_ack_0 : boolean;
  signal ptr_deref_346_base_resize_req_0 : boolean;
  signal ptr_deref_346_base_resize_ack_0 : boolean;
  signal ptr_deref_346_root_address_inst_req_0 : boolean;
  signal ptr_deref_346_root_address_inst_ack_0 : boolean;
  signal ptr_deref_346_addr_0_req_0 : boolean;
  signal ptr_deref_346_addr_0_ack_0 : boolean;
  signal ptr_deref_346_load_0_req_0 : boolean;
  signal ptr_deref_346_load_0_ack_0 : boolean;
  signal ptr_deref_346_load_0_req_1 : boolean;
  signal ptr_deref_346_load_0_ack_1 : boolean;
  signal ptr_deref_346_gather_scatter_req_0 : boolean;
  signal ptr_deref_346_gather_scatter_ack_0 : boolean;
  signal binary_352_inst_req_0 : boolean;
  signal binary_352_inst_ack_0 : boolean;
  signal binary_352_inst_req_1 : boolean;
  signal binary_352_inst_ack_1 : boolean;
  signal ptr_deref_355_base_resize_req_0 : boolean;
  signal ptr_deref_355_base_resize_ack_0 : boolean;
  signal ptr_deref_355_root_address_inst_req_0 : boolean;
  signal ptr_deref_355_root_address_inst_ack_0 : boolean;
  signal ptr_deref_355_addr_0_req_0 : boolean;
  signal ptr_deref_355_addr_0_ack_0 : boolean;
  signal ptr_deref_355_gather_scatter_req_0 : boolean;
  signal ptr_deref_355_gather_scatter_ack_0 : boolean;
  signal ptr_deref_355_store_0_req_0 : boolean;
  signal ptr_deref_355_store_0_ack_0 : boolean;
  signal ptr_deref_355_store_0_req_1 : boolean;
  signal ptr_deref_355_store_0_ack_1 : boolean;
  signal memory_space_5_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(0 downto 0);
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"sendResult start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"sendResult start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"sendResult fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"sendResult fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  sendResult_CP_1524: Block -- control-path 
    signal cp_elements: BooleanArray(106 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(39);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(39), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 5 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296__entry__
      -- 	branch_block_stmt_281/branch_block_stmt_281__entry__
      -- 	branch_block_stmt_281/$entry
      -- 	$entry
      -- 
    -- CP-element group 1 branch  place  bypass 
    -- predecessors 30 
    -- successors 31 34 
    -- members (2) 
      -- 	branch_block_stmt_281/if_stmt_311__entry__
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310__exit__
      -- 
    cp_elements(1) <= cp_elements(30);
    -- CP-element group 2 merge  place  bypass 
    -- predecessors 37 106 
    -- successors 40 
    -- members (2) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338__entry__
      -- 	branch_block_stmt_281/merge_stmt_317__exit__
      -- 
    cp_elements(2) <= OrReduce(cp_elements(37) & cp_elements(106));
    -- CP-element group 3 transition  place  output  bypass 
    -- predecessors 78 
    -- successors 79 
    -- members (11) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338__exit__
      -- 	branch_block_stmt_281/assign_stmt_341__entry__
      -- 	branch_block_stmt_281/assign_stmt_341/$entry
      -- 	branch_block_stmt_281/assign_stmt_341/assign_stmt_341_trigger_
      -- 	branch_block_stmt_281/assign_stmt_341/assign_stmt_341_active_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_340_trigger_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_340_active_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_340_completed_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_trigger_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_complete/pipe_wreq
      -- 
    cp_elements(3) <= cp_elements(78);
    pipe_wreq_1982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_339_inst_req_0); -- 
    -- CP-element group 4 transition  place  bypass 
    -- predecessors 102 
    -- successors 103 
    -- members (4) 
      -- 	branch_block_stmt_281/bb_3_bb_1
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357__exit__
      -- 	branch_block_stmt_281/bb_3_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_281/bb_3_bb_1_PhiReq/$exit
      -- 
    cp_elements(4) <= cp_elements(102);
    -- CP-element group 5 fork  transition  bypass 
    -- predecessors 0 
    -- successors 6 8 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/$entry
      -- 
    cp_elements(5) <= cp_elements(0);
    -- CP-element group 6 transition  bypass 
    -- predecessors 5 
    -- successors 7 
    -- members (2) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/assign_stmt_296_active_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/assign_stmt_296_trigger_
      -- 
    cp_elements(6) <= cp_elements(5);
    -- CP-element group 7 join  transition  output  no-bypass 
    -- predecessors 6 11 
    -- successors 12 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_trigger_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/split_req
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/$entry
      -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(6);
      predecessors(1) <= cp_elements(11);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(7)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_1588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_293_gather_scatter_req_0); -- 
    -- CP-element group 8 transition  output  bypass 
    -- predecessors 5 
    -- successors 9 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/simple_obj_ref_292_trigger_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/simple_obj_ref_292_completed_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/simple_obj_ref_292_active_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_addr_resize/$entry
      -- 
    cp_elements(8) <= cp_elements(5);
    base_resize_req_1573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => ptr_deref_293_base_resize_req_0); -- 
    -- CP-element group 9 transition  input  output  no-bypass 
    -- predecessors 8 
    -- successors 10 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_addr_resize/$exit
      -- 
    base_resize_ack_1574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_base_resize_ack_0, ack => cp_elements(9)); -- 
    sum_rename_req_1578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => ptr_deref_293_root_address_inst_req_0); -- 
    -- CP-element group 10 transition  input  output  no-bypass 
    -- predecessors 9 
    -- successors 11 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_word_addrgen/root_register_req
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_root_address_inst_ack_0, ack => cp_elements(10)); -- 
    root_register_req_1583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_293_addr_0_req_0); -- 
    -- CP-element group 11 transition  input  no-bypass 
    -- predecessors 10 
    -- successors 7 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_word_addrgen/root_register_ack
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_word_address_calculated
      -- 
    root_register_ack_1584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_addr_0_ack_0, ack => cp_elements(11)); -- 
    -- CP-element group 12 transition  input  output  no-bypass 
    -- predecessors 7 
    -- successors 13 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/split_ack
      -- 
    split_ack_1589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_gather_scatter_ack_0, ack => cp_elements(12)); -- 
    rr_1596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => ptr_deref_293_store_0_req_0); -- 
    -- CP-element group 13 transition  input  output  no-bypass 
    -- predecessors 12 
    -- successors 14 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_active_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/$entry
      -- 
    ra_1597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_store_0_ack_0, ack => cp_elements(13)); -- 
    cr_1607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_293_store_0_req_1); -- 
    -- CP-element group 14 transition  place  input  no-bypass 
    -- predecessors 13 
    -- successors 103 
    -- members (11) 
      -- 	branch_block_stmt_281/bb_0_bb_1
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_completed_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296__exit__
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/assign_stmt_296_completed_
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/$exit
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_287_to_assign_stmt_296/ptr_deref_293_complete/$exit
      -- 	branch_block_stmt_281/bb_0_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_281/bb_0_bb_1_PhiReq/$exit
      -- 
    ca_1608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_293_store_0_ack_1, ack => cp_elements(14)); -- 
    -- CP-element group 15 fork  transition  bypass 
    -- predecessors 104 
    -- successors 16 23 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/$entry
      -- 
    cp_elements(15) <= cp_elements(104);
    -- CP-element group 16 transition  output  bypass 
    -- predecessors 15 
    -- successors 17 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_300_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_300_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_300_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_address_calculated
      -- 
    cp_elements(16) <= cp_elements(15);
    base_resize_req_1628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_301_base_resize_req_0); -- 
    -- CP-element group 17 transition  input  output  no-bypass 
    -- predecessors 16 
    -- successors 18 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_1629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_base_resize_ack_0, ack => cp_elements(17)); -- 
    sum_rename_req_1633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_301_root_address_inst_req_0); -- 
    -- CP-element group 18 transition  input  output  no-bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_word_addrgen/root_register_req
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_base_plus_offset/$exit
      -- 
    sum_rename_ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_root_address_inst_ack_0, ack => cp_elements(18)); -- 
    root_register_req_1638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_301_addr_0_req_0); -- 
    -- CP-element group 19 transition  input  output  no-bypass 
    -- predecessors 18 
    -- successors 20 
    -- members (8) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_word_addrgen/root_register_ack
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/$entry
      -- 
    root_register_ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_addr_0_ack_0, ack => cp_elements(19)); -- 
    rr_1649_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_301_load_0_req_0); -- 
    -- CP-element group 20 transition  input  output  no-bypass 
    -- predecessors 19 
    -- successors 21 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/word_access_0/cr
      -- 
    ra_1650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_load_0_ack_0, ack => cp_elements(20)); -- 
    cr_1660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_301_load_0_req_1); -- 
    -- CP-element group 21 transition  input  output  no-bypass 
    -- predecessors 20 
    -- successors 22 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/merge_req
      -- 
    ca_1661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_load_0_ack_1, ack => cp_elements(21)); -- 
    merge_req_1662_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_301_gather_scatter_req_0); -- 
    -- CP-element group 22 transition  input  output  no-bypass 
    -- predecessors 21 
    -- successors 27 
    -- members (12) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_302_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_302_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_302_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/ptr_deref_301_complete/merge_ack
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_304_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_304_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/simple_obj_ref_304_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_complete/req
      -- 
    merge_ack_1663_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_301_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    req_1683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => type_cast_305_inst_req_0); -- 
    -- CP-element group 23 transition  bypass 
    -- predecessors 15 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_active_
      -- 
    cp_elements(23) <= cp_elements(15);
    -- CP-element group 24 join  transition  bypass 
    -- predecessors 28 29 
    -- successors 30 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_310_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_310_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/assign_stmt_310_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_completed_
      -- 
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(28);
      predecessors(1) <= cp_elements(29);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(24)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 25 transition  output  bypass 
    -- predecessors 27 
    -- successors 28 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_sample_start_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Sample/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Sample/rr
      -- 
    cp_elements(25) <= cp_elements(27);
    rr_1688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => binary_309_inst_req_0); -- 
    -- CP-element group 26 transition  output  bypass 
    -- predecessors 27 
    -- successors 29 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_update_start_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Update/$entry
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Update/cr
      -- 
    cp_elements(26) <= cp_elements(27);
    cr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_309_inst_req_1); -- 
    -- CP-element group 27 fork  transition  input  no-bypass 
    -- predecessors 22 
    -- successors 25 26 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_trigger_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_active_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/type_cast_305_complete/ack
      -- 
    ack_1684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_305_inst_ack_0, ack => cp_elements(27)); -- 
    -- CP-element group 28 transition  input  no-bypass 
    -- predecessors 25 
    -- successors 24 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_sample_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Sample/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Sample/ra
      -- 
    ra_1689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_309_inst_ack_0, ack => cp_elements(28)); -- 
    -- CP-element group 29 transition  input  no-bypass 
    -- predecessors 26 
    -- successors 24 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_update_completed_
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Update/$exit
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/binary_309_Update/ca
      -- 
    ca_1694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_309_inst_ack_1, ack => cp_elements(29)); -- 
    -- CP-element group 30 join  transition  no-bypass 
    -- predecessors 23 24 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310/$exit
      -- 
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(23);
      predecessors(1) <= cp_elements(24);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(30)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 31 transition  bypass 
    -- predecessors 1 
    -- successors 32 
    -- members (1) 
      -- 	branch_block_stmt_281/if_stmt_311_dead_link/$entry
      -- 
    cp_elements(31) <= cp_elements(1);
    -- CP-element group 32 transition  dead  bypass 
    -- predecessors 31 
    -- successors 33 
    -- members (1) 
      -- 	branch_block_stmt_281/if_stmt_311_dead_link/dead_transition
      -- 
    cp_elements(32) <= false;
    -- CP-element group 33 transition  place  bypass 
    -- predecessors 32 
    -- successors 105 
    -- members (4) 
      -- 	branch_block_stmt_281/merge_stmt_317__entry__
      -- 	branch_block_stmt_281/if_stmt_311__exit__
      -- 	branch_block_stmt_281/if_stmt_311_dead_link/$exit
      -- 	branch_block_stmt_281/merge_stmt_317_dead_link/$entry
      -- 
    cp_elements(33) <= cp_elements(32);
    -- CP-element group 34 transition  output  bypass 
    -- predecessors 1 
    -- successors 35 
    -- members (3) 
      -- 	branch_block_stmt_281/if_stmt_311_eval_test/$entry
      -- 	branch_block_stmt_281/if_stmt_311_eval_test/$exit
      -- 	branch_block_stmt_281/if_stmt_311_eval_test/branch_req
      -- 
    cp_elements(34) <= cp_elements(1);
    branch_req_1702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => if_stmt_311_branch_req_0); -- 
    -- CP-element group 35 branch  place  bypass 
    -- predecessors 34 
    -- successors 36 38 
    -- members (1) 
      -- 	branch_block_stmt_281/simple_obj_ref_312_place
      -- 
    cp_elements(35) <= cp_elements(34);
    -- CP-element group 36 transition  bypass 
    -- predecessors 35 
    -- successors 37 
    -- members (1) 
      -- 	branch_block_stmt_281/if_stmt_311_if_link/$entry
      -- 
    cp_elements(36) <= cp_elements(35);
    -- CP-element group 37 transition  place  input  no-bypass 
    -- predecessors 36 
    -- successors 2 
    -- members (9) 
      -- 	branch_block_stmt_281/if_stmt_311_if_link/$exit
      -- 	branch_block_stmt_281/if_stmt_311_if_link/if_choice_transition
      -- 	branch_block_stmt_281/bb_1_bb_2
      -- 	branch_block_stmt_281/bb_1_bb_2_PhiReq/$entry
      -- 	branch_block_stmt_281/bb_1_bb_2_PhiReq/$exit
      -- 	branch_block_stmt_281/merge_stmt_317_PhiReqMerge
      -- 	branch_block_stmt_281/merge_stmt_317_PhiAck/$entry
      -- 	branch_block_stmt_281/merge_stmt_317_PhiAck/$exit
      -- 	branch_block_stmt_281/merge_stmt_317_PhiAck/dummy
      -- 
    if_choice_transition_1707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_311_branch_ack_1, ack => cp_elements(37)); -- 
    -- CP-element group 38 transition  bypass 
    -- predecessors 35 
    -- successors 39 
    -- members (1) 
      -- 	branch_block_stmt_281/if_stmt_311_else_link/$entry
      -- 
    cp_elements(38) <= cp_elements(35);
    -- CP-element group 39 transition  place  input  no-bypass 
    -- predecessors 38 
    -- successors 
    -- members (21) 
      -- 	branch_block_stmt_281/branch_block_stmt_281__exit__
      -- 	branch_block_stmt_281/$exit
      -- 	branch_block_stmt_281/merge_stmt_361__exit__
      -- 	branch_block_stmt_281/return__
      -- 	branch_block_stmt_281/merge_stmt_359__exit__
      -- 	$exit
      -- 	branch_block_stmt_281/if_stmt_311_else_link/$exit
      -- 	branch_block_stmt_281/if_stmt_311_else_link/else_choice_transition
      -- 	branch_block_stmt_281/bb_1_bb_4
      -- 	branch_block_stmt_281/bb_1_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_281/bb_1_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_281/merge_stmt_359_PhiReqMerge
      -- 	branch_block_stmt_281/merge_stmt_359_PhiAck/$entry
      -- 	branch_block_stmt_281/merge_stmt_359_PhiAck/$exit
      -- 	branch_block_stmt_281/merge_stmt_359_PhiAck/dummy
      -- 	branch_block_stmt_281/return___PhiReq/$entry
      -- 	branch_block_stmt_281/return___PhiReq/$exit
      -- 	branch_block_stmt_281/merge_stmt_361_PhiReqMerge
      -- 	branch_block_stmt_281/merge_stmt_361_PhiAck/$entry
      -- 	branch_block_stmt_281/merge_stmt_361_PhiAck/$exit
      -- 	branch_block_stmt_281/merge_stmt_361_PhiAck/dummy
      -- 
    else_choice_transition_1711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_311_branch_ack_0, ack => cp_elements(39)); -- 
    -- CP-element group 40 fork  transition  bypass 
    -- predecessors 2 
    -- successors 41 48 62 71 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/$entry
      -- 
    cp_elements(40) <= cp_elements(2);
    -- CP-element group 41 transition  output  bypass 
    -- predecessors 40 
    -- successors 42 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_319_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_319_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_319_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_addr_resize/base_resize_req
      -- 
    cp_elements(41) <= cp_elements(40);
    base_resize_req_1733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_320_base_resize_req_0); -- 
    -- CP-element group 42 transition  input  output  no-bypass 
    -- predecessors 41 
    -- successors 43 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_base_resize_ack_0, ack => cp_elements(42)); -- 
    sum_rename_req_1738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_320_root_address_inst_req_0); -- 
    -- CP-element group 43 transition  input  output  no-bypass 
    -- predecessors 42 
    -- successors 44 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_root_address_inst_ack_0, ack => cp_elements(43)); -- 
    root_register_req_1743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_320_addr_0_req_0); -- 
    -- CP-element group 44 transition  input  output  no-bypass 
    -- predecessors 43 
    -- successors 45 
    -- members (8) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_word_addrgen/root_register_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/word_access_0/rr
      -- 
    root_register_ack_1744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_addr_0_ack_0, ack => cp_elements(44)); -- 
    rr_1754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_320_load_0_req_0); -- 
    -- CP-element group 45 transition  input  output  no-bypass 
    -- predecessors 44 
    -- successors 46 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/word_access_0/cr
      -- 
    ra_1755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_load_0_ack_0, ack => cp_elements(45)); -- 
    cr_1765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_320_load_0_req_1); -- 
    -- CP-element group 46 transition  input  output  no-bypass 
    -- predecessors 45 
    -- successors 47 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/merge_req
      -- 
    ca_1766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_load_0_ack_1, ack => cp_elements(46)); -- 
    merge_req_1767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_320_gather_scatter_req_0); -- 
    -- CP-element group 47 transition  input  output  no-bypass 
    -- predecessors 46 
    -- successors 50 
    -- members (12) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_321_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_321_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_321_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_320_complete/merge_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_computed_0
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_323_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_323_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_323_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_resize_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_resize_0/index_resize_req
      -- 
    merge_ack_1768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_320_gather_scatter_ack_0, ack => cp_elements(47)); -- 
    index_resize_req_1786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => array_obj_ref_324_index_0_resize_req_0); -- 
    -- CP-element group 48 transition  bypass 
    -- predecessors 40 
    -- successors 49 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_trigger_
      -- 
    cp_elements(48) <= cp_elements(40);
    -- CP-element group 49 join  transition  output  no-bypass 
    -- predecessors 48 53 
    -- successors 54 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_complete/final_reg_req
      -- 
    cpelement_group_49 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(48);
      predecessors(1) <= cp_elements(53);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(49)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(49),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => addr_of_325_final_reg_req_0); -- 
    -- CP-element group 50 transition  input  output  no-bypass 
    -- predecessors 47 
    -- successors 51 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_resized_0
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_resize_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_scale_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_1787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_324_index_0_resize_ack_0, ack => cp_elements(50)); -- 
    scale_rename_req_1791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => array_obj_ref_324_index_0_rename_req_0); -- 
    -- CP-element group 51 transition  input  output  no-bypass 
    -- predecessors 50 
    -- successors 52 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_indices_scaled
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_scale_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_add_indices/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_add_indices/final_index_req
      -- 
    scale_rename_ack_1792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_324_index_0_rename_ack_0, ack => cp_elements(51)); -- 
    final_index_req_1796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_324_offset_inst_req_0); -- 
    -- CP-element group 52 transition  input  output  no-bypass 
    -- predecessors 51 
    -- successors 53 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_offset_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_add_indices/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_add_indices/final_index_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_1797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_324_offset_inst_ack_0, ack => cp_elements(52)); -- 
    sum_rename_req_1801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_324_root_address_inst_req_0); -- 
    -- CP-element group 53 transition  input  no-bypass 
    -- predecessors 52 
    -- successors 49 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/array_obj_ref_324_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_324_root_address_inst_ack_0, ack => cp_elements(53)); -- 
    -- CP-element group 54 transition  input  output  no-bypass 
    -- predecessors 49 
    -- successors 55 
    -- members (12) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_326_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_326_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_326_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/addr_of_325_complete/final_reg_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_328_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_328_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_328_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_325_final_reg_ack_0, ack => cp_elements(54)); -- 
    base_resize_req_1824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_329_base_resize_req_0); -- 
    -- CP-element group 55 transition  input  output  no-bypass 
    -- predecessors 54 
    -- successors 56 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_base_resize_ack_0, ack => cp_elements(55)); -- 
    sum_rename_req_1829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_329_root_address_inst_req_0); -- 
    -- CP-element group 56 transition  input  output  no-bypass 
    -- predecessors 55 
    -- successors 57 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_root_address_inst_ack_0, ack => cp_elements(56)); -- 
    root_register_req_1834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_329_addr_0_req_0); -- 
    -- CP-element group 57 transition  input  output  no-bypass 
    -- predecessors 56 
    -- successors 58 
    -- members (8) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_word_addrgen/root_register_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/word_access_0/rr
      -- 
    root_register_ack_1835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_addr_0_ack_0, ack => cp_elements(57)); -- 
    rr_1845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => ptr_deref_329_load_0_req_0); -- 
    -- CP-element group 58 transition  input  output  no-bypass 
    -- predecessors 57 
    -- successors 59 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/word_access_0/cr
      -- 
    ra_1846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_load_0_ack_0, ack => cp_elements(58)); -- 
    cr_1856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_329_load_0_req_1); -- 
    -- CP-element group 59 transition  input  output  no-bypass 
    -- predecessors 58 
    -- successors 60 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/merge_req
      -- 
    ca_1857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_load_0_ack_1, ack => cp_elements(59)); -- 
    merge_req_1858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_329_gather_scatter_req_0); -- 
    -- CP-element group 60 transition  input  no-bypass 
    -- predecessors 59 
    -- successors 61 
    -- members (11) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_330_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_330_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_330_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_329_complete/merge_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_334_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_334_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_333_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_333_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_333_completed_
      -- 
    merge_ack_1859_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_329_gather_scatter_ack_0, ack => cp_elements(60)); -- 
    -- CP-element group 61 join  transition  output  bypass 
    -- predecessors 60 65 
    -- successors 66 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/split_req
      -- 
    cpelement_group_61 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(60);
      predecessors(1) <= cp_elements(65);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(61)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(61),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_332_gather_scatter_req_0); -- 
    -- CP-element group 62 transition  output  bypass 
    -- predecessors 40 
    -- successors 63 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_331_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_331_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_331_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_addr_resize/base_resize_req
      -- 
    cp_elements(62) <= cp_elements(40);
    base_resize_req_1879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_332_base_resize_req_0); -- 
    -- CP-element group 63 transition  input  output  no-bypass 
    -- predecessors 62 
    -- successors 64 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1880_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_base_resize_ack_0, ack => cp_elements(63)); -- 
    sum_rename_req_1884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_332_root_address_inst_req_0); -- 
    -- CP-element group 64 transition  input  output  no-bypass 
    -- predecessors 63 
    -- successors 65 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_root_address_inst_ack_0, ack => cp_elements(64)); -- 
    root_register_req_1889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_332_addr_0_req_0); -- 
    -- CP-element group 65 transition  input  no-bypass 
    -- predecessors 64 
    -- successors 61 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_word_addrgen/root_register_ack
      -- 
    root_register_ack_1890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_addr_0_ack_0, ack => cp_elements(65)); -- 
    -- CP-element group 66 transition  input  output  no-bypass 
    -- predecessors 61 
    -- successors 67 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/split_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/word_access_0/rr
      -- 
    split_ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_gather_scatter_ack_0, ack => cp_elements(66)); -- 
    rr_1902_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => ptr_deref_332_store_0_req_0); -- 
    -- CP-element group 67 fork  transition  input  no-bypass 
    -- predecessors 66 
    -- successors 68 70 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_request/word_access/word_access_0/ra
      -- 
    ra_1903_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_store_0_ack_0, ack => cp_elements(67)); -- 
    -- CP-element group 68 transition  output  bypass 
    -- predecessors 67 
    -- successors 69 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/word_access_0/cr
      -- 
    cp_elements(68) <= cp_elements(67);
    cr_1913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_332_store_0_req_1); -- 
    -- CP-element group 69 transition  input  no-bypass 
    -- predecessors 68 
    -- successors 78 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_334_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_332_complete/word_access/word_access_0/ca
      -- 
    ca_1914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_332_store_0_ack_1, ack => cp_elements(69)); -- 
    -- CP-element group 70 join  transition  output  bypass 
    -- predecessors 67 74 
    -- successors 75 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/word_access_0/rr
      -- 
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(67);
      predecessors(1) <= cp_elements(74);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(70)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1952_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_337_load_0_req_0); -- 
    -- CP-element group 71 transition  output  bypass 
    -- predecessors 40 
    -- successors 72 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_336_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_336_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/simple_obj_ref_336_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_addr_resize/base_resize_req
      -- 
    cp_elements(71) <= cp_elements(40);
    base_resize_req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_337_base_resize_req_0); -- 
    -- CP-element group 72 transition  input  output  no-bypass 
    -- predecessors 71 
    -- successors 73 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_1932_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_base_resize_ack_0, ack => cp_elements(72)); -- 
    sum_rename_req_1936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_337_root_address_inst_req_0); -- 
    -- CP-element group 73 transition  input  output  no-bypass 
    -- predecessors 72 
    -- successors 74 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_word_addrgen/root_register_req
      -- 
    sum_rename_ack_1937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_root_address_inst_ack_0, ack => cp_elements(73)); -- 
    root_register_req_1941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => ptr_deref_337_addr_0_req_0); -- 
    -- CP-element group 74 transition  input  no-bypass 
    -- predecessors 73 
    -- successors 70 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_word_addrgen/root_register_ack
      -- 
    root_register_ack_1942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_addr_0_ack_0, ack => cp_elements(74)); -- 
    -- CP-element group 75 transition  input  output  no-bypass 
    -- predecessors 70 
    -- successors 76 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/word_access_0/cr
      -- 
    ra_1953_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_load_0_ack_0, ack => cp_elements(75)); -- 
    cr_1963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => ptr_deref_337_load_0_req_1); -- 
    -- CP-element group 76 transition  input  output  no-bypass 
    -- predecessors 75 
    -- successors 77 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/merge_req
      -- 
    ca_1964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_load_0_ack_1, ack => cp_elements(76)); -- 
    merge_req_1965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_337_gather_scatter_req_0); -- 
    -- CP-element group 77 transition  input  no-bypass 
    -- predecessors 76 
    -- successors 78 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_338_trigger_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_338_active_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/assign_stmt_338_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_completed_
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/ptr_deref_337_complete/merge_ack
      -- 
    merge_ack_1966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_337_gather_scatter_ack_0, ack => cp_elements(77)); -- 
    -- CP-element group 78 join  transition  bypass 
    -- predecessors 69 77 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_321_to_assign_stmt_338/$exit
      -- 
    cpelement_group_78 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(69);
      predecessors(1) <= cp_elements(77);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(78)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(78),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 79 transition  place  input  no-bypass 
    -- predecessors 3 
    -- successors 80 
    -- members (16) 
      -- 	branch_block_stmt_281/bb_2_bb_3
      -- 	branch_block_stmt_281/merge_stmt_343__exit__
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357__entry__
      -- 	branch_block_stmt_281/assign_stmt_341__exit__
      -- 	branch_block_stmt_281/assign_stmt_341/$exit
      -- 	branch_block_stmt_281/assign_stmt_341/assign_stmt_341_completed_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_active_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_completed_
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_341/simple_obj_ref_339_complete/pipe_wack
      -- 	branch_block_stmt_281/bb_2_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_281/bb_2_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_281/merge_stmt_343_PhiReqMerge
      -- 	branch_block_stmt_281/merge_stmt_343_PhiAck/$entry
      -- 	branch_block_stmt_281/merge_stmt_343_PhiAck/$exit
      -- 	branch_block_stmt_281/merge_stmt_343_PhiAck/dummy
      -- 
    pipe_wack_1983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_339_inst_ack_0, ack => cp_elements(79)); -- 
    -- CP-element group 80 fork  transition  bypass 
    -- predecessors 79 
    -- successors 81 88 95 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/$entry
      -- 
    cp_elements(80) <= cp_elements(79);
    -- CP-element group 81 transition  output  bypass 
    -- predecessors 80 
    -- successors 82 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_345_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_345_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_345_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_addr_resize/base_resize_req
      -- 
    cp_elements(81) <= cp_elements(80);
    base_resize_req_2003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_346_base_resize_req_0); -- 
    -- CP-element group 82 transition  input  output  no-bypass 
    -- predecessors 81 
    -- successors 83 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_base_resize_ack_0, ack => cp_elements(82)); -- 
    sum_rename_req_2008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_346_root_address_inst_req_0); -- 
    -- CP-element group 83 transition  input  output  no-bypass 
    -- predecessors 82 
    -- successors 84 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_root_address_inst_ack_0, ack => cp_elements(83)); -- 
    root_register_req_2013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_346_addr_0_req_0); -- 
    -- CP-element group 84 transition  input  output  no-bypass 
    -- predecessors 83 
    -- successors 85 
    -- members (8) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_word_addrgen/root_register_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/word_access_0/rr
      -- 
    root_register_ack_2014_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_addr_0_ack_0, ack => cp_elements(84)); -- 
    rr_2024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_346_load_0_req_0); -- 
    -- CP-element group 85 transition  input  output  no-bypass 
    -- predecessors 84 
    -- successors 86 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/word_access_0/cr
      -- 
    ra_2025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_load_0_ack_0, ack => cp_elements(85)); -- 
    cr_2035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_346_load_0_req_1); -- 
    -- CP-element group 86 transition  input  output  no-bypass 
    -- predecessors 85 
    -- successors 87 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/merge_req
      -- 
    ca_2036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_load_0_ack_1, ack => cp_elements(86)); -- 
    merge_req_2037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_346_gather_scatter_req_0); -- 
    -- CP-element group 87 fork  transition  input  no-bypass 
    -- predecessors 86 
    -- successors 90 91 
    -- members (10) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_347_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_347_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_347_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_346_complete/merge_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_349_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_349_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_349_completed_
      -- 
    merge_ack_2038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_346_gather_scatter_ack_0, ack => cp_elements(87)); -- 
    -- CP-element group 88 transition  bypass 
    -- predecessors 80 
    -- successors 102 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_active_
      -- 
    cp_elements(88) <= cp_elements(80);
    -- CP-element group 89 join  transition  bypass 
    -- predecessors 92 93 
    -- successors 94 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_353_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_353_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_353_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_357_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_357_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_356_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_356_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_356_completed_
      -- 
    cpelement_group_89 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(92);
      predecessors(1) <= cp_elements(93);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(89)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(89),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 90 transition  output  bypass 
    -- predecessors 87 
    -- successors 92 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_sample_start_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Sample/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Sample/rr
      -- 
    cp_elements(90) <= cp_elements(87);
    rr_2055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => binary_352_inst_req_0); -- 
    -- CP-element group 91 transition  output  bypass 
    -- predecessors 87 
    -- successors 93 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_update_start_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Update/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Update/cr
      -- 
    cp_elements(91) <= cp_elements(87);
    cr_2060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => binary_352_inst_req_1); -- 
    -- CP-element group 92 transition  input  no-bypass 
    -- predecessors 90 
    -- successors 89 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_sample_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Sample/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Sample/ra
      -- 
    ra_2056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_352_inst_ack_0, ack => cp_elements(92)); -- 
    -- CP-element group 93 transition  input  no-bypass 
    -- predecessors 91 
    -- successors 89 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_update_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Update/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/binary_352_Update/ca
      -- 
    ca_2061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_352_inst_ack_1, ack => cp_elements(93)); -- 
    -- CP-element group 94 join  transition  output  bypass 
    -- predecessors 89 98 
    -- successors 99 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/split_req
      -- 
    cpelement_group_94 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(89);
      predecessors(1) <= cp_elements(98);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(94)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(94),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_355_gather_scatter_req_0); -- 
    -- CP-element group 95 transition  output  bypass 
    -- predecessors 80 
    -- successors 96 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_354_trigger_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_354_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/simple_obj_ref_354_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_addr_resize/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_addr_resize/base_resize_req
      -- 
    cp_elements(95) <= cp_elements(80);
    base_resize_req_2081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_355_base_resize_req_0); -- 
    -- CP-element group 96 transition  input  output  no-bypass 
    -- predecessors 95 
    -- successors 97 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_address_resized
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_addr_resize/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_plus_offset/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_base_resize_ack_0, ack => cp_elements(96)); -- 
    sum_rename_req_2086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_355_root_address_inst_req_0); -- 
    -- CP-element group 97 transition  input  output  no-bypass 
    -- predecessors 96 
    -- successors 98 
    -- members (5) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_root_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_plus_offset/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_word_addrgen/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_root_address_inst_ack_0, ack => cp_elements(97)); -- 
    root_register_req_2091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_355_addr_0_req_0); -- 
    -- CP-element group 98 transition  input  no-bypass 
    -- predecessors 97 
    -- successors 94 
    -- members (3) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_word_address_calculated
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_word_addrgen/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_word_addrgen/root_register_ack
      -- 
    root_register_ack_2092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_addr_0_ack_0, ack => cp_elements(98)); -- 
    -- CP-element group 99 transition  input  output  no-bypass 
    -- predecessors 94 
    -- successors 100 
    -- members (4) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/split_ack
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/word_access_0/rr
      -- 
    split_ack_2097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_gather_scatter_ack_0, ack => cp_elements(99)); -- 
    rr_2104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => ptr_deref_355_store_0_req_0); -- 
    -- CP-element group 100 transition  input  output  no-bypass 
    -- predecessors 99 
    -- successors 101 
    -- members (9) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_active_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/word_access_0/cr
      -- 
    ra_2105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_store_0_ack_0, ack => cp_elements(100)); -- 
    cr_2115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_355_store_0_req_1); -- 
    -- CP-element group 101 transition  input  no-bypass 
    -- predecessors 100 
    -- successors 102 
    -- members (6) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/assign_stmt_357_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_completed_
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/ptr_deref_355_complete/word_access/word_access_0/ca
      -- 
    ca_2116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_355_store_0_ack_1, ack => cp_elements(101)); -- 
    -- CP-element group 102 join  transition  bypass 
    -- predecessors 88 101 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_281/assign_stmt_347_to_assign_stmt_357/$exit
      -- 
    cpelement_group_102 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(88);
      predecessors(1) <= cp_elements(101);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(102)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(102),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 103 merge  place  bypass 
    -- predecessors 4 14 
    -- successors 104 
    -- members (1) 
      -- 	branch_block_stmt_281/merge_stmt_298_PhiReqMerge
      -- 
    cp_elements(103) <= OrReduce(cp_elements(4) & cp_elements(14));
    -- CP-element group 104 transition  place  bypass 
    -- predecessors 103 
    -- successors 15 
    -- members (5) 
      -- 	branch_block_stmt_281/merge_stmt_298__exit__
      -- 	branch_block_stmt_281/assign_stmt_302_to_assign_stmt_310__entry__
      -- 	branch_block_stmt_281/merge_stmt_298_PhiAck/$entry
      -- 	branch_block_stmt_281/merge_stmt_298_PhiAck/$exit
      -- 	branch_block_stmt_281/merge_stmt_298_PhiAck/dummy
      -- 
    cp_elements(104) <= cp_elements(103);
    -- CP-element group 105 transition  dead  bypass 
    -- predecessors 33 
    -- successors 106 
    -- members (1) 
      -- 	branch_block_stmt_281/merge_stmt_317_dead_link/dead_transition
      -- 
    cp_elements(105) <= false;
    -- CP-element group 106 transition  bypass 
    -- predecessors 105 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_281/merge_stmt_317_dead_link/$exit
      -- 
    cp_elements(106) <= cp_elements(105);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_324_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_324_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_324_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_324_root_address : std_logic_vector(6 downto 0);
    signal iNsTr_14_347 : std_logic_vector(31 downto 0);
    signal iNsTr_15_353 : std_logic_vector(31 downto 0);
    signal iNsTr_2_302 : std_logic_vector(31 downto 0);
    signal iNsTr_3_310 : std_logic_vector(0 downto 0);
    signal iNsTr_5_321 : std_logic_vector(31 downto 0);
    signal iNsTr_6_326 : std_logic_vector(31 downto 0);
    signal iNsTr_7_330 : std_logic_vector(31 downto 0);
    signal iNsTr_9_338 : std_logic_vector(31 downto 0);
    signal idx_287 : std_logic_vector(31 downto 0);
    signal ptr_deref_293_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_293_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_293_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_293_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_293_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_293_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_301_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_301_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_301_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_301_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_301_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_320_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_320_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_320_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_320_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_320_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_329_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_329_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_329_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_329_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_329_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_332_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_332_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_332_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_332_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_332_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_332_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_337_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_337_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_337_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_337_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_337_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_346_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_346_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_346_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_346_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_346_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_355_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_355_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_355_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_355_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_355_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_355_word_offset_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_323_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_323_scaled : std_logic_vector(6 downto 0);
    signal type_cast_295_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_305_wire : std_logic_vector(31 downto 0);
    signal type_cast_308_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_351_wire_constant : std_logic_vector(31 downto 0);
    signal val_291 : std_logic_vector(31 downto 0);
    signal xxsendResultxxbodyxxidx_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxsendResultxxbodyxxval_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_324_offset_scale_factor_0 <= "0000001";
    array_obj_ref_324_resized_base_address <= "0000000";
    idx_287 <= "00000000000000000000000000000000";
    ptr_deref_293_word_offset_0 <= "0";
    ptr_deref_301_word_offset_0 <= "0";
    ptr_deref_320_word_offset_0 <= "0";
    ptr_deref_329_word_offset_0 <= "0000000";
    ptr_deref_332_word_offset_0 <= "0";
    ptr_deref_337_word_offset_0 <= "0";
    ptr_deref_346_word_offset_0 <= "0";
    ptr_deref_355_word_offset_0 <= "0";
    type_cast_295_wire_constant <= "00000000000000000000000000000000";
    type_cast_308_wire_constant <= "00000000000000000000000001000000";
    type_cast_351_wire_constant <= "00000000000000000000000000000001";
    val_291 <= "00000000000000000000000000000000";
    xxsendResultxxbodyxxidx_alloc_base_address <= "0";
    xxsendResultxxbodyxxval_alloc_base_address <= "0";
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_325_final_reg_req_0,addr_of_325_final_reg_ack_0,sl_one,"addr_of_325_final_reg ",false,array_obj_ref_324_root_address,
    false,iNsTr_6_326);
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_325_final_reg_req_0;
      addr_of_325_final_reg_ack_0 <= ack; 
      addr_of_325_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_324_root_address, dout => iNsTr_6_326, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_305_inst_req_0,type_cast_305_inst_ack_0,sl_one,"type_cast_305_inst ",false,iNsTr_2_302,
    false,type_cast_305_wire);
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_305_inst_req_0;
      type_cast_305_inst_ack_0 <= ack; 
      type_cast_305_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_2_302, dout => type_cast_305_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_324_index_0_rename_req_0,array_obj_ref_324_index_0_rename_ack_0,sl_one,"array_obj_ref_324_index_0_rename ",false,simple_obj_ref_323_resized,
    false,simple_obj_ref_323_scaled);
    array_obj_ref_324_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_324_index_0_rename_ack_0 <= array_obj_ref_324_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_323_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_323_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_324_index_0_resize_req_0,array_obj_ref_324_index_0_resize_ack_0,sl_one,"array_obj_ref_324_index_0_resize ",false,iNsTr_5_321,
    false,simple_obj_ref_323_resized);
    array_obj_ref_324_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_324_index_0_resize_ack_0 <= array_obj_ref_324_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_5_321;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_323_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_324_offset_inst_req_0,array_obj_ref_324_offset_inst_ack_0,sl_one,"array_obj_ref_324_offset_inst ",false,simple_obj_ref_323_scaled,
    false,array_obj_ref_324_final_offset);
    array_obj_ref_324_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_324_offset_inst_ack_0 <= array_obj_ref_324_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_323_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_324_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_324_root_address_inst_req_0,array_obj_ref_324_root_address_inst_ack_0,sl_one,"array_obj_ref_324_root_address_inst ",false,array_obj_ref_324_final_offset,
    false,array_obj_ref_324_root_address);
    array_obj_ref_324_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_324_root_address_inst_ack_0 <= array_obj_ref_324_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_324_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_324_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_293_addr_0_req_0,ptr_deref_293_addr_0_ack_0,sl_one,"ptr_deref_293_addr_0 ",false,ptr_deref_293_root_address,
    false,ptr_deref_293_word_address_0);
    ptr_deref_293_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_293_addr_0_ack_0 <= ptr_deref_293_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_293_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_293_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_293_base_resize_req_0,ptr_deref_293_base_resize_ack_0,sl_one,"ptr_deref_293_base_resize ",false,idx_287,
    false,ptr_deref_293_resized_base_address);
    ptr_deref_293_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_293_base_resize_ack_0 <= ptr_deref_293_base_resize_req_0;
      in_aggregated_sig <= idx_287;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_293_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_293_gather_scatter_req_0,ptr_deref_293_gather_scatter_ack_0,sl_one,"ptr_deref_293_gather_scatter ",false,type_cast_295_wire_constant,
    false,ptr_deref_293_data_0);
    ptr_deref_293_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_293_gather_scatter_ack_0 <= ptr_deref_293_gather_scatter_req_0;
      in_aggregated_sig <= type_cast_295_wire_constant;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_293_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_293_root_address_inst_req_0,ptr_deref_293_root_address_inst_ack_0,sl_one,"ptr_deref_293_root_address_inst ",false,ptr_deref_293_resized_base_address,
    false,ptr_deref_293_root_address);
    ptr_deref_293_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_293_root_address_inst_ack_0 <= ptr_deref_293_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_293_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_293_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_301_addr_0_req_0,ptr_deref_301_addr_0_ack_0,sl_one,"ptr_deref_301_addr_0 ",false,ptr_deref_301_root_address,
    false,ptr_deref_301_word_address_0);
    ptr_deref_301_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_301_addr_0_ack_0 <= ptr_deref_301_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_301_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_301_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_301_base_resize_req_0,ptr_deref_301_base_resize_ack_0,sl_one,"ptr_deref_301_base_resize ",false,idx_287,
    false,ptr_deref_301_resized_base_address);
    ptr_deref_301_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_301_base_resize_ack_0 <= ptr_deref_301_base_resize_req_0;
      in_aggregated_sig <= idx_287;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_301_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_301_gather_scatter_req_0,ptr_deref_301_gather_scatter_ack_0,sl_one,"ptr_deref_301_gather_scatter ",false,ptr_deref_301_data_0,
    false,iNsTr_2_302);
    ptr_deref_301_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_301_gather_scatter_ack_0 <= ptr_deref_301_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_301_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_2_302 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_301_root_address_inst_req_0,ptr_deref_301_root_address_inst_ack_0,sl_one,"ptr_deref_301_root_address_inst ",false,ptr_deref_301_resized_base_address,
    false,ptr_deref_301_root_address);
    ptr_deref_301_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_301_root_address_inst_ack_0 <= ptr_deref_301_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_301_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_301_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_320_addr_0_req_0,ptr_deref_320_addr_0_ack_0,sl_one,"ptr_deref_320_addr_0 ",false,ptr_deref_320_root_address,
    false,ptr_deref_320_word_address_0);
    ptr_deref_320_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_320_addr_0_ack_0 <= ptr_deref_320_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_320_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_320_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_320_base_resize_req_0,ptr_deref_320_base_resize_ack_0,sl_one,"ptr_deref_320_base_resize ",false,idx_287,
    false,ptr_deref_320_resized_base_address);
    ptr_deref_320_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_320_base_resize_ack_0 <= ptr_deref_320_base_resize_req_0;
      in_aggregated_sig <= idx_287;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_320_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_320_gather_scatter_req_0,ptr_deref_320_gather_scatter_ack_0,sl_one,"ptr_deref_320_gather_scatter ",false,ptr_deref_320_data_0,
    false,iNsTr_5_321);
    ptr_deref_320_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_320_gather_scatter_ack_0 <= ptr_deref_320_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_320_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_5_321 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_320_root_address_inst_req_0,ptr_deref_320_root_address_inst_ack_0,sl_one,"ptr_deref_320_root_address_inst ",false,ptr_deref_320_resized_base_address,
    false,ptr_deref_320_root_address);
    ptr_deref_320_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_320_root_address_inst_ack_0 <= ptr_deref_320_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_320_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_320_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_329_addr_0_req_0,ptr_deref_329_addr_0_ack_0,sl_one,"ptr_deref_329_addr_0 ",false,ptr_deref_329_root_address,
    false,ptr_deref_329_word_address_0);
    ptr_deref_329_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_329_addr_0_ack_0 <= ptr_deref_329_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_329_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_329_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_329_base_resize_req_0,ptr_deref_329_base_resize_ack_0,sl_one,"ptr_deref_329_base_resize ",false,iNsTr_6_326,
    false,ptr_deref_329_resized_base_address);
    ptr_deref_329_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_329_base_resize_ack_0 <= ptr_deref_329_base_resize_req_0;
      in_aggregated_sig <= iNsTr_6_326;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_329_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_329_gather_scatter_req_0,ptr_deref_329_gather_scatter_ack_0,sl_one,"ptr_deref_329_gather_scatter ",false,ptr_deref_329_data_0,
    false,iNsTr_7_330);
    ptr_deref_329_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_329_gather_scatter_ack_0 <= ptr_deref_329_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_329_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_7_330 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_329_root_address_inst_req_0,ptr_deref_329_root_address_inst_ack_0,sl_one,"ptr_deref_329_root_address_inst ",false,ptr_deref_329_resized_base_address,
    false,ptr_deref_329_root_address);
    ptr_deref_329_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_329_root_address_inst_ack_0 <= ptr_deref_329_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_329_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_329_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_332_addr_0_req_0,ptr_deref_332_addr_0_ack_0,sl_one,"ptr_deref_332_addr_0 ",false,ptr_deref_332_root_address,
    false,ptr_deref_332_word_address_0);
    ptr_deref_332_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_332_addr_0_ack_0 <= ptr_deref_332_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_332_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_332_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_332_base_resize_req_0,ptr_deref_332_base_resize_ack_0,sl_one,"ptr_deref_332_base_resize ",false,val_291,
    false,ptr_deref_332_resized_base_address);
    ptr_deref_332_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_332_base_resize_ack_0 <= ptr_deref_332_base_resize_req_0;
      in_aggregated_sig <= val_291;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_332_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_332_gather_scatter_req_0,ptr_deref_332_gather_scatter_ack_0,sl_one,"ptr_deref_332_gather_scatter ",false,iNsTr_7_330,
    false,ptr_deref_332_data_0);
    ptr_deref_332_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_332_gather_scatter_ack_0 <= ptr_deref_332_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_7_330;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_332_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_332_root_address_inst_req_0,ptr_deref_332_root_address_inst_ack_0,sl_one,"ptr_deref_332_root_address_inst ",false,ptr_deref_332_resized_base_address,
    false,ptr_deref_332_root_address);
    ptr_deref_332_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_332_root_address_inst_ack_0 <= ptr_deref_332_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_332_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_332_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_337_addr_0_req_0,ptr_deref_337_addr_0_ack_0,sl_one,"ptr_deref_337_addr_0 ",false,ptr_deref_337_root_address,
    false,ptr_deref_337_word_address_0);
    ptr_deref_337_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_337_addr_0_ack_0 <= ptr_deref_337_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_337_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_337_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_337_base_resize_req_0,ptr_deref_337_base_resize_ack_0,sl_one,"ptr_deref_337_base_resize ",false,val_291,
    false,ptr_deref_337_resized_base_address);
    ptr_deref_337_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_337_base_resize_ack_0 <= ptr_deref_337_base_resize_req_0;
      in_aggregated_sig <= val_291;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_337_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_337_gather_scatter_req_0,ptr_deref_337_gather_scatter_ack_0,sl_one,"ptr_deref_337_gather_scatter ",false,ptr_deref_337_data_0,
    false,iNsTr_9_338);
    ptr_deref_337_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_337_gather_scatter_ack_0 <= ptr_deref_337_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_337_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_9_338 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_337_root_address_inst_req_0,ptr_deref_337_root_address_inst_ack_0,sl_one,"ptr_deref_337_root_address_inst ",false,ptr_deref_337_resized_base_address,
    false,ptr_deref_337_root_address);
    ptr_deref_337_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_337_root_address_inst_ack_0 <= ptr_deref_337_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_337_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_337_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_346_addr_0_req_0,ptr_deref_346_addr_0_ack_0,sl_one,"ptr_deref_346_addr_0 ",false,ptr_deref_346_root_address,
    false,ptr_deref_346_word_address_0);
    ptr_deref_346_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_346_addr_0_ack_0 <= ptr_deref_346_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_346_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_346_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_346_base_resize_req_0,ptr_deref_346_base_resize_ack_0,sl_one,"ptr_deref_346_base_resize ",false,idx_287,
    false,ptr_deref_346_resized_base_address);
    ptr_deref_346_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_346_base_resize_ack_0 <= ptr_deref_346_base_resize_req_0;
      in_aggregated_sig <= idx_287;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_346_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_346_gather_scatter_req_0,ptr_deref_346_gather_scatter_ack_0,sl_one,"ptr_deref_346_gather_scatter ",false,ptr_deref_346_data_0,
    false,iNsTr_14_347);
    ptr_deref_346_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_346_gather_scatter_ack_0 <= ptr_deref_346_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_346_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_14_347 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_346_root_address_inst_req_0,ptr_deref_346_root_address_inst_ack_0,sl_one,"ptr_deref_346_root_address_inst ",false,ptr_deref_346_resized_base_address,
    false,ptr_deref_346_root_address);
    ptr_deref_346_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_346_root_address_inst_ack_0 <= ptr_deref_346_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_346_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_346_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_355_addr_0_req_0,ptr_deref_355_addr_0_ack_0,sl_one,"ptr_deref_355_addr_0 ",false,ptr_deref_355_root_address,
    false,ptr_deref_355_word_address_0);
    ptr_deref_355_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_355_addr_0_ack_0 <= ptr_deref_355_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_355_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_355_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_355_base_resize_req_0,ptr_deref_355_base_resize_ack_0,sl_one,"ptr_deref_355_base_resize ",false,idx_287,
    false,ptr_deref_355_resized_base_address);
    ptr_deref_355_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_355_base_resize_ack_0 <= ptr_deref_355_base_resize_req_0;
      in_aggregated_sig <= idx_287;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_355_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_355_gather_scatter_req_0,ptr_deref_355_gather_scatter_ack_0,sl_one,"ptr_deref_355_gather_scatter ",false,iNsTr_15_353,
    false,ptr_deref_355_data_0);
    ptr_deref_355_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_355_gather_scatter_ack_0 <= ptr_deref_355_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_15_353;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_355_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_355_root_address_inst_req_0,ptr_deref_355_root_address_inst_ack_0,sl_one,"ptr_deref_355_root_address_inst ",false,ptr_deref_355_resized_base_address,
    false,ptr_deref_355_root_address);
    ptr_deref_355_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_355_root_address_inst_ack_0 <= ptr_deref_355_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_355_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_355_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_311_branch_req_0," req0 if_stmt_311_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_311_branch_ack_0," ack0 if_stmt_311_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_311_branch_ack_1," ack1 if_stmt_311_branch");
    if_stmt_311_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_310;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_311_branch_req_0,
          ack0 => if_stmt_311_branch_ack_0,
          ack1 => if_stmt_311_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_309_inst_req_0,binary_309_inst_ack_0,binary_309_inst_req_1,binary_309_inst_ack_1,sl_one,"binary_309_inst",false,type_cast_305_wire & type_cast_308_wire_constant,
    false,iNsTr_3_310);
    -- shared split operator group (0) : binary_309_inst 
    ApIntSlt_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_305_wire;
      iNsTr_3_310 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_309_inst_req_0;
      reqR(0) <= binary_309_inst_req_1;
      binary_309_inst_ack_0 <= ackL(0); 
      binary_309_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_352_inst_req_0,binary_352_inst_ack_0,binary_352_inst_req_1,binary_352_inst_ack_1,sl_one,"binary_352_inst",false,iNsTr_14_347 & type_cast_351_wire_constant,
    false,iNsTr_15_353);
    -- shared split operator group (1) : binary_352_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_14_347;
      iNsTr_15_353 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_352_inst_req_0;
      reqR(0) <= binary_352_inst_req_1;
      binary_352_inst_ack_0 <= ackL(0); 
      binary_352_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_301_load_0_req_0,ptr_deref_301_load_0_ack_0,ptr_deref_301_load_0_req_1,ptr_deref_301_load_0_ack_1,sl_one,"ptr_deref_301_load_0",false,ptr_deref_301_word_address_0,
    false,ptr_deref_301_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_320_load_0_req_0,ptr_deref_320_load_0_ack_0,ptr_deref_320_load_0_req_1,ptr_deref_320_load_0_ack_1,sl_one,"ptr_deref_320_load_0",false,ptr_deref_320_word_address_0,
    false,ptr_deref_320_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_346_load_0_req_0,ptr_deref_346_load_0_ack_0,ptr_deref_346_load_0_req_1,ptr_deref_346_load_0_ack_1,sl_one,"ptr_deref_346_load_0",false,ptr_deref_346_word_address_0,
    false,ptr_deref_346_data_0);
    -- shared load operator group (0) : ptr_deref_301_load_0 ptr_deref_320_load_0 ptr_deref_346_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_301_load_0_req_0,
        ptr_deref_301_load_0_ack_0,
        ptr_deref_301_load_0_req_1,
        ptr_deref_301_load_0_ack_1,
        "ptr_deref_301_load_0",
        "memory_space_5" ,
        ptr_deref_301_data_0,
        ptr_deref_301_word_address_0,
        "ptr_deref_301_data_0",
        "ptr_deref_301_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_320_load_0_req_0,
        ptr_deref_320_load_0_ack_0,
        ptr_deref_320_load_0_req_1,
        ptr_deref_320_load_0_ack_1,
        "ptr_deref_320_load_0",
        "memory_space_5" ,
        ptr_deref_320_data_0,
        ptr_deref_320_word_address_0,
        "ptr_deref_320_data_0",
        "ptr_deref_320_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_346_load_0_req_0,
        ptr_deref_346_load_0_ack_0,
        ptr_deref_346_load_0_req_1,
        ptr_deref_346_load_0_ack_1,
        "ptr_deref_346_load_0",
        "memory_space_5" ,
        ptr_deref_346_data_0,
        ptr_deref_346_word_address_0,
        "ptr_deref_346_data_0",
        "ptr_deref_346_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_301_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_320_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_346_load_0_req_0;
      ptr_deref_301_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_320_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_346_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_301_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_320_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_346_load_0_req_1;
      ptr_deref_301_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_320_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_346_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_301_word_address_0 & ptr_deref_320_word_address_0 & ptr_deref_346_word_address_0;
      ptr_deref_301_data_0 <= data_out(95 downto 64);
      ptr_deref_320_data_0 <= data_out(63 downto 32);
      ptr_deref_346_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(0 downto 0),
          mtag => memory_space_5_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(31 downto 0),
          mtag => memory_space_5_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_329_load_0_req_0,ptr_deref_329_load_0_ack_0,ptr_deref_329_load_0_req_1,ptr_deref_329_load_0_ack_1,sl_one,"ptr_deref_329_load_0",false,ptr_deref_329_word_address_0,
    false,ptr_deref_329_data_0);
    -- shared load operator group (1) : ptr_deref_329_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_329_load_0_req_0,
        ptr_deref_329_load_0_ack_0,
        ptr_deref_329_load_0_req_1,
        ptr_deref_329_load_0_ack_1,
        "ptr_deref_329_load_0",
        "memory_space_2" ,
        ptr_deref_329_data_0,
        ptr_deref_329_word_address_0,
        "ptr_deref_329_data_0",
        "ptr_deref_329_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_329_load_0_req_0;
      ptr_deref_329_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_329_load_0_req_1;
      ptr_deref_329_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_329_word_address_0;
      ptr_deref_329_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_337_load_0_req_0,ptr_deref_337_load_0_ack_0,ptr_deref_337_load_0_req_1,ptr_deref_337_load_0_ack_1,sl_one,"ptr_deref_337_load_0",false,ptr_deref_337_word_address_0,
    false,ptr_deref_337_data_0);
    -- shared load operator group (2) : ptr_deref_337_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_337_load_0_req_0,
        ptr_deref_337_load_0_ack_0,
        ptr_deref_337_load_0_req_1,
        ptr_deref_337_load_0_ack_1,
        "ptr_deref_337_load_0",
        "memory_space_6" ,
        ptr_deref_337_data_0,
        ptr_deref_337_word_address_0,
        "ptr_deref_337_data_0",
        "ptr_deref_337_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_337_load_0_req_0;
      ptr_deref_337_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_337_load_0_req_1;
      ptr_deref_337_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_337_word_address_0;
      ptr_deref_337_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_355_store_0_req_0,ptr_deref_355_store_0_ack_0,ptr_deref_355_store_0_req_1,ptr_deref_355_store_0_ack_1,sl_one,"ptr_deref_355_store_0",false,ptr_deref_355_word_address_0 & ptr_deref_355_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_293_store_0_req_0,ptr_deref_293_store_0_ack_0,ptr_deref_293_store_0_req_1,ptr_deref_293_store_0_ack_1,sl_one,"ptr_deref_293_store_0",false,ptr_deref_293_word_address_0 & ptr_deref_293_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_355_store_0_req_0,
      ptr_deref_355_store_0_ack_0,
      ptr_deref_355_store_0_req_1,
      ptr_deref_355_store_0_ack_1,
      "ptr_deref_355_store_0",
      "memory_space_5" ,
      ptr_deref_355_data_0,
      ptr_deref_355_word_address_0,
      "ptr_deref_355_data_0",
      "ptr_deref_355_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_293_store_0_req_0,
      ptr_deref_293_store_0_ack_0,
      ptr_deref_293_store_0_req_1,
      ptr_deref_293_store_0_ack_1,
      "ptr_deref_293_store_0",
      "memory_space_5" ,
      ptr_deref_293_data_0,
      ptr_deref_293_word_address_0,
      "ptr_deref_293_data_0",
      "ptr_deref_293_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_355_store_0 ptr_deref_293_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_355_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_293_store_0_req_0;
      ptr_deref_355_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_293_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_355_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_293_store_0_req_1;
      ptr_deref_355_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_293_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_355_word_address_0 & ptr_deref_293_word_address_0;
      data_in <= ptr_deref_355_data_0 & ptr_deref_293_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(0 downto 0),
          mdata => memory_space_5_sr_data(31 downto 0),
          mtag => memory_space_5_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_332_store_0_req_0,ptr_deref_332_store_0_ack_0,ptr_deref_332_store_0_req_1,ptr_deref_332_store_0_ack_1,sl_one,"ptr_deref_332_store_0",false,ptr_deref_332_word_address_0 & ptr_deref_332_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_332_store_0_req_0,
      ptr_deref_332_store_0_ack_0,
      ptr_deref_332_store_0_req_1,
      ptr_deref_332_store_0_ack_1,
      "ptr_deref_332_store_0",
      "memory_space_6" ,
      ptr_deref_332_data_0,
      ptr_deref_332_word_address_0,
      "ptr_deref_332_data_0",
      "ptr_deref_332_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_332_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_332_store_0_req_0;
      ptr_deref_332_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_332_store_0_req_1;
      ptr_deref_332_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_332_word_address_0;
      data_in <= ptr_deref_332_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_339_inst_req_0,simple_obj_ref_339_inst_ack_0,sl_one,"simple_obj_ref_339_inst  PipeWrite to out_data_pipe",false,iNsTr_9_338,
    true, slv_zero);
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_339_inst_ack_0 then -- 
          assert false report " WritePipe out_data_pipe from wire iNsTr_9_338 value="  &  convert_slv_to_hex_string(iNsTr_9_338) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_339_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      req_unguarded(0) <= simple_obj_ref_339_inst_req_0;
      simple_obj_ref_339_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      data_in <= iNsTr_9_338;
      out_data_pipe_write_0: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_pipe_write_req(0),
          oack => out_data_pipe_pipe_write_ack(0),
          odata => out_data_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity vectorSum is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    x_vectorSum_x_call_reqs : out  std_logic_vector(0 downto 0);
    x_vectorSum_x_call_acks : in   std_logic_vector(0 downto 0);
    x_vectorSum_x_call_tag  :  out  std_logic_vector(0 downto 0);
    x_vectorSum_x_return_reqs : out  std_logic_vector(0 downto 0);
    x_vectorSum_x_return_acks : in   std_logic_vector(0 downto 0);
    x_vectorSum_x_return_tag :  in   std_logic_vector(0 downto 0);
    getData_call_reqs : out  std_logic_vector(0 downto 0);
    getData_call_acks : in   std_logic_vector(0 downto 0);
    getData_call_tag  :  out  std_logic_vector(0 downto 0);
    getData_return_reqs : out  std_logic_vector(0 downto 0);
    getData_return_acks : in   std_logic_vector(0 downto 0);
    getData_return_tag :  in   std_logic_vector(0 downto 0);
    sendResult_call_reqs : out  std_logic_vector(0 downto 0);
    sendResult_call_acks : in   std_logic_vector(0 downto 0);
    sendResult_call_tag  :  out  std_logic_vector(0 downto 0);
    sendResult_return_reqs : out  std_logic_vector(0 downto 0);
    sendResult_return_acks : in   std_logic_vector(0 downto 0);
    sendResult_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity vectorSum;
architecture Default of vectorSum is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal vectorSum_CP_8539_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_368_call_req_0 : boolean;
  signal call_stmt_368_call_ack_0 : boolean;
  signal call_stmt_368_call_req_1 : boolean;
  signal call_stmt_368_call_ack_1 : boolean;
  signal call_stmt_369_call_req_0 : boolean;
  signal call_stmt_369_call_ack_0 : boolean;
  signal call_stmt_369_call_req_1 : boolean;
  signal call_stmt_369_call_ack_1 : boolean;
  signal call_stmt_370_call_req_0 : boolean;
  signal call_stmt_370_call_ack_0 : boolean;
  signal call_stmt_370_call_req_1 : boolean;
  signal call_stmt_370_call_ack_1 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"vectorSum start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"vectorSum start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"vectorSum fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"vectorSum fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  vectorSum_CP_8539: Block -- control-path 
    signal cp_elements: BooleanArray(9 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 8 
    -- members (6) 
      -- 	$entry
      -- 	branch_block_stmt_365/$entry
      -- 	branch_block_stmt_365/branch_block_stmt_365__entry__
      -- 	branch_block_stmt_365/bb_0_bb_1
      -- 	branch_block_stmt_365/bb_0_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_365/bb_0_bb_1_PhiReq/$exit
      -- 
    -- CP-element group 1 transition  place  bypass 
    -- predecessors 
    -- successors 
    -- members (11) 
      -- 	$exit
      -- 	branch_block_stmt_365/$exit
      -- 	branch_block_stmt_365/branch_block_stmt_365__exit__
      -- 	branch_block_stmt_365/return__
      -- 	branch_block_stmt_365/merge_stmt_373__exit__
      -- 	branch_block_stmt_365/return___PhiReq/$entry
      -- 	branch_block_stmt_365/return___PhiReq/$exit
      -- 	branch_block_stmt_365/merge_stmt_373_PhiReqMerge
      -- 	branch_block_stmt_365/merge_stmt_373_PhiAck/$entry
      -- 	branch_block_stmt_365/merge_stmt_373_PhiAck/$exit
      -- 	branch_block_stmt_365/merge_stmt_373_PhiAck/dummy
      -- 
    cp_elements(1) <= false; 
    -- CP-element group 2 transition  input  output  no-bypass 
    -- predecessors 9 
    -- successors 3 
    -- members (5) 
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_active_
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_start/$exit
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_start/cra
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_complete/$entry
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_complete/ccr
      -- 
    cra_8569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_368_call_ack_0, ack => cp_elements(2)); -- 
    ccr_8573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_368_call_req_1); -- 
    -- CP-element group 3 transition  place  input  output  no-bypass 
    -- predecessors 2 
    -- successors 4 
    -- members (11) 
      -- 	branch_block_stmt_365/call_stmt_368__exit__
      -- 	branch_block_stmt_365/call_stmt_369__entry__
      -- 	branch_block_stmt_365/call_stmt_368/$exit
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_call_complete
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_completed_
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_complete/$exit
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_complete/cca
      -- 	branch_block_stmt_365/call_stmt_369/$entry
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_trigger_
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_start/$entry
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_start/crr
      -- 
    cca_8574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_368_call_ack_1, ack => cp_elements(3)); -- 
    crr_8585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => call_stmt_369_call_req_0); -- 
    -- CP-element group 4 transition  input  output  no-bypass 
    -- predecessors 3 
    -- successors 5 
    -- members (5) 
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_active_
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_start/$exit
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_start/cra
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_complete/$entry
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_complete/ccr
      -- 
    cra_8586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_369_call_ack_0, ack => cp_elements(4)); -- 
    ccr_8590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_369_call_req_1); -- 
    -- CP-element group 5 transition  place  input  output  no-bypass 
    -- predecessors 4 
    -- successors 6 
    -- members (11) 
      -- 	branch_block_stmt_365/call_stmt_369__exit__
      -- 	branch_block_stmt_365/call_stmt_370__entry__
      -- 	branch_block_stmt_365/call_stmt_369/$exit
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_call_complete
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_completed_
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_complete/$exit
      -- 	branch_block_stmt_365/call_stmt_369/call_stmt_369_complete/cca
      -- 	branch_block_stmt_365/call_stmt_370/$entry
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_trigger_
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_start/$entry
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_start/crr
      -- 
    cca_8591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_369_call_ack_1, ack => cp_elements(5)); -- 
    crr_8602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_370_call_req_0); -- 
    -- CP-element group 6 transition  input  output  no-bypass 
    -- predecessors 5 
    -- successors 7 
    -- members (5) 
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_active_
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_start/$exit
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_start/cra
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_complete/$entry
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_complete/ccr
      -- 
    cra_8603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_370_call_ack_0, ack => cp_elements(6)); -- 
    ccr_8607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => call_stmt_370_call_req_1); -- 
    -- CP-element group 7 transition  place  input  no-bypass 
    -- predecessors 6 
    -- successors 8 
    -- members (9) 
      -- 	branch_block_stmt_365/call_stmt_370__exit__
      -- 	branch_block_stmt_365/bb_1_bb_1
      -- 	branch_block_stmt_365/call_stmt_370/$exit
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_call_complete
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_completed_
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_complete/$exit
      -- 	branch_block_stmt_365/call_stmt_370/call_stmt_370_complete/cca
      -- 	branch_block_stmt_365/bb_1_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_365/bb_1_bb_1_PhiReq/$exit
      -- 
    cca_8608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_370_call_ack_1, ack => cp_elements(7)); -- 
    -- CP-element group 8 merge  place  bypass 
    -- predecessors 0 7 
    -- successors 9 
    -- members (1) 
      -- 	branch_block_stmt_365/merge_stmt_367_PhiReqMerge
      -- 
    cp_elements(8) <= OrReduce(cp_elements(0) & cp_elements(7));
    -- CP-element group 9 transition  place  output  bypass 
    -- predecessors 8 
    -- successors 2 
    -- members (9) 
      -- 	branch_block_stmt_365/merge_stmt_367__exit__
      -- 	branch_block_stmt_365/call_stmt_368__entry__
      -- 	branch_block_stmt_365/call_stmt_368/$entry
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_trigger_
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_start/$entry
      -- 	branch_block_stmt_365/call_stmt_368/call_stmt_368_start/crr
      -- 	branch_block_stmt_365/merge_stmt_367_PhiAck/$entry
      -- 	branch_block_stmt_365/merge_stmt_367_PhiAck/$exit
      -- 	branch_block_stmt_365/merge_stmt_367_PhiAck/dummy
      -- 
    cp_elements(9) <= cp_elements(8);
    crr_8568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => call_stmt_368_call_req_0); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    LogSplitOperator(clk,reset,global_clock_cycle_count,call_stmt_368_call_req_0,call_stmt_368_call_ack_0,call_stmt_368_call_req_1,call_stmt_368_call_ack_1,sl_one,"call_stmt_368_call",true, slv_zero,
    true, slv_zero);
    -- shared call operator group (0) : call_stmt_368_call 
    getData_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_368_call_req_0;
      call_stmt_368_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_368_call_req_1;
      call_stmt_368_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => getData_call_reqs(0),
          ackR => getData_call_acks(0),
          tagR => getData_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1, no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => getData_return_acks(0), -- cross-over
          ackL => getData_return_reqs(0), -- cross-over
          tagL => getData_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,call_stmt_369_call_req_0,call_stmt_369_call_ack_0,call_stmt_369_call_req_1,call_stmt_369_call_ack_1,sl_one,"call_stmt_369_call",true, slv_zero,
    true, slv_zero);
    -- shared call operator group (1) : call_stmt_369_call 
    x_vectorSum_x_call_group_1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_369_call_req_0;
      call_stmt_369_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_369_call_req_1;
      call_stmt_369_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => x_vectorSum_x_call_reqs(0),
          ackR => x_vectorSum_x_call_acks(0),
          tagR => x_vectorSum_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1, no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => x_vectorSum_x_return_acks(0), -- cross-over
          ackL => x_vectorSum_x_return_reqs(0), -- cross-over
          tagL => x_vectorSum_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,call_stmt_370_call_req_0,call_stmt_370_call_ack_0,call_stmt_370_call_req_1,call_stmt_370_call_ack_1,sl_one,"call_stmt_370_call",true, slv_zero,
    true, slv_zero);
    -- shared call operator group (2) : call_stmt_370_call 
    sendResult_call_group_2: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_370_call_req_0;
      call_stmt_370_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_370_call_req_1;
      call_stmt_370_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => sendResult_call_reqs(0),
          ackR => sendResult_call_acks(0),
          tagR => sendResult_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1, no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => sendResult_return_acks(0), -- cross-over
          ackL => sendResult_return_reqs(0), -- cross-over
          tagL => sendResult_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity x_vectorSum_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity x_vectorSum_x;
architecture Default of x_vectorSum_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal x_vectorSum_x_xCP_2164_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_512_base_resize_ack_0 : boolean;
  signal ptr_deref_529_base_resize_req_0 : boolean;
  signal ptr_deref_529_base_resize_ack_0 : boolean;
  signal binary_522_inst_req_0 : boolean;
  signal ptr_deref_512_load_0_ack_0 : boolean;
  signal ptr_deref_551_store_0_req_1 : boolean;
  signal binary_522_inst_ack_0 : boolean;
  signal binary_544_inst_req_1 : boolean;
  signal ptr_deref_639_store_0_ack_1 : boolean;
  signal ptr_deref_639_base_resize_req_0 : boolean;
  signal ptr_deref_644_base_resize_ack_0 : boolean;
  signal ptr_deref_529_gather_scatter_ack_0 : boolean;
  signal type_cast_648_inst_req_0 : boolean;
  signal ptr_deref_529_addr_0_req_0 : boolean;
  signal binary_544_inst_ack_0 : boolean;
  signal ptr_deref_512_root_address_inst_req_0 : boolean;
  signal ptr_deref_639_gather_scatter_ack_0 : boolean;
  signal ptr_deref_639_gather_scatter_req_0 : boolean;
  signal ptr_deref_534_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_652_index_0_resize_req_0 : boolean;
  signal binary_522_inst_ack_1 : boolean;
  signal ptr_deref_507_base_resize_req_0 : boolean;
  signal ptr_deref_507_base_resize_ack_0 : boolean;
  signal ptr_deref_507_root_address_inst_req_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal binary_522_inst_req_1 : boolean;
  signal ptr_deref_512_load_0_req_0 : boolean;
  signal ptr_deref_551_store_0_req_0 : boolean;
  signal ptr_deref_512_base_resize_req_0 : boolean;
  signal ptr_deref_512_load_0_req_1 : boolean;
  signal ptr_deref_507_gather_scatter_req_0 : boolean;
  signal ptr_deref_534_base_resize_ack_0 : boolean;
  signal ptr_deref_529_addr_0_ack_0 : boolean;
  signal ptr_deref_507_addr_0_ack_0 : boolean;
  signal ptr_deref_551_store_0_ack_1 : boolean;
  signal ptr_deref_529_store_0_ack_1 : boolean;
  signal ptr_deref_534_base_resize_req_0 : boolean;
  signal ptr_deref_551_base_resize_ack_0 : boolean;
  signal type_cast_526_inst_req_0 : boolean;
  signal ptr_deref_529_store_0_req_1 : boolean;
  signal ptr_deref_551_root_address_inst_req_0 : boolean;
  signal ptr_deref_644_load_0_ack_1 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal ptr_deref_534_load_0_req_0 : boolean;
  signal ptr_deref_512_addr_0_req_0 : boolean;
  signal array_obj_ref_652_index_0_resize_ack_0 : boolean;
  signal ptr_deref_644_root_address_inst_req_0 : boolean;
  signal ptr_deref_551_addr_0_req_0 : boolean;
  signal binary_544_inst_ack_1 : boolean;
  signal type_cast_648_inst_ack_0 : boolean;
  signal ptr_deref_512_addr_0_ack_0 : boolean;
  signal ptr_deref_644_root_address_inst_ack_0 : boolean;
  signal ptr_deref_534_load_0_req_1 : boolean;
  signal ptr_deref_534_load_0_ack_1 : boolean;
  signal ptr_deref_507_addr_0_req_0 : boolean;
  signal ptr_deref_534_addr_0_req_0 : boolean;
  signal ptr_deref_534_addr_0_ack_0 : boolean;
  signal ptr_deref_507_root_address_inst_ack_0 : boolean;
  signal ptr_deref_507_gather_scatter_ack_0 : boolean;
  signal ptr_deref_529_store_0_req_0 : boolean;
  signal ptr_deref_551_root_address_inst_ack_0 : boolean;
  signal type_cast_548_inst_req_0 : boolean;
  signal ptr_deref_551_store_0_ack_0 : boolean;
  signal ptr_deref_507_store_0_req_0 : boolean;
  signal ptr_deref_512_load_0_ack_1 : boolean;
  signal ptr_deref_512_gather_scatter_req_0 : boolean;
  signal ptr_deref_507_store_0_ack_0 : boolean;
  signal ptr_deref_512_gather_scatter_ack_0 : boolean;
  signal ptr_deref_529_store_0_ack_0 : boolean;
  signal ptr_deref_551_base_resize_req_0 : boolean;
  signal type_cast_526_inst_ack_0 : boolean;
  signal ptr_deref_534_gather_scatter_req_0 : boolean;
  signal type_cast_548_inst_ack_0 : boolean;
  signal ptr_deref_507_store_0_req_1 : boolean;
  signal ptr_deref_551_gather_scatter_req_0 : boolean;
  signal ptr_deref_507_store_0_ack_1 : boolean;
  signal ptr_deref_551_addr_0_ack_0 : boolean;
  signal ptr_deref_551_gather_scatter_ack_0 : boolean;
  signal ptr_deref_534_root_address_inst_req_0 : boolean;
  signal type_cast_516_inst_req_0 : boolean;
  signal ptr_deref_529_root_address_inst_req_0 : boolean;
  signal binary_544_inst_req_0 : boolean;
  signal ptr_deref_529_gather_scatter_req_0 : boolean;
  signal type_cast_516_inst_ack_0 : boolean;
  signal ptr_deref_534_root_address_inst_ack_0 : boolean;
  signal ptr_deref_529_root_address_inst_ack_0 : boolean;
  signal ptr_deref_512_root_address_inst_ack_0 : boolean;
  signal ptr_deref_534_load_0_ack_0 : boolean;
  signal ptr_deref_639_base_resize_ack_0 : boolean;
  signal array_obj_ref_652_root_address_inst_ack_0 : boolean;
  signal addr_of_653_final_reg_req_0 : boolean;
  signal ptr_deref_644_addr_0_req_0 : boolean;
  signal array_obj_ref_652_offset_inst_req_0 : boolean;
  signal addr_of_653_final_reg_ack_0 : boolean;
  signal ptr_deref_639_root_address_inst_req_0 : boolean;
  signal ptr_deref_644_addr_0_ack_0 : boolean;
  signal ptr_deref_639_root_address_inst_ack_0 : boolean;
  signal ptr_deref_459_base_resize_req_0 : boolean;
  signal ptr_deref_459_base_resize_ack_0 : boolean;
  signal ptr_deref_459_root_address_inst_req_0 : boolean;
  signal ptr_deref_459_root_address_inst_ack_0 : boolean;
  signal ptr_deref_459_addr_0_req_0 : boolean;
  signal ptr_deref_459_addr_0_ack_0 : boolean;
  signal array_obj_ref_652_index_0_rename_req_0 : boolean;
  signal ptr_deref_459_gather_scatter_req_0 : boolean;
  signal ptr_deref_459_gather_scatter_ack_0 : boolean;
  signal ptr_deref_459_store_0_req_0 : boolean;
  signal ptr_deref_459_store_0_ack_0 : boolean;
  signal ptr_deref_459_store_0_req_1 : boolean;
  signal ptr_deref_459_store_0_ack_1 : boolean;
  signal ptr_deref_644_gather_scatter_req_0 : boolean;
  signal ptr_deref_639_store_0_req_0 : boolean;
  signal ptr_deref_639_store_0_ack_0 : boolean;
  signal array_obj_ref_652_root_address_inst_req_0 : boolean;
  signal ptr_deref_467_base_resize_req_0 : boolean;
  signal ptr_deref_467_base_resize_ack_0 : boolean;
  signal array_obj_ref_652_index_0_rename_ack_0 : boolean;
  signal ptr_deref_467_root_address_inst_req_0 : boolean;
  signal ptr_deref_467_root_address_inst_ack_0 : boolean;
  signal ptr_deref_644_load_0_req_1 : boolean;
  signal ptr_deref_467_addr_0_req_0 : boolean;
  signal ptr_deref_467_addr_0_ack_0 : boolean;
  signal ptr_deref_639_addr_0_req_0 : boolean;
  signal ptr_deref_644_base_resize_req_0 : boolean;
  signal ptr_deref_467_load_0_req_0 : boolean;
  signal ptr_deref_467_load_0_ack_0 : boolean;
  signal ptr_deref_639_store_0_req_1 : boolean;
  signal ptr_deref_467_load_0_req_1 : boolean;
  signal ptr_deref_467_load_0_ack_1 : boolean;
  signal ptr_deref_467_gather_scatter_req_0 : boolean;
  signal ptr_deref_467_gather_scatter_ack_0 : boolean;
  signal ptr_deref_639_addr_0_ack_0 : boolean;
  signal ptr_deref_644_load_0_req_0 : boolean;
  signal ptr_deref_644_load_0_ack_0 : boolean;
  signal ptr_deref_644_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_652_offset_inst_ack_0 : boolean;
  signal type_cast_471_inst_req_0 : boolean;
  signal type_cast_471_inst_ack_0 : boolean;
  signal type_cast_475_inst_req_0 : boolean;
  signal type_cast_475_inst_ack_0 : boolean;
  signal binary_479_inst_req_0 : boolean;
  signal binary_479_inst_ack_0 : boolean;
  signal binary_479_inst_req_1 : boolean;
  signal binary_479_inst_ack_1 : boolean;
  signal if_stmt_481_branch_req_0 : boolean;
  signal if_stmt_481_branch_ack_1 : boolean;
  signal if_stmt_481_branch_ack_0 : boolean;
  signal ptr_deref_490_base_resize_req_0 : boolean;
  signal ptr_deref_490_base_resize_ack_0 : boolean;
  signal ptr_deref_490_root_address_inst_req_0 : boolean;
  signal ptr_deref_490_root_address_inst_ack_0 : boolean;
  signal ptr_deref_490_addr_0_req_0 : boolean;
  signal ptr_deref_490_addr_0_ack_0 : boolean;
  signal ptr_deref_490_load_0_req_0 : boolean;
  signal ptr_deref_490_load_0_ack_0 : boolean;
  signal ptr_deref_490_load_0_req_1 : boolean;
  signal ptr_deref_490_load_0_ack_1 : boolean;
  signal ptr_deref_490_gather_scatter_req_0 : boolean;
  signal ptr_deref_490_gather_scatter_ack_0 : boolean;
  signal type_cast_494_inst_req_0 : boolean;
  signal type_cast_494_inst_ack_0 : boolean;
  signal binary_500_inst_req_0 : boolean;
  signal binary_500_inst_ack_0 : boolean;
  signal binary_500_inst_req_1 : boolean;
  signal binary_500_inst_ack_1 : boolean;
  signal type_cast_504_inst_req_0 : boolean;
  signal type_cast_504_inst_ack_0 : boolean;
  signal ptr_deref_556_base_resize_req_0 : boolean;
  signal ptr_deref_556_base_resize_ack_0 : boolean;
  signal ptr_deref_556_root_address_inst_req_0 : boolean;
  signal ptr_deref_556_root_address_inst_ack_0 : boolean;
  signal ptr_deref_556_addr_0_req_0 : boolean;
  signal ptr_deref_556_addr_0_ack_0 : boolean;
  signal ptr_deref_556_load_0_req_0 : boolean;
  signal ptr_deref_556_load_0_ack_0 : boolean;
  signal ptr_deref_556_load_0_req_1 : boolean;
  signal ptr_deref_556_load_0_ack_1 : boolean;
  signal ptr_deref_556_gather_scatter_req_0 : boolean;
  signal ptr_deref_556_gather_scatter_ack_0 : boolean;
  signal type_cast_560_inst_req_0 : boolean;
  signal type_cast_560_inst_ack_0 : boolean;
  signal binary_566_inst_req_0 : boolean;
  signal binary_566_inst_ack_0 : boolean;
  signal binary_566_inst_req_1 : boolean;
  signal binary_566_inst_ack_1 : boolean;
  signal type_cast_570_inst_req_0 : boolean;
  signal type_cast_570_inst_ack_0 : boolean;
  signal ptr_deref_786_base_resize_req_0 : boolean;
  signal ptr_deref_573_base_resize_req_0 : boolean;
  signal ptr_deref_573_base_resize_ack_0 : boolean;
  signal ptr_deref_773_load_0_req_1 : boolean;
  signal ptr_deref_573_root_address_inst_req_0 : boolean;
  signal ptr_deref_573_root_address_inst_ack_0 : boolean;
  signal ptr_deref_573_addr_0_req_0 : boolean;
  signal ptr_deref_573_addr_0_ack_0 : boolean;
  signal ptr_deref_573_gather_scatter_req_0 : boolean;
  signal ptr_deref_573_gather_scatter_ack_0 : boolean;
  signal ptr_deref_573_store_0_req_0 : boolean;
  signal ptr_deref_573_store_0_ack_0 : boolean;
  signal ptr_deref_773_load_0_ack_1 : boolean;
  signal ptr_deref_573_store_0_req_1 : boolean;
  signal ptr_deref_573_store_0_ack_1 : boolean;
  signal ptr_deref_773_gather_scatter_req_0 : boolean;
  signal ptr_deref_578_base_resize_req_0 : boolean;
  signal ptr_deref_578_base_resize_ack_0 : boolean;
  signal ptr_deref_578_root_address_inst_req_0 : boolean;
  signal ptr_deref_578_root_address_inst_ack_0 : boolean;
  signal ptr_deref_578_addr_0_req_0 : boolean;
  signal ptr_deref_578_addr_0_ack_0 : boolean;
  signal addr_of_782_final_reg_req_0 : boolean;
  signal addr_of_782_final_reg_ack_0 : boolean;
  signal ptr_deref_578_load_0_req_0 : boolean;
  signal ptr_deref_578_load_0_ack_0 : boolean;
  signal ptr_deref_773_gather_scatter_ack_0 : boolean;
  signal ptr_deref_578_load_0_req_1 : boolean;
  signal ptr_deref_578_load_0_ack_1 : boolean;
  signal ptr_deref_578_gather_scatter_req_0 : boolean;
  signal ptr_deref_578_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_781_root_address_inst_req_0 : boolean;
  signal type_cast_582_inst_req_0 : boolean;
  signal type_cast_582_inst_ack_0 : boolean;
  signal array_obj_ref_781_index_0_resize_req_0 : boolean;
  signal binary_588_inst_req_0 : boolean;
  signal binary_588_inst_ack_0 : boolean;
  signal binary_588_inst_req_1 : boolean;
  signal binary_588_inst_ack_1 : boolean;
  signal ptr_deref_786_root_address_inst_req_0 : boolean;
  signal ptr_deref_786_root_address_inst_ack_0 : boolean;
  signal ptr_deref_773_base_resize_req_0 : boolean;
  signal array_obj_ref_781_offset_inst_req_0 : boolean;
  signal ptr_deref_773_base_resize_ack_0 : boolean;
  signal type_cast_592_inst_req_0 : boolean;
  signal type_cast_592_inst_ack_0 : boolean;
  signal array_obj_ref_781_index_0_resize_ack_0 : boolean;
  signal ptr_deref_773_root_address_inst_req_0 : boolean;
  signal array_obj_ref_781_offset_inst_ack_0 : boolean;
  signal ptr_deref_773_root_address_inst_ack_0 : boolean;
  signal ptr_deref_595_base_resize_req_0 : boolean;
  signal ptr_deref_595_base_resize_ack_0 : boolean;
  signal ptr_deref_595_root_address_inst_req_0 : boolean;
  signal ptr_deref_595_root_address_inst_ack_0 : boolean;
  signal ptr_deref_595_addr_0_req_0 : boolean;
  signal ptr_deref_595_addr_0_ack_0 : boolean;
  signal ptr_deref_595_gather_scatter_req_0 : boolean;
  signal ptr_deref_595_gather_scatter_ack_0 : boolean;
  signal ptr_deref_595_store_0_req_0 : boolean;
  signal ptr_deref_595_store_0_ack_0 : boolean;
  signal ptr_deref_595_store_0_req_1 : boolean;
  signal ptr_deref_595_store_0_ack_1 : boolean;
  signal array_obj_ref_781_root_address_inst_ack_0 : boolean;
  signal ptr_deref_773_addr_0_req_0 : boolean;
  signal ptr_deref_786_base_resize_ack_0 : boolean;
  signal type_cast_777_inst_req_0 : boolean;
  signal ptr_deref_773_addr_0_ack_0 : boolean;
  signal ptr_deref_600_base_resize_req_0 : boolean;
  signal ptr_deref_600_base_resize_ack_0 : boolean;
  signal ptr_deref_600_root_address_inst_req_0 : boolean;
  signal ptr_deref_600_root_address_inst_ack_0 : boolean;
  signal ptr_deref_600_addr_0_req_0 : boolean;
  signal ptr_deref_600_addr_0_ack_0 : boolean;
  signal type_cast_777_inst_ack_0 : boolean;
  signal ptr_deref_600_load_0_req_0 : boolean;
  signal ptr_deref_600_load_0_ack_0 : boolean;
  signal ptr_deref_600_load_0_req_1 : boolean;
  signal ptr_deref_600_load_0_ack_1 : boolean;
  signal ptr_deref_600_gather_scatter_req_0 : boolean;
  signal ptr_deref_600_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_781_index_0_rename_req_0 : boolean;
  signal ptr_deref_773_load_0_req_0 : boolean;
  signal ptr_deref_773_load_0_ack_0 : boolean;
  signal array_obj_ref_781_index_0_rename_ack_0 : boolean;
  signal type_cast_604_inst_req_0 : boolean;
  signal type_cast_604_inst_ack_0 : boolean;
  signal binary_610_inst_req_0 : boolean;
  signal binary_610_inst_ack_0 : boolean;
  signal binary_610_inst_req_1 : boolean;
  signal binary_610_inst_ack_1 : boolean;
  signal type_cast_614_inst_req_0 : boolean;
  signal type_cast_614_inst_ack_0 : boolean;
  signal ptr_deref_617_base_resize_req_0 : boolean;
  signal ptr_deref_617_base_resize_ack_0 : boolean;
  signal ptr_deref_617_root_address_inst_req_0 : boolean;
  signal ptr_deref_617_root_address_inst_ack_0 : boolean;
  signal ptr_deref_617_addr_0_req_0 : boolean;
  signal ptr_deref_617_addr_0_ack_0 : boolean;
  signal ptr_deref_617_gather_scatter_req_0 : boolean;
  signal ptr_deref_617_gather_scatter_ack_0 : boolean;
  signal ptr_deref_617_store_0_req_0 : boolean;
  signal ptr_deref_617_store_0_ack_0 : boolean;
  signal ptr_deref_617_store_0_req_1 : boolean;
  signal ptr_deref_617_store_0_ack_1 : boolean;
  signal ptr_deref_622_base_resize_req_0 : boolean;
  signal ptr_deref_622_base_resize_ack_0 : boolean;
  signal ptr_deref_622_root_address_inst_req_0 : boolean;
  signal ptr_deref_622_root_address_inst_ack_0 : boolean;
  signal ptr_deref_622_addr_0_req_0 : boolean;
  signal ptr_deref_622_addr_0_ack_0 : boolean;
  signal ptr_deref_622_load_0_req_0 : boolean;
  signal ptr_deref_622_load_0_ack_0 : boolean;
  signal ptr_deref_622_load_0_req_1 : boolean;
  signal ptr_deref_622_load_0_ack_1 : boolean;
  signal ptr_deref_622_gather_scatter_req_0 : boolean;
  signal ptr_deref_622_gather_scatter_ack_0 : boolean;
  signal type_cast_626_inst_req_0 : boolean;
  signal type_cast_626_inst_ack_0 : boolean;
  signal binary_632_inst_req_0 : boolean;
  signal binary_632_inst_ack_0 : boolean;
  signal binary_632_inst_req_1 : boolean;
  signal binary_632_inst_ack_1 : boolean;
  signal type_cast_636_inst_req_0 : boolean;
  signal type_cast_636_inst_ack_0 : boolean;
  signal ptr_deref_786_addr_0_req_0 : boolean;
  signal ptr_deref_786_addr_0_ack_0 : boolean;
  signal ptr_deref_657_base_resize_req_0 : boolean;
  signal ptr_deref_657_base_resize_ack_0 : boolean;
  signal ptr_deref_657_root_address_inst_req_0 : boolean;
  signal ptr_deref_657_root_address_inst_ack_0 : boolean;
  signal ptr_deref_657_addr_0_req_0 : boolean;
  signal ptr_deref_657_addr_0_ack_0 : boolean;
  signal ptr_deref_657_load_0_req_0 : boolean;
  signal ptr_deref_657_load_0_ack_0 : boolean;
  signal ptr_deref_657_load_0_req_1 : boolean;
  signal ptr_deref_657_load_0_ack_1 : boolean;
  signal ptr_deref_657_gather_scatter_req_0 : boolean;
  signal ptr_deref_657_gather_scatter_ack_0 : boolean;
  signal ptr_deref_661_base_resize_req_0 : boolean;
  signal ptr_deref_661_base_resize_ack_0 : boolean;
  signal ptr_deref_661_root_address_inst_req_0 : boolean;
  signal ptr_deref_661_root_address_inst_ack_0 : boolean;
  signal ptr_deref_661_addr_0_req_0 : boolean;
  signal ptr_deref_661_addr_0_ack_0 : boolean;
  signal ptr_deref_661_load_0_req_0 : boolean;
  signal ptr_deref_661_load_0_ack_0 : boolean;
  signal ptr_deref_661_load_0_req_1 : boolean;
  signal ptr_deref_661_load_0_ack_1 : boolean;
  signal ptr_deref_661_gather_scatter_req_0 : boolean;
  signal ptr_deref_661_gather_scatter_ack_0 : boolean;
  signal type_cast_665_inst_req_0 : boolean;
  signal type_cast_665_inst_ack_0 : boolean;
  signal array_obj_ref_669_index_0_resize_req_0 : boolean;
  signal array_obj_ref_669_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_669_index_0_rename_req_0 : boolean;
  signal array_obj_ref_669_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_669_offset_inst_req_0 : boolean;
  signal array_obj_ref_669_offset_inst_ack_0 : boolean;
  signal array_obj_ref_669_root_address_inst_req_0 : boolean;
  signal array_obj_ref_669_root_address_inst_ack_0 : boolean;
  signal addr_of_670_final_reg_req_0 : boolean;
  signal addr_of_670_final_reg_ack_0 : boolean;
  signal ptr_deref_674_base_resize_req_0 : boolean;
  signal ptr_deref_674_base_resize_ack_0 : boolean;
  signal ptr_deref_674_root_address_inst_req_0 : boolean;
  signal ptr_deref_674_root_address_inst_ack_0 : boolean;
  signal ptr_deref_674_addr_0_req_0 : boolean;
  signal ptr_deref_674_addr_0_ack_0 : boolean;
  signal ptr_deref_674_load_0_req_0 : boolean;
  signal ptr_deref_674_load_0_ack_0 : boolean;
  signal ptr_deref_674_load_0_req_1 : boolean;
  signal ptr_deref_674_load_0_ack_1 : boolean;
  signal ptr_deref_674_gather_scatter_req_0 : boolean;
  signal ptr_deref_674_gather_scatter_ack_0 : boolean;
  signal binary_679_inst_req_0 : boolean;
  signal binary_679_inst_ack_0 : boolean;
  signal binary_679_inst_req_1 : boolean;
  signal binary_679_inst_ack_1 : boolean;
  signal ptr_deref_682_base_resize_req_0 : boolean;
  signal ptr_deref_682_base_resize_ack_0 : boolean;
  signal ptr_deref_682_root_address_inst_req_0 : boolean;
  signal ptr_deref_682_root_address_inst_ack_0 : boolean;
  signal ptr_deref_682_addr_0_req_0 : boolean;
  signal ptr_deref_682_addr_0_ack_0 : boolean;
  signal ptr_deref_682_gather_scatter_req_0 : boolean;
  signal ptr_deref_682_gather_scatter_ack_0 : boolean;
  signal ptr_deref_682_store_0_req_0 : boolean;
  signal ptr_deref_682_store_0_ack_0 : boolean;
  signal ptr_deref_682_store_0_req_1 : boolean;
  signal ptr_deref_682_store_0_ack_1 : boolean;
  signal ptr_deref_687_base_resize_req_0 : boolean;
  signal ptr_deref_687_base_resize_ack_0 : boolean;
  signal ptr_deref_687_root_address_inst_req_0 : boolean;
  signal ptr_deref_687_root_address_inst_ack_0 : boolean;
  signal ptr_deref_687_addr_0_req_0 : boolean;
  signal ptr_deref_687_addr_0_ack_0 : boolean;
  signal ptr_deref_687_load_0_req_0 : boolean;
  signal ptr_deref_687_load_0_ack_0 : boolean;
  signal ptr_deref_687_load_0_req_1 : boolean;
  signal ptr_deref_687_load_0_ack_1 : boolean;
  signal ptr_deref_687_gather_scatter_req_0 : boolean;
  signal ptr_deref_687_gather_scatter_ack_0 : boolean;
  signal type_cast_691_inst_req_0 : boolean;
  signal type_cast_691_inst_ack_0 : boolean;
  signal ptr_deref_889_addr_0_ack_0 : boolean;
  signal array_obj_ref_695_index_0_resize_req_0 : boolean;
  signal array_obj_ref_695_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_695_index_0_rename_req_0 : boolean;
  signal array_obj_ref_695_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_695_offset_inst_req_0 : boolean;
  signal array_obj_ref_695_offset_inst_ack_0 : boolean;
  signal array_obj_ref_695_root_address_inst_req_0 : boolean;
  signal array_obj_ref_695_root_address_inst_ack_0 : boolean;
  signal addr_of_696_final_reg_req_0 : boolean;
  signal addr_of_696_final_reg_ack_0 : boolean;
  signal ptr_deref_700_base_resize_req_0 : boolean;
  signal ptr_deref_700_base_resize_ack_0 : boolean;
  signal ptr_deref_700_root_address_inst_req_0 : boolean;
  signal ptr_deref_700_root_address_inst_ack_0 : boolean;
  signal ptr_deref_700_addr_0_req_0 : boolean;
  signal ptr_deref_700_addr_0_ack_0 : boolean;
  signal ptr_deref_700_load_0_req_0 : boolean;
  signal ptr_deref_700_load_0_ack_0 : boolean;
  signal ptr_deref_700_load_0_req_1 : boolean;
  signal ptr_deref_700_load_0_ack_1 : boolean;
  signal ptr_deref_700_gather_scatter_req_0 : boolean;
  signal ptr_deref_700_gather_scatter_ack_0 : boolean;
  signal ptr_deref_704_base_resize_req_0 : boolean;
  signal ptr_deref_704_base_resize_ack_0 : boolean;
  signal ptr_deref_704_root_address_inst_req_0 : boolean;
  signal ptr_deref_704_root_address_inst_ack_0 : boolean;
  signal ptr_deref_704_addr_0_req_0 : boolean;
  signal ptr_deref_704_addr_0_ack_0 : boolean;
  signal ptr_deref_704_load_0_req_0 : boolean;
  signal ptr_deref_704_load_0_ack_0 : boolean;
  signal ptr_deref_704_load_0_req_1 : boolean;
  signal ptr_deref_704_load_0_ack_1 : boolean;
  signal ptr_deref_704_gather_scatter_req_0 : boolean;
  signal ptr_deref_704_gather_scatter_ack_0 : boolean;
  signal ptr_deref_889_load_0_req_0 : boolean;
  signal ptr_deref_889_load_0_ack_0 : boolean;
  signal type_cast_708_inst_req_0 : boolean;
  signal type_cast_708_inst_ack_0 : boolean;
  signal ptr_deref_889_base_resize_req_0 : boolean;
  signal ptr_deref_889_base_resize_ack_0 : boolean;
  signal array_obj_ref_712_index_0_resize_req_0 : boolean;
  signal array_obj_ref_712_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_712_index_0_rename_req_0 : boolean;
  signal array_obj_ref_712_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_712_offset_inst_req_0 : boolean;
  signal array_obj_ref_712_offset_inst_ack_0 : boolean;
  signal array_obj_ref_712_root_address_inst_req_0 : boolean;
  signal array_obj_ref_712_root_address_inst_ack_0 : boolean;
  signal addr_of_713_final_reg_req_0 : boolean;
  signal addr_of_713_final_reg_ack_0 : boolean;
  signal ptr_deref_889_gather_scatter_ack_0 : boolean;
  signal ptr_deref_889_root_address_inst_req_0 : boolean;
  signal ptr_deref_889_root_address_inst_ack_0 : boolean;
  signal ptr_deref_889_load_0_req_1 : boolean;
  signal ptr_deref_889_load_0_ack_1 : boolean;
  signal ptr_deref_889_addr_0_req_0 : boolean;
  signal ptr_deref_889_gather_scatter_req_0 : boolean;
  signal ptr_deref_717_base_resize_req_0 : boolean;
  signal ptr_deref_717_base_resize_ack_0 : boolean;
  signal ptr_deref_717_root_address_inst_req_0 : boolean;
  signal ptr_deref_717_root_address_inst_ack_0 : boolean;
  signal ptr_deref_717_addr_0_req_0 : boolean;
  signal ptr_deref_717_addr_0_ack_0 : boolean;
  signal ptr_deref_717_load_0_req_0 : boolean;
  signal ptr_deref_717_load_0_ack_0 : boolean;
  signal ptr_deref_717_load_0_req_1 : boolean;
  signal ptr_deref_717_load_0_ack_1 : boolean;
  signal ptr_deref_717_gather_scatter_req_0 : boolean;
  signal ptr_deref_717_gather_scatter_ack_0 : boolean;
  signal binary_722_inst_req_0 : boolean;
  signal binary_722_inst_ack_0 : boolean;
  signal binary_722_inst_req_1 : boolean;
  signal binary_722_inst_ack_1 : boolean;
  signal ptr_deref_725_base_resize_req_0 : boolean;
  signal ptr_deref_725_base_resize_ack_0 : boolean;
  signal ptr_deref_725_root_address_inst_req_0 : boolean;
  signal ptr_deref_725_root_address_inst_ack_0 : boolean;
  signal ptr_deref_725_addr_0_req_0 : boolean;
  signal ptr_deref_725_addr_0_ack_0 : boolean;
  signal ptr_deref_725_gather_scatter_req_0 : boolean;
  signal ptr_deref_725_gather_scatter_ack_0 : boolean;
  signal ptr_deref_725_store_0_req_0 : boolean;
  signal ptr_deref_725_store_0_ack_0 : boolean;
  signal ptr_deref_725_store_0_req_1 : boolean;
  signal ptr_deref_725_store_0_ack_1 : boolean;
  signal ptr_deref_730_base_resize_req_0 : boolean;
  signal ptr_deref_730_base_resize_ack_0 : boolean;
  signal ptr_deref_730_root_address_inst_req_0 : boolean;
  signal ptr_deref_730_root_address_inst_ack_0 : boolean;
  signal ptr_deref_730_addr_0_req_0 : boolean;
  signal ptr_deref_730_addr_0_ack_0 : boolean;
  signal ptr_deref_730_load_0_req_0 : boolean;
  signal ptr_deref_730_load_0_ack_0 : boolean;
  signal ptr_deref_730_load_0_req_1 : boolean;
  signal ptr_deref_730_load_0_ack_1 : boolean;
  signal ptr_deref_730_gather_scatter_req_0 : boolean;
  signal ptr_deref_730_gather_scatter_ack_0 : boolean;
  signal type_cast_734_inst_req_0 : boolean;
  signal type_cast_734_inst_ack_0 : boolean;
  signal array_obj_ref_738_index_0_resize_req_0 : boolean;
  signal array_obj_ref_738_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_738_index_0_rename_req_0 : boolean;
  signal array_obj_ref_738_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_738_offset_inst_req_0 : boolean;
  signal array_obj_ref_738_offset_inst_ack_0 : boolean;
  signal array_obj_ref_738_root_address_inst_req_0 : boolean;
  signal array_obj_ref_738_root_address_inst_ack_0 : boolean;
  signal addr_of_739_final_reg_req_0 : boolean;
  signal addr_of_739_final_reg_ack_0 : boolean;
  signal ptr_deref_743_base_resize_req_0 : boolean;
  signal ptr_deref_743_base_resize_ack_0 : boolean;
  signal ptr_deref_743_root_address_inst_req_0 : boolean;
  signal ptr_deref_743_root_address_inst_ack_0 : boolean;
  signal ptr_deref_743_addr_0_req_0 : boolean;
  signal ptr_deref_743_addr_0_ack_0 : boolean;
  signal ptr_deref_743_load_0_req_0 : boolean;
  signal ptr_deref_743_load_0_ack_0 : boolean;
  signal ptr_deref_743_load_0_req_1 : boolean;
  signal ptr_deref_743_load_0_ack_1 : boolean;
  signal ptr_deref_743_gather_scatter_req_0 : boolean;
  signal ptr_deref_743_gather_scatter_ack_0 : boolean;
  signal ptr_deref_747_base_resize_req_0 : boolean;
  signal ptr_deref_747_base_resize_ack_0 : boolean;
  signal ptr_deref_747_root_address_inst_req_0 : boolean;
  signal ptr_deref_747_root_address_inst_ack_0 : boolean;
  signal ptr_deref_747_addr_0_req_0 : boolean;
  signal ptr_deref_747_addr_0_ack_0 : boolean;
  signal ptr_deref_747_load_0_req_0 : boolean;
  signal ptr_deref_747_load_0_ack_0 : boolean;
  signal ptr_deref_747_load_0_req_1 : boolean;
  signal ptr_deref_747_load_0_ack_1 : boolean;
  signal ptr_deref_747_gather_scatter_req_0 : boolean;
  signal ptr_deref_747_gather_scatter_ack_0 : boolean;
  signal type_cast_751_inst_req_0 : boolean;
  signal type_cast_751_inst_ack_0 : boolean;
  signal array_obj_ref_755_index_0_resize_req_0 : boolean;
  signal array_obj_ref_755_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_755_index_0_rename_req_0 : boolean;
  signal array_obj_ref_755_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_755_offset_inst_req_0 : boolean;
  signal array_obj_ref_755_offset_inst_ack_0 : boolean;
  signal array_obj_ref_755_root_address_inst_req_0 : boolean;
  signal array_obj_ref_755_root_address_inst_ack_0 : boolean;
  signal addr_of_756_final_reg_req_0 : boolean;
  signal addr_of_756_final_reg_ack_0 : boolean;
  signal ptr_deref_760_base_resize_req_0 : boolean;
  signal ptr_deref_760_base_resize_ack_0 : boolean;
  signal ptr_deref_760_root_address_inst_req_0 : boolean;
  signal ptr_deref_760_root_address_inst_ack_0 : boolean;
  signal ptr_deref_760_addr_0_req_0 : boolean;
  signal ptr_deref_760_addr_0_ack_0 : boolean;
  signal ptr_deref_760_load_0_req_0 : boolean;
  signal ptr_deref_760_load_0_ack_0 : boolean;
  signal ptr_deref_760_load_0_req_1 : boolean;
  signal ptr_deref_760_load_0_ack_1 : boolean;
  signal ptr_deref_760_gather_scatter_req_0 : boolean;
  signal ptr_deref_760_gather_scatter_ack_0 : boolean;
  signal binary_765_inst_req_0 : boolean;
  signal binary_765_inst_ack_0 : boolean;
  signal binary_765_inst_req_1 : boolean;
  signal binary_765_inst_ack_1 : boolean;
  signal ptr_deref_768_base_resize_req_0 : boolean;
  signal ptr_deref_768_base_resize_ack_0 : boolean;
  signal ptr_deref_768_root_address_inst_req_0 : boolean;
  signal ptr_deref_768_root_address_inst_ack_0 : boolean;
  signal ptr_deref_768_addr_0_req_0 : boolean;
  signal ptr_deref_768_addr_0_ack_0 : boolean;
  signal ptr_deref_768_gather_scatter_req_0 : boolean;
  signal ptr_deref_768_gather_scatter_ack_0 : boolean;
  signal ptr_deref_768_store_0_req_0 : boolean;
  signal ptr_deref_768_store_0_ack_0 : boolean;
  signal ptr_deref_768_store_0_req_1 : boolean;
  signal ptr_deref_768_store_0_ack_1 : boolean;
  signal ptr_deref_1051_gather_scatter_ack_0 : boolean;
  signal ptr_deref_786_load_0_req_0 : boolean;
  signal ptr_deref_786_load_0_ack_0 : boolean;
  signal ptr_deref_786_load_0_req_1 : boolean;
  signal ptr_deref_786_load_0_ack_1 : boolean;
  signal ptr_deref_786_gather_scatter_req_0 : boolean;
  signal ptr_deref_786_gather_scatter_ack_0 : boolean;
  signal ptr_deref_790_base_resize_req_0 : boolean;
  signal ptr_deref_790_base_resize_ack_0 : boolean;
  signal ptr_deref_790_root_address_inst_req_0 : boolean;
  signal ptr_deref_790_root_address_inst_ack_0 : boolean;
  signal ptr_deref_790_addr_0_req_0 : boolean;
  signal ptr_deref_790_addr_0_ack_0 : boolean;
  signal ptr_deref_790_load_0_req_0 : boolean;
  signal ptr_deref_790_load_0_ack_0 : boolean;
  signal ptr_deref_790_load_0_req_1 : boolean;
  signal ptr_deref_790_load_0_ack_1 : boolean;
  signal ptr_deref_790_gather_scatter_req_0 : boolean;
  signal ptr_deref_790_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1034_gather_scatter_ack_0 : boolean;
  signal type_cast_794_inst_req_0 : boolean;
  signal type_cast_794_inst_ack_0 : boolean;
  signal type_cast_1038_inst_ack_0 : boolean;
  signal array_obj_ref_798_index_0_resize_req_0 : boolean;
  signal array_obj_ref_798_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_798_index_0_rename_req_0 : boolean;
  signal array_obj_ref_798_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_798_offset_inst_req_0 : boolean;
  signal array_obj_ref_798_offset_inst_ack_0 : boolean;
  signal array_obj_ref_798_root_address_inst_req_0 : boolean;
  signal array_obj_ref_798_root_address_inst_ack_0 : boolean;
  signal addr_of_799_final_reg_req_0 : boolean;
  signal addr_of_799_final_reg_ack_0 : boolean;
  signal ptr_deref_1030_load_0_ack_0 : boolean;
  signal ptr_deref_803_base_resize_req_0 : boolean;
  signal ptr_deref_803_base_resize_ack_0 : boolean;
  signal ptr_deref_803_root_address_inst_req_0 : boolean;
  signal ptr_deref_803_root_address_inst_ack_0 : boolean;
  signal ptr_deref_803_addr_0_req_0 : boolean;
  signal ptr_deref_803_addr_0_ack_0 : boolean;
  signal ptr_deref_803_load_0_req_0 : boolean;
  signal ptr_deref_803_load_0_ack_0 : boolean;
  signal ptr_deref_803_load_0_req_1 : boolean;
  signal ptr_deref_803_load_0_ack_1 : boolean;
  signal ptr_deref_803_gather_scatter_req_0 : boolean;
  signal ptr_deref_803_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1034_base_resize_ack_0 : boolean;
  signal ptr_deref_1034_base_resize_req_0 : boolean;
  signal binary_808_inst_req_0 : boolean;
  signal binary_808_inst_ack_0 : boolean;
  signal binary_808_inst_req_1 : boolean;
  signal binary_808_inst_ack_1 : boolean;
  signal ptr_deref_988_load_0_req_1 : boolean;
  signal ptr_deref_988_load_0_ack_1 : boolean;
  signal ptr_deref_1034_gather_scatter_req_0 : boolean;
  signal ptr_deref_811_base_resize_req_0 : boolean;
  signal ptr_deref_811_base_resize_ack_0 : boolean;
  signal ptr_deref_811_root_address_inst_req_0 : boolean;
  signal ptr_deref_811_root_address_inst_ack_0 : boolean;
  signal ptr_deref_811_addr_0_req_0 : boolean;
  signal ptr_deref_811_addr_0_ack_0 : boolean;
  signal ptr_deref_811_gather_scatter_req_0 : boolean;
  signal ptr_deref_811_gather_scatter_ack_0 : boolean;
  signal ptr_deref_811_store_0_req_0 : boolean;
  signal ptr_deref_811_store_0_ack_0 : boolean;
  signal ptr_deref_811_store_0_req_1 : boolean;
  signal ptr_deref_811_store_0_ack_1 : boolean;
  signal ptr_deref_992_base_resize_ack_0 : boolean;
  signal ptr_deref_988_gather_scatter_req_0 : boolean;
  signal ptr_deref_816_base_resize_req_0 : boolean;
  signal ptr_deref_816_base_resize_ack_0 : boolean;
  signal ptr_deref_988_gather_scatter_ack_0 : boolean;
  signal ptr_deref_816_root_address_inst_req_0 : boolean;
  signal ptr_deref_816_root_address_inst_ack_0 : boolean;
  signal ptr_deref_992_base_resize_req_0 : boolean;
  signal ptr_deref_816_addr_0_req_0 : boolean;
  signal ptr_deref_816_addr_0_ack_0 : boolean;
  signal ptr_deref_816_load_0_req_0 : boolean;
  signal ptr_deref_816_load_0_ack_0 : boolean;
  signal ptr_deref_816_load_0_req_1 : boolean;
  signal ptr_deref_816_load_0_ack_1 : boolean;
  signal ptr_deref_816_gather_scatter_req_0 : boolean;
  signal ptr_deref_816_gather_scatter_ack_0 : boolean;
  signal type_cast_820_inst_req_0 : boolean;
  signal type_cast_820_inst_ack_0 : boolean;
  signal array_obj_ref_824_index_0_resize_req_0 : boolean;
  signal array_obj_ref_824_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_824_index_0_rename_req_0 : boolean;
  signal array_obj_ref_824_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_824_offset_inst_req_0 : boolean;
  signal array_obj_ref_824_offset_inst_ack_0 : boolean;
  signal array_obj_ref_824_root_address_inst_req_0 : boolean;
  signal array_obj_ref_824_root_address_inst_ack_0 : boolean;
  signal addr_of_825_final_reg_req_0 : boolean;
  signal addr_of_825_final_reg_ack_0 : boolean;
  signal ptr_deref_829_base_resize_req_0 : boolean;
  signal ptr_deref_829_base_resize_ack_0 : boolean;
  signal ptr_deref_829_root_address_inst_req_0 : boolean;
  signal ptr_deref_829_root_address_inst_ack_0 : boolean;
  signal ptr_deref_829_addr_0_req_0 : boolean;
  signal ptr_deref_829_addr_0_ack_0 : boolean;
  signal ptr_deref_829_load_0_req_0 : boolean;
  signal ptr_deref_829_load_0_ack_0 : boolean;
  signal ptr_deref_829_load_0_req_1 : boolean;
  signal ptr_deref_829_load_0_ack_1 : boolean;
  signal ptr_deref_829_gather_scatter_req_0 : boolean;
  signal ptr_deref_829_gather_scatter_ack_0 : boolean;
  signal ptr_deref_833_base_resize_req_0 : boolean;
  signal ptr_deref_833_base_resize_ack_0 : boolean;
  signal ptr_deref_833_root_address_inst_req_0 : boolean;
  signal ptr_deref_833_root_address_inst_ack_0 : boolean;
  signal ptr_deref_833_addr_0_req_0 : boolean;
  signal ptr_deref_833_addr_0_ack_0 : boolean;
  signal ptr_deref_833_load_0_req_0 : boolean;
  signal ptr_deref_833_load_0_ack_0 : boolean;
  signal ptr_deref_833_load_0_req_1 : boolean;
  signal ptr_deref_833_load_0_ack_1 : boolean;
  signal ptr_deref_833_gather_scatter_req_0 : boolean;
  signal ptr_deref_833_gather_scatter_ack_0 : boolean;
  signal type_cast_837_inst_req_0 : boolean;
  signal type_cast_837_inst_ack_0 : boolean;
  signal array_obj_ref_841_index_0_resize_req_0 : boolean;
  signal array_obj_ref_841_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_841_index_0_rename_req_0 : boolean;
  signal array_obj_ref_841_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_841_offset_inst_req_0 : boolean;
  signal array_obj_ref_841_offset_inst_ack_0 : boolean;
  signal array_obj_ref_841_root_address_inst_req_0 : boolean;
  signal array_obj_ref_841_root_address_inst_ack_0 : boolean;
  signal addr_of_842_final_reg_req_0 : boolean;
  signal addr_of_842_final_reg_ack_0 : boolean;
  signal ptr_deref_846_base_resize_req_0 : boolean;
  signal ptr_deref_846_base_resize_ack_0 : boolean;
  signal ptr_deref_846_root_address_inst_req_0 : boolean;
  signal ptr_deref_846_root_address_inst_ack_0 : boolean;
  signal ptr_deref_846_addr_0_req_0 : boolean;
  signal ptr_deref_846_addr_0_ack_0 : boolean;
  signal ptr_deref_846_load_0_req_0 : boolean;
  signal ptr_deref_846_load_0_ack_0 : boolean;
  signal ptr_deref_846_load_0_req_1 : boolean;
  signal ptr_deref_846_load_0_ack_1 : boolean;
  signal ptr_deref_846_gather_scatter_req_0 : boolean;
  signal ptr_deref_846_gather_scatter_ack_0 : boolean;
  signal binary_851_inst_req_0 : boolean;
  signal binary_851_inst_ack_0 : boolean;
  signal binary_851_inst_req_1 : boolean;
  signal binary_851_inst_ack_1 : boolean;
  signal ptr_deref_854_base_resize_req_0 : boolean;
  signal ptr_deref_854_base_resize_ack_0 : boolean;
  signal ptr_deref_854_root_address_inst_req_0 : boolean;
  signal ptr_deref_854_root_address_inst_ack_0 : boolean;
  signal ptr_deref_854_addr_0_req_0 : boolean;
  signal ptr_deref_854_addr_0_ack_0 : boolean;
  signal ptr_deref_854_gather_scatter_req_0 : boolean;
  signal ptr_deref_854_gather_scatter_ack_0 : boolean;
  signal ptr_deref_854_store_0_req_0 : boolean;
  signal ptr_deref_854_store_0_ack_0 : boolean;
  signal ptr_deref_854_store_0_req_1 : boolean;
  signal ptr_deref_854_store_0_ack_1 : boolean;
  signal ptr_deref_859_base_resize_req_0 : boolean;
  signal ptr_deref_859_base_resize_ack_0 : boolean;
  signal ptr_deref_859_root_address_inst_req_0 : boolean;
  signal ptr_deref_859_root_address_inst_ack_0 : boolean;
  signal ptr_deref_859_addr_0_req_0 : boolean;
  signal ptr_deref_859_addr_0_ack_0 : boolean;
  signal ptr_deref_859_load_0_req_0 : boolean;
  signal ptr_deref_859_load_0_ack_0 : boolean;
  signal ptr_deref_859_load_0_req_1 : boolean;
  signal ptr_deref_859_load_0_ack_1 : boolean;
  signal ptr_deref_859_gather_scatter_req_0 : boolean;
  signal ptr_deref_859_gather_scatter_ack_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal array_obj_ref_867_index_0_resize_req_0 : boolean;
  signal array_obj_ref_867_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_867_index_0_rename_req_0 : boolean;
  signal array_obj_ref_867_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_867_offset_inst_req_0 : boolean;
  signal array_obj_ref_867_offset_inst_ack_0 : boolean;
  signal array_obj_ref_867_root_address_inst_req_0 : boolean;
  signal array_obj_ref_867_root_address_inst_ack_0 : boolean;
  signal addr_of_868_final_reg_req_0 : boolean;
  signal addr_of_868_final_reg_ack_0 : boolean;
  signal ptr_deref_872_base_resize_req_0 : boolean;
  signal ptr_deref_872_base_resize_ack_0 : boolean;
  signal ptr_deref_872_root_address_inst_req_0 : boolean;
  signal ptr_deref_872_root_address_inst_ack_0 : boolean;
  signal ptr_deref_872_addr_0_req_0 : boolean;
  signal ptr_deref_872_addr_0_ack_0 : boolean;
  signal ptr_deref_872_load_0_req_0 : boolean;
  signal ptr_deref_872_load_0_ack_0 : boolean;
  signal ptr_deref_872_load_0_req_1 : boolean;
  signal ptr_deref_872_load_0_ack_1 : boolean;
  signal ptr_deref_872_gather_scatter_req_0 : boolean;
  signal ptr_deref_872_gather_scatter_ack_0 : boolean;
  signal ptr_deref_876_base_resize_req_0 : boolean;
  signal ptr_deref_876_base_resize_ack_0 : boolean;
  signal ptr_deref_876_root_address_inst_req_0 : boolean;
  signal ptr_deref_876_root_address_inst_ack_0 : boolean;
  signal ptr_deref_876_addr_0_req_0 : boolean;
  signal ptr_deref_876_addr_0_ack_0 : boolean;
  signal ptr_deref_876_load_0_req_0 : boolean;
  signal ptr_deref_876_load_0_ack_0 : boolean;
  signal ptr_deref_876_load_0_req_1 : boolean;
  signal ptr_deref_876_load_0_ack_1 : boolean;
  signal ptr_deref_876_gather_scatter_req_0 : boolean;
  signal ptr_deref_876_gather_scatter_ack_0 : boolean;
  signal type_cast_880_inst_req_0 : boolean;
  signal type_cast_880_inst_ack_0 : boolean;
  signal array_obj_ref_884_index_0_resize_req_0 : boolean;
  signal array_obj_ref_884_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_884_index_0_rename_req_0 : boolean;
  signal array_obj_ref_884_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_884_offset_inst_req_0 : boolean;
  signal array_obj_ref_884_offset_inst_ack_0 : boolean;
  signal array_obj_ref_884_root_address_inst_req_0 : boolean;
  signal array_obj_ref_884_root_address_inst_ack_0 : boolean;
  signal addr_of_885_final_reg_req_0 : boolean;
  signal addr_of_885_final_reg_ack_0 : boolean;
  signal binary_894_inst_req_0 : boolean;
  signal binary_894_inst_ack_0 : boolean;
  signal binary_894_inst_req_1 : boolean;
  signal binary_894_inst_ack_1 : boolean;
  signal ptr_deref_897_base_resize_req_0 : boolean;
  signal ptr_deref_897_base_resize_ack_0 : boolean;
  signal ptr_deref_897_root_address_inst_req_0 : boolean;
  signal ptr_deref_897_root_address_inst_ack_0 : boolean;
  signal ptr_deref_897_addr_0_req_0 : boolean;
  signal ptr_deref_897_addr_0_ack_0 : boolean;
  signal ptr_deref_897_gather_scatter_req_0 : boolean;
  signal ptr_deref_897_gather_scatter_ack_0 : boolean;
  signal ptr_deref_897_store_0_req_0 : boolean;
  signal ptr_deref_897_store_0_ack_0 : boolean;
  signal ptr_deref_1034_load_0_req_0 : boolean;
  signal ptr_deref_897_store_0_req_1 : boolean;
  signal ptr_deref_897_store_0_ack_1 : boolean;
  signal array_obj_ref_1042_offset_inst_req_0 : boolean;
  signal ptr_deref_1046_base_resize_req_0 : boolean;
  signal ptr_deref_1051_root_address_inst_ack_0 : boolean;
  signal ptr_deref_902_base_resize_req_0 : boolean;
  signal ptr_deref_902_base_resize_ack_0 : boolean;
  signal ptr_deref_902_root_address_inst_req_0 : boolean;
  signal ptr_deref_902_root_address_inst_ack_0 : boolean;
  signal ptr_deref_902_addr_0_req_0 : boolean;
  signal ptr_deref_902_addr_0_ack_0 : boolean;
  signal ptr_deref_1046_store_0_ack_0 : boolean;
  signal ptr_deref_1034_load_0_ack_0 : boolean;
  signal ptr_deref_902_load_0_req_0 : boolean;
  signal ptr_deref_902_load_0_ack_0 : boolean;
  signal ptr_deref_902_load_0_req_1 : boolean;
  signal ptr_deref_902_load_0_ack_1 : boolean;
  signal ptr_deref_902_gather_scatter_req_0 : boolean;
  signal ptr_deref_902_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1046_store_0_req_0 : boolean;
  signal ptr_deref_1030_load_0_req_1 : boolean;
  signal ptr_deref_1051_base_resize_ack_0 : boolean;
  signal type_cast_906_inst_req_0 : boolean;
  signal type_cast_906_inst_ack_0 : boolean;
  signal array_obj_ref_1042_offset_inst_ack_0 : boolean;
  signal ptr_deref_1030_load_0_ack_1 : boolean;
  signal ptr_deref_1030_gather_scatter_req_0 : boolean;
  signal ptr_deref_1030_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_910_index_0_resize_req_0 : boolean;
  signal array_obj_ref_910_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_910_index_0_rename_req_0 : boolean;
  signal array_obj_ref_910_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1046_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1042_index_0_rename_req_0 : boolean;
  signal array_obj_ref_910_offset_inst_req_0 : boolean;
  signal array_obj_ref_910_offset_inst_ack_0 : boolean;
  signal array_obj_ref_910_root_address_inst_req_0 : boolean;
  signal array_obj_ref_910_root_address_inst_ack_0 : boolean;
  signal addr_of_911_final_reg_req_0 : boolean;
  signal addr_of_911_final_reg_ack_0 : boolean;
  signal ptr_deref_1034_root_address_inst_req_0 : boolean;
  signal ptr_deref_1034_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1046_root_address_inst_req_0 : boolean;
  signal ptr_deref_915_base_resize_req_0 : boolean;
  signal ptr_deref_915_base_resize_ack_0 : boolean;
  signal array_obj_ref_1042_index_0_rename_ack_0 : boolean;
  signal ptr_deref_915_root_address_inst_req_0 : boolean;
  signal ptr_deref_915_root_address_inst_ack_0 : boolean;
  signal ptr_deref_915_addr_0_req_0 : boolean;
  signal ptr_deref_915_addr_0_ack_0 : boolean;
  signal ptr_deref_915_load_0_req_0 : boolean;
  signal ptr_deref_915_load_0_ack_0 : boolean;
  signal ptr_deref_915_load_0_req_1 : boolean;
  signal ptr_deref_915_load_0_ack_1 : boolean;
  signal ptr_deref_915_gather_scatter_req_0 : boolean;
  signal ptr_deref_915_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1051_root_address_inst_req_0 : boolean;
  signal ptr_deref_1034_load_0_req_1 : boolean;
  signal ptr_deref_919_base_resize_req_0 : boolean;
  signal ptr_deref_919_base_resize_ack_0 : boolean;
  signal ptr_deref_919_root_address_inst_req_0 : boolean;
  signal ptr_deref_919_root_address_inst_ack_0 : boolean;
  signal ptr_deref_919_addr_0_req_0 : boolean;
  signal ptr_deref_919_addr_0_ack_0 : boolean;
  signal ptr_deref_1034_load_0_ack_1 : boolean;
  signal ptr_deref_919_load_0_req_0 : boolean;
  signal ptr_deref_919_load_0_ack_0 : boolean;
  signal type_cast_1038_inst_req_0 : boolean;
  signal ptr_deref_919_load_0_req_1 : boolean;
  signal ptr_deref_919_load_0_ack_1 : boolean;
  signal ptr_deref_919_gather_scatter_req_0 : boolean;
  signal ptr_deref_919_gather_scatter_ack_0 : boolean;
  signal type_cast_923_inst_req_0 : boolean;
  signal type_cast_923_inst_ack_0 : boolean;
  signal array_obj_ref_927_index_0_resize_req_0 : boolean;
  signal array_obj_ref_927_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_927_index_0_rename_req_0 : boolean;
  signal array_obj_ref_927_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_927_offset_inst_req_0 : boolean;
  signal array_obj_ref_927_offset_inst_ack_0 : boolean;
  signal array_obj_ref_927_root_address_inst_req_0 : boolean;
  signal array_obj_ref_927_root_address_inst_ack_0 : boolean;
  signal addr_of_928_final_reg_req_0 : boolean;
  signal addr_of_928_final_reg_ack_0 : boolean;
  signal ptr_deref_932_base_resize_req_0 : boolean;
  signal ptr_deref_932_base_resize_ack_0 : boolean;
  signal ptr_deref_932_root_address_inst_req_0 : boolean;
  signal ptr_deref_932_root_address_inst_ack_0 : boolean;
  signal ptr_deref_932_addr_0_req_0 : boolean;
  signal ptr_deref_932_addr_0_ack_0 : boolean;
  signal ptr_deref_932_load_0_req_0 : boolean;
  signal ptr_deref_932_load_0_ack_0 : boolean;
  signal ptr_deref_932_load_0_req_1 : boolean;
  signal ptr_deref_932_load_0_ack_1 : boolean;
  signal ptr_deref_932_gather_scatter_req_0 : boolean;
  signal ptr_deref_932_gather_scatter_ack_0 : boolean;
  signal binary_937_inst_req_0 : boolean;
  signal binary_937_inst_ack_0 : boolean;
  signal binary_937_inst_req_1 : boolean;
  signal binary_937_inst_ack_1 : boolean;
  signal ptr_deref_940_base_resize_req_0 : boolean;
  signal ptr_deref_940_base_resize_ack_0 : boolean;
  signal ptr_deref_940_root_address_inst_req_0 : boolean;
  signal ptr_deref_940_root_address_inst_ack_0 : boolean;
  signal ptr_deref_940_addr_0_req_0 : boolean;
  signal ptr_deref_940_addr_0_ack_0 : boolean;
  signal ptr_deref_940_gather_scatter_req_0 : boolean;
  signal ptr_deref_940_gather_scatter_ack_0 : boolean;
  signal ptr_deref_940_store_0_req_0 : boolean;
  signal ptr_deref_940_store_0_ack_0 : boolean;
  signal ptr_deref_940_store_0_req_1 : boolean;
  signal ptr_deref_940_store_0_ack_1 : boolean;
  signal ptr_deref_945_base_resize_req_0 : boolean;
  signal ptr_deref_945_base_resize_ack_0 : boolean;
  signal ptr_deref_945_root_address_inst_req_0 : boolean;
  signal ptr_deref_945_root_address_inst_ack_0 : boolean;
  signal ptr_deref_945_addr_0_req_0 : boolean;
  signal ptr_deref_945_addr_0_ack_0 : boolean;
  signal ptr_deref_945_load_0_req_0 : boolean;
  signal ptr_deref_945_load_0_ack_0 : boolean;
  signal ptr_deref_945_load_0_req_1 : boolean;
  signal ptr_deref_945_load_0_ack_1 : boolean;
  signal ptr_deref_945_gather_scatter_req_0 : boolean;
  signal ptr_deref_945_gather_scatter_ack_0 : boolean;
  signal type_cast_949_inst_req_0 : boolean;
  signal type_cast_949_inst_ack_0 : boolean;
  signal array_obj_ref_953_index_0_resize_req_0 : boolean;
  signal array_obj_ref_953_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_953_index_0_rename_req_0 : boolean;
  signal array_obj_ref_953_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_953_offset_inst_req_0 : boolean;
  signal array_obj_ref_953_offset_inst_ack_0 : boolean;
  signal array_obj_ref_953_root_address_inst_req_0 : boolean;
  signal array_obj_ref_953_root_address_inst_ack_0 : boolean;
  signal addr_of_954_final_reg_req_0 : boolean;
  signal addr_of_954_final_reg_ack_0 : boolean;
  signal ptr_deref_958_base_resize_req_0 : boolean;
  signal ptr_deref_958_base_resize_ack_0 : boolean;
  signal ptr_deref_958_root_address_inst_req_0 : boolean;
  signal ptr_deref_958_root_address_inst_ack_0 : boolean;
  signal ptr_deref_958_addr_0_req_0 : boolean;
  signal ptr_deref_958_addr_0_ack_0 : boolean;
  signal ptr_deref_958_load_0_req_0 : boolean;
  signal ptr_deref_958_load_0_ack_0 : boolean;
  signal ptr_deref_958_load_0_req_1 : boolean;
  signal ptr_deref_958_load_0_ack_1 : boolean;
  signal ptr_deref_958_gather_scatter_req_0 : boolean;
  signal ptr_deref_958_gather_scatter_ack_0 : boolean;
  signal ptr_deref_962_base_resize_req_0 : boolean;
  signal ptr_deref_962_base_resize_ack_0 : boolean;
  signal ptr_deref_962_root_address_inst_req_0 : boolean;
  signal ptr_deref_962_root_address_inst_ack_0 : boolean;
  signal ptr_deref_962_addr_0_req_0 : boolean;
  signal ptr_deref_962_addr_0_ack_0 : boolean;
  signal ptr_deref_962_load_0_req_0 : boolean;
  signal ptr_deref_962_load_0_ack_0 : boolean;
  signal ptr_deref_962_load_0_req_1 : boolean;
  signal ptr_deref_962_load_0_ack_1 : boolean;
  signal ptr_deref_962_gather_scatter_req_0 : boolean;
  signal ptr_deref_962_gather_scatter_ack_0 : boolean;
  signal type_cast_966_inst_req_0 : boolean;
  signal type_cast_966_inst_ack_0 : boolean;
  signal array_obj_ref_970_index_0_resize_req_0 : boolean;
  signal array_obj_ref_970_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_970_index_0_rename_req_0 : boolean;
  signal array_obj_ref_970_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_970_offset_inst_req_0 : boolean;
  signal array_obj_ref_970_offset_inst_ack_0 : boolean;
  signal array_obj_ref_970_root_address_inst_req_0 : boolean;
  signal array_obj_ref_970_root_address_inst_ack_0 : boolean;
  signal addr_of_971_final_reg_req_0 : boolean;
  signal addr_of_971_final_reg_ack_0 : boolean;
  signal ptr_deref_975_base_resize_req_0 : boolean;
  signal ptr_deref_975_base_resize_ack_0 : boolean;
  signal ptr_deref_975_root_address_inst_req_0 : boolean;
  signal ptr_deref_975_root_address_inst_ack_0 : boolean;
  signal ptr_deref_975_addr_0_req_0 : boolean;
  signal ptr_deref_975_addr_0_ack_0 : boolean;
  signal ptr_deref_975_load_0_req_0 : boolean;
  signal ptr_deref_975_load_0_ack_0 : boolean;
  signal ptr_deref_975_load_0_req_1 : boolean;
  signal ptr_deref_975_load_0_ack_1 : boolean;
  signal ptr_deref_975_gather_scatter_req_0 : boolean;
  signal ptr_deref_975_gather_scatter_ack_0 : boolean;
  signal binary_980_inst_req_0 : boolean;
  signal binary_980_inst_ack_0 : boolean;
  signal binary_980_inst_req_1 : boolean;
  signal binary_980_inst_ack_1 : boolean;
  signal ptr_deref_983_base_resize_req_0 : boolean;
  signal ptr_deref_983_base_resize_ack_0 : boolean;
  signal ptr_deref_983_root_address_inst_req_0 : boolean;
  signal ptr_deref_983_root_address_inst_ack_0 : boolean;
  signal ptr_deref_983_addr_0_req_0 : boolean;
  signal ptr_deref_983_addr_0_ack_0 : boolean;
  signal ptr_deref_983_gather_scatter_req_0 : boolean;
  signal ptr_deref_983_gather_scatter_ack_0 : boolean;
  signal ptr_deref_983_store_0_req_0 : boolean;
  signal ptr_deref_983_store_0_ack_0 : boolean;
  signal ptr_deref_983_store_0_req_1 : boolean;
  signal ptr_deref_983_store_0_ack_1 : boolean;
  signal ptr_deref_988_base_resize_req_0 : boolean;
  signal ptr_deref_988_base_resize_ack_0 : boolean;
  signal ptr_deref_988_root_address_inst_req_0 : boolean;
  signal ptr_deref_988_root_address_inst_ack_0 : boolean;
  signal ptr_deref_988_addr_0_req_0 : boolean;
  signal ptr_deref_988_addr_0_ack_0 : boolean;
  signal ptr_deref_988_load_0_req_0 : boolean;
  signal ptr_deref_988_load_0_ack_0 : boolean;
  signal ptr_deref_992_root_address_inst_req_0 : boolean;
  signal ptr_deref_992_root_address_inst_ack_0 : boolean;
  signal ptr_deref_992_addr_0_req_0 : boolean;
  signal ptr_deref_992_addr_0_ack_0 : boolean;
  signal ptr_deref_992_load_0_req_0 : boolean;
  signal ptr_deref_992_load_0_ack_0 : boolean;
  signal ptr_deref_992_load_0_req_1 : boolean;
  signal ptr_deref_992_load_0_ack_1 : boolean;
  signal ptr_deref_992_gather_scatter_req_0 : boolean;
  signal ptr_deref_992_gather_scatter_ack_0 : boolean;
  signal type_cast_996_inst_req_0 : boolean;
  signal type_cast_996_inst_ack_0 : boolean;
  signal array_obj_ref_1000_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1000_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1000_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1000_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1051_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1000_offset_inst_req_0 : boolean;
  signal array_obj_ref_1000_offset_inst_ack_0 : boolean;
  signal ptr_deref_1051_load_0_req_1 : boolean;
  signal array_obj_ref_1000_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1000_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1051_load_0_ack_1 : boolean;
  signal ptr_deref_1051_addr_0_ack_0 : boolean;
  signal addr_of_1001_final_reg_req_0 : boolean;
  signal addr_of_1001_final_reg_ack_0 : boolean;
  signal ptr_deref_1030_load_0_req_0 : boolean;
  signal ptr_deref_1051_base_resize_req_0 : boolean;
  signal ptr_deref_1046_base_resize_ack_0 : boolean;
  signal ptr_deref_1046_addr_0_ack_0 : boolean;
  signal ptr_deref_1004_base_resize_req_0 : boolean;
  signal ptr_deref_1004_base_resize_ack_0 : boolean;
  signal ptr_deref_1046_store_0_ack_1 : boolean;
  signal ptr_deref_1004_root_address_inst_req_0 : boolean;
  signal ptr_deref_1004_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1046_store_0_req_1 : boolean;
  signal ptr_deref_1030_addr_0_ack_0 : boolean;
  signal ptr_deref_1004_addr_0_req_0 : boolean;
  signal ptr_deref_1004_addr_0_ack_0 : boolean;
  signal ptr_deref_1030_addr_0_req_0 : boolean;
  signal ptr_deref_1004_gather_scatter_req_0 : boolean;
  signal ptr_deref_1004_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1004_store_0_req_0 : boolean;
  signal ptr_deref_1004_store_0_ack_0 : boolean;
  signal ptr_deref_1046_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1004_store_0_req_1 : boolean;
  signal ptr_deref_1004_store_0_ack_1 : boolean;
  signal ptr_deref_1051_load_0_ack_0 : boolean;
  signal ptr_deref_1051_load_0_req_0 : boolean;
  signal ptr_deref_1051_addr_0_req_0 : boolean;
  signal array_obj_ref_1042_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1030_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1030_root_address_inst_req_0 : boolean;
  signal ptr_deref_1046_addr_0_req_0 : boolean;
  signal ptr_deref_1046_gather_scatter_req_0 : boolean;
  signal ptr_deref_1030_base_resize_ack_0 : boolean;
  signal addr_of_1043_final_reg_ack_0 : boolean;
  signal ptr_deref_1009_base_resize_req_0 : boolean;
  signal ptr_deref_1009_base_resize_ack_0 : boolean;
  signal ptr_deref_1030_base_resize_req_0 : boolean;
  signal array_obj_ref_1042_index_0_resize_req_0 : boolean;
  signal addr_of_1043_final_reg_req_0 : boolean;
  signal ptr_deref_1009_root_address_inst_req_0 : boolean;
  signal ptr_deref_1009_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1009_addr_0_req_0 : boolean;
  signal ptr_deref_1009_addr_0_ack_0 : boolean;
  signal ptr_deref_1009_load_0_req_0 : boolean;
  signal ptr_deref_1009_load_0_ack_0 : boolean;
  signal array_obj_ref_1042_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1042_root_address_inst_req_0 : boolean;
  signal ptr_deref_1009_load_0_req_1 : boolean;
  signal ptr_deref_1009_load_0_ack_1 : boolean;
  signal ptr_deref_1009_gather_scatter_req_0 : boolean;
  signal ptr_deref_1009_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1034_addr_0_ack_0 : boolean;
  signal ptr_deref_1034_addr_0_req_0 : boolean;
  signal ptr_deref_1013_base_resize_req_0 : boolean;
  signal ptr_deref_1013_base_resize_ack_0 : boolean;
  signal ptr_deref_1175_base_resize_ack_0 : boolean;
  signal ptr_deref_1013_root_address_inst_req_0 : boolean;
  signal ptr_deref_1013_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1013_addr_0_req_0 : boolean;
  signal ptr_deref_1013_addr_0_ack_0 : boolean;
  signal ptr_deref_1175_addr_0_req_0 : boolean;
  signal ptr_deref_1013_load_0_req_0 : boolean;
  signal ptr_deref_1013_load_0_ack_0 : boolean;
  signal ptr_deref_1013_load_0_req_1 : boolean;
  signal ptr_deref_1013_load_0_ack_1 : boolean;
  signal ptr_deref_1013_gather_scatter_req_0 : boolean;
  signal ptr_deref_1013_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1175_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1175_root_address_inst_req_0 : boolean;
  signal ptr_deref_1175_root_address_inst_ack_0 : boolean;
  signal type_cast_1017_inst_req_0 : boolean;
  signal type_cast_1017_inst_ack_0 : boolean;
  signal ptr_deref_1175_gather_scatter_req_0 : boolean;
  signal ptr_deref_1175_base_resize_req_0 : boolean;
  signal array_obj_ref_1021_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1021_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1175_store_0_req_0 : boolean;
  signal array_obj_ref_1021_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1021_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1021_offset_inst_req_0 : boolean;
  signal array_obj_ref_1021_offset_inst_ack_0 : boolean;
  signal ptr_deref_1175_addr_0_ack_0 : boolean;
  signal array_obj_ref_1021_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1021_root_address_inst_ack_0 : boolean;
  signal addr_of_1022_final_reg_req_0 : boolean;
  signal addr_of_1022_final_reg_ack_0 : boolean;
  signal ptr_deref_1025_base_resize_req_0 : boolean;
  signal ptr_deref_1025_base_resize_ack_0 : boolean;
  signal ptr_deref_1025_root_address_inst_req_0 : boolean;
  signal ptr_deref_1025_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1025_addr_0_req_0 : boolean;
  signal ptr_deref_1025_addr_0_ack_0 : boolean;
  signal ptr_deref_1025_gather_scatter_req_0 : boolean;
  signal ptr_deref_1025_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1025_store_0_req_0 : boolean;
  signal ptr_deref_1025_store_0_ack_0 : boolean;
  signal ptr_deref_1025_store_0_req_1 : boolean;
  signal ptr_deref_1025_store_0_ack_1 : boolean;
  signal ptr_deref_1055_base_resize_req_0 : boolean;
  signal ptr_deref_1055_base_resize_ack_0 : boolean;
  signal ptr_deref_1055_root_address_inst_req_0 : boolean;
  signal ptr_deref_1055_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1055_addr_0_req_0 : boolean;
  signal ptr_deref_1055_addr_0_ack_0 : boolean;
  signal ptr_deref_1055_load_0_req_0 : boolean;
  signal ptr_deref_1055_load_0_ack_0 : boolean;
  signal ptr_deref_1055_load_0_req_1 : boolean;
  signal ptr_deref_1055_load_0_ack_1 : boolean;
  signal ptr_deref_1055_gather_scatter_req_0 : boolean;
  signal ptr_deref_1055_gather_scatter_ack_0 : boolean;
  signal type_cast_1059_inst_req_0 : boolean;
  signal type_cast_1059_inst_ack_0 : boolean;
  signal array_obj_ref_1063_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1063_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1063_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1063_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1063_offset_inst_req_0 : boolean;
  signal array_obj_ref_1063_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1063_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1063_root_address_inst_ack_0 : boolean;
  signal addr_of_1064_final_reg_req_0 : boolean;
  signal addr_of_1064_final_reg_ack_0 : boolean;
  signal ptr_deref_1067_base_resize_req_0 : boolean;
  signal ptr_deref_1067_base_resize_ack_0 : boolean;
  signal ptr_deref_1067_root_address_inst_req_0 : boolean;
  signal ptr_deref_1067_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1067_addr_0_req_0 : boolean;
  signal ptr_deref_1067_addr_0_ack_0 : boolean;
  signal ptr_deref_1067_gather_scatter_req_0 : boolean;
  signal ptr_deref_1067_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1067_store_0_req_0 : boolean;
  signal ptr_deref_1067_store_0_ack_0 : boolean;
  signal ptr_deref_1067_store_0_req_1 : boolean;
  signal ptr_deref_1067_store_0_ack_1 : boolean;
  signal ptr_deref_1072_base_resize_req_0 : boolean;
  signal ptr_deref_1072_base_resize_ack_0 : boolean;
  signal ptr_deref_1072_root_address_inst_req_0 : boolean;
  signal ptr_deref_1072_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1072_addr_0_req_0 : boolean;
  signal ptr_deref_1072_addr_0_ack_0 : boolean;
  signal ptr_deref_1072_load_0_req_0 : boolean;
  signal ptr_deref_1072_load_0_ack_0 : boolean;
  signal ptr_deref_1072_load_0_req_1 : boolean;
  signal ptr_deref_1072_load_0_ack_1 : boolean;
  signal ptr_deref_1072_gather_scatter_req_0 : boolean;
  signal ptr_deref_1072_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1076_base_resize_req_0 : boolean;
  signal ptr_deref_1076_base_resize_ack_0 : boolean;
  signal ptr_deref_1076_root_address_inst_req_0 : boolean;
  signal ptr_deref_1076_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1076_addr_0_req_0 : boolean;
  signal ptr_deref_1076_addr_0_ack_0 : boolean;
  signal ptr_deref_1076_load_0_req_0 : boolean;
  signal ptr_deref_1076_load_0_ack_0 : boolean;
  signal ptr_deref_1076_load_0_req_1 : boolean;
  signal ptr_deref_1076_load_0_ack_1 : boolean;
  signal ptr_deref_1076_gather_scatter_req_0 : boolean;
  signal ptr_deref_1076_gather_scatter_ack_0 : boolean;
  signal type_cast_1080_inst_req_0 : boolean;
  signal type_cast_1080_inst_ack_0 : boolean;
  signal array_obj_ref_1084_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1084_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1084_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1084_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1084_offset_inst_req_0 : boolean;
  signal array_obj_ref_1084_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1084_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1084_root_address_inst_ack_0 : boolean;
  signal addr_of_1085_final_reg_req_0 : boolean;
  signal addr_of_1085_final_reg_ack_0 : boolean;
  signal ptr_deref_1088_base_resize_req_0 : boolean;
  signal ptr_deref_1088_base_resize_ack_0 : boolean;
  signal ptr_deref_1088_root_address_inst_req_0 : boolean;
  signal ptr_deref_1088_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1088_addr_0_req_0 : boolean;
  signal ptr_deref_1088_addr_0_ack_0 : boolean;
  signal ptr_deref_1088_gather_scatter_req_0 : boolean;
  signal ptr_deref_1088_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1088_store_0_req_0 : boolean;
  signal ptr_deref_1088_store_0_ack_0 : boolean;
  signal ptr_deref_1088_store_0_req_1 : boolean;
  signal ptr_deref_1088_store_0_ack_1 : boolean;
  signal ptr_deref_1093_base_resize_req_0 : boolean;
  signal ptr_deref_1093_base_resize_ack_0 : boolean;
  signal ptr_deref_1093_root_address_inst_req_0 : boolean;
  signal ptr_deref_1093_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1093_addr_0_req_0 : boolean;
  signal ptr_deref_1093_addr_0_ack_0 : boolean;
  signal ptr_deref_1093_load_0_req_0 : boolean;
  signal ptr_deref_1093_load_0_ack_0 : boolean;
  signal ptr_deref_1093_load_0_req_1 : boolean;
  signal ptr_deref_1093_load_0_ack_1 : boolean;
  signal ptr_deref_1093_gather_scatter_req_0 : boolean;
  signal ptr_deref_1093_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1097_base_resize_req_0 : boolean;
  signal ptr_deref_1097_base_resize_ack_0 : boolean;
  signal ptr_deref_1097_root_address_inst_req_0 : boolean;
  signal ptr_deref_1097_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1097_addr_0_req_0 : boolean;
  signal ptr_deref_1097_addr_0_ack_0 : boolean;
  signal ptr_deref_1097_load_0_req_0 : boolean;
  signal ptr_deref_1097_load_0_ack_0 : boolean;
  signal ptr_deref_1097_load_0_req_1 : boolean;
  signal ptr_deref_1097_load_0_ack_1 : boolean;
  signal ptr_deref_1097_gather_scatter_req_0 : boolean;
  signal ptr_deref_1097_gather_scatter_ack_0 : boolean;
  signal type_cast_1101_inst_req_0 : boolean;
  signal type_cast_1101_inst_ack_0 : boolean;
  signal array_obj_ref_1105_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1105_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1105_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1105_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1105_offset_inst_req_0 : boolean;
  signal array_obj_ref_1105_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1105_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1105_root_address_inst_ack_0 : boolean;
  signal addr_of_1106_final_reg_req_0 : boolean;
  signal addr_of_1106_final_reg_ack_0 : boolean;
  signal ptr_deref_1109_base_resize_req_0 : boolean;
  signal ptr_deref_1109_base_resize_ack_0 : boolean;
  signal ptr_deref_1109_root_address_inst_req_0 : boolean;
  signal ptr_deref_1109_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1109_addr_0_req_0 : boolean;
  signal ptr_deref_1109_addr_0_ack_0 : boolean;
  signal ptr_deref_1109_gather_scatter_req_0 : boolean;
  signal ptr_deref_1109_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1109_store_0_req_0 : boolean;
  signal ptr_deref_1109_store_0_ack_0 : boolean;
  signal ptr_deref_1109_store_0_req_1 : boolean;
  signal ptr_deref_1109_store_0_ack_1 : boolean;
  signal ptr_deref_1114_base_resize_req_0 : boolean;
  signal ptr_deref_1114_base_resize_ack_0 : boolean;
  signal ptr_deref_1114_root_address_inst_req_0 : boolean;
  signal ptr_deref_1114_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1114_addr_0_req_0 : boolean;
  signal ptr_deref_1114_addr_0_ack_0 : boolean;
  signal ptr_deref_1114_load_0_req_0 : boolean;
  signal ptr_deref_1114_load_0_ack_0 : boolean;
  signal ptr_deref_1114_load_0_req_1 : boolean;
  signal ptr_deref_1114_load_0_ack_1 : boolean;
  signal ptr_deref_1114_gather_scatter_req_0 : boolean;
  signal ptr_deref_1114_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1118_base_resize_req_0 : boolean;
  signal ptr_deref_1118_base_resize_ack_0 : boolean;
  signal ptr_deref_1118_root_address_inst_req_0 : boolean;
  signal ptr_deref_1118_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1118_addr_0_req_0 : boolean;
  signal ptr_deref_1118_addr_0_ack_0 : boolean;
  signal ptr_deref_1118_load_0_req_0 : boolean;
  signal ptr_deref_1118_load_0_ack_0 : boolean;
  signal ptr_deref_1118_load_0_req_1 : boolean;
  signal ptr_deref_1118_load_0_ack_1 : boolean;
  signal ptr_deref_1118_gather_scatter_req_0 : boolean;
  signal ptr_deref_1118_gather_scatter_ack_0 : boolean;
  signal type_cast_1122_inst_req_0 : boolean;
  signal type_cast_1122_inst_ack_0 : boolean;
  signal array_obj_ref_1126_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1126_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1126_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1126_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1126_offset_inst_req_0 : boolean;
  signal array_obj_ref_1126_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1126_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1126_root_address_inst_ack_0 : boolean;
  signal addr_of_1127_final_reg_req_0 : boolean;
  signal addr_of_1127_final_reg_ack_0 : boolean;
  signal ptr_deref_1130_base_resize_req_0 : boolean;
  signal ptr_deref_1130_base_resize_ack_0 : boolean;
  signal ptr_deref_1130_root_address_inst_req_0 : boolean;
  signal ptr_deref_1130_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1130_addr_0_req_0 : boolean;
  signal ptr_deref_1130_addr_0_ack_0 : boolean;
  signal ptr_deref_1130_gather_scatter_req_0 : boolean;
  signal ptr_deref_1130_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1130_store_0_req_0 : boolean;
  signal ptr_deref_1130_store_0_ack_0 : boolean;
  signal ptr_deref_1130_store_0_req_1 : boolean;
  signal ptr_deref_1130_store_0_ack_1 : boolean;
  signal ptr_deref_1135_base_resize_req_0 : boolean;
  signal ptr_deref_1135_base_resize_ack_0 : boolean;
  signal ptr_deref_1135_root_address_inst_req_0 : boolean;
  signal ptr_deref_1135_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1135_addr_0_req_0 : boolean;
  signal ptr_deref_1135_addr_0_ack_0 : boolean;
  signal ptr_deref_1135_load_0_req_0 : boolean;
  signal ptr_deref_1135_load_0_ack_0 : boolean;
  signal ptr_deref_1135_load_0_req_1 : boolean;
  signal ptr_deref_1135_load_0_ack_1 : boolean;
  signal ptr_deref_1135_gather_scatter_req_0 : boolean;
  signal ptr_deref_1135_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1139_base_resize_req_0 : boolean;
  signal ptr_deref_1139_base_resize_ack_0 : boolean;
  signal ptr_deref_1139_root_address_inst_req_0 : boolean;
  signal ptr_deref_1139_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1139_addr_0_req_0 : boolean;
  signal ptr_deref_1139_addr_0_ack_0 : boolean;
  signal ptr_deref_1139_load_0_req_0 : boolean;
  signal ptr_deref_1139_load_0_ack_0 : boolean;
  signal ptr_deref_1139_load_0_req_1 : boolean;
  signal ptr_deref_1139_load_0_ack_1 : boolean;
  signal ptr_deref_1139_gather_scatter_req_0 : boolean;
  signal ptr_deref_1139_gather_scatter_ack_0 : boolean;
  signal type_cast_1143_inst_req_0 : boolean;
  signal type_cast_1143_inst_ack_0 : boolean;
  signal array_obj_ref_1147_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1147_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1147_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1147_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1147_offset_inst_req_0 : boolean;
  signal array_obj_ref_1147_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1147_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1147_root_address_inst_ack_0 : boolean;
  signal addr_of_1148_final_reg_req_0 : boolean;
  signal addr_of_1148_final_reg_ack_0 : boolean;
  signal ptr_deref_1151_base_resize_req_0 : boolean;
  signal ptr_deref_1151_base_resize_ack_0 : boolean;
  signal ptr_deref_1151_root_address_inst_req_0 : boolean;
  signal ptr_deref_1151_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1151_addr_0_req_0 : boolean;
  signal ptr_deref_1151_addr_0_ack_0 : boolean;
  signal ptr_deref_1151_gather_scatter_req_0 : boolean;
  signal ptr_deref_1151_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1151_store_0_req_0 : boolean;
  signal ptr_deref_1151_store_0_ack_0 : boolean;
  signal ptr_deref_1151_store_0_req_1 : boolean;
  signal ptr_deref_1151_store_0_ack_1 : boolean;
  signal ptr_deref_1158_base_resize_req_0 : boolean;
  signal ptr_deref_1158_base_resize_ack_0 : boolean;
  signal ptr_deref_1158_root_address_inst_req_0 : boolean;
  signal ptr_deref_1158_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1158_addr_0_req_0 : boolean;
  signal ptr_deref_1158_addr_0_ack_0 : boolean;
  signal ptr_deref_1158_load_0_req_0 : boolean;
  signal ptr_deref_1158_load_0_ack_0 : boolean;
  signal ptr_deref_1158_load_0_req_1 : boolean;
  signal ptr_deref_1158_load_0_ack_1 : boolean;
  signal ptr_deref_1158_gather_scatter_req_0 : boolean;
  signal ptr_deref_1158_gather_scatter_ack_0 : boolean;
  signal type_cast_1162_inst_req_0 : boolean;
  signal type_cast_1162_inst_ack_0 : boolean;
  signal ptr_deref_1175_store_0_ack_0 : boolean;
  signal binary_1168_inst_req_0 : boolean;
  signal binary_1168_inst_ack_0 : boolean;
  signal binary_1168_inst_req_1 : boolean;
  signal binary_1168_inst_ack_1 : boolean;
  signal type_cast_1172_inst_req_0 : boolean;
  signal type_cast_1172_inst_ack_0 : boolean;
  signal ptr_deref_1175_store_0_req_1 : boolean;
  signal ptr_deref_1175_store_0_ack_1 : boolean;
  signal memory_space_10_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_10_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_10_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_10_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_10_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_10_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_10_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_10_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_10_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_10_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_11_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_11_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_11_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_11_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_11_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_11_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_11_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_11_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_11_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_11_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_12_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_12_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_12_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_12_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_12_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_12_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_12_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_12_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_12_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_12_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_13_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_13_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_13_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_13_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_13_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_13_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_13_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_13_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_13_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_13_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_14_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_14_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_14_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_14_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_14_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_14_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_14_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_14_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_14_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_14_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_14_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_15_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_15_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_15_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_15_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_15_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_15_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_15_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_15_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_15_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_15_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_15_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_16_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_16_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_16_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_16_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_16_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_16_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_16_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_16_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_16_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_17_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_17_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_17_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_17_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_17_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_17_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_17_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_17_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_17_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_18_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_18_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_18_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_18_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_18_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_18_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_18_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_18_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_18_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_18_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_18_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_18_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_18_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_18_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_18_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_18_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_19_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_19_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_19_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_19_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_19_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_19_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_19_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_19_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_19_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_19_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_19_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_19_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_19_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_19_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_19_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_19_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_20_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_20_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_20_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_20_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_20_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_20_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_20_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_20_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_20_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_20_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_20_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_20_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_20_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_20_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_20_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_20_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_21_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_21_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_21_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_21_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_21_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_21_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_21_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_21_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_21_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_21_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_21_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_21_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_21_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_21_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_21_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_21_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_22_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_22_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_22_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_22_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_22_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_22_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_22_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_22_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_22_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_22_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_22_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_22_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_22_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_22_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_22_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_22_sc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(1 downto 0);
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"x_vectorSum_x start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"x_vectorSum_x start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"x_vectorSum_x fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"x_vectorSum_x fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  x_vectorSum_x_xCP_2164: Block -- control-path 
    signal cp_elements: BooleanArray(971 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(40);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(40), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  bypass 
    -- predecessors 
    -- successors 5 
    -- members (4) 
      -- 	$entry
      -- 	branch_block_stmt_377/$entry
      -- 	branch_block_stmt_377/branch_block_stmt_377__entry__
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462__entry__
      -- 
    -- CP-element group 1 branch  place  bypass 
    -- predecessors 31 
    -- successors 32 35 
    -- members (2) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480__exit__
      -- 	branch_block_stmt_377/if_stmt_481__entry__
      -- 
    cp_elements(1) <= cp_elements(31);
    -- CP-element group 2 merge  place  bypass 
    -- predecessors 38 971 
    -- successors 41 
    -- members (2) 
      -- 	branch_block_stmt_377/merge_stmt_487__exit__
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153__entry__
      -- 
    cp_elements(2) <= OrReduce(cp_elements(38) & cp_elements(971));
    -- CP-element group 3 transition  place  bypass 
    -- predecessors 942 
    -- successors 943 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153__exit__
      -- 	branch_block_stmt_377/bb_2_bb_3
      -- 	branch_block_stmt_377/merge_stmt_1155__exit__
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177__entry__
      -- 	branch_block_stmt_377/merge_stmt_1155_PhiReqMerge
      -- 	branch_block_stmt_377/bb_2_bb_3_PhiReq/$entry
      -- 	branch_block_stmt_377/bb_2_bb_3_PhiReq/$exit
      -- 	branch_block_stmt_377/merge_stmt_1155_PhiAck/$entry
      -- 	branch_block_stmt_377/merge_stmt_1155_PhiAck/$exit
      -- 	branch_block_stmt_377/merge_stmt_1155_PhiAck/dummy
      -- 
    cp_elements(3) <= cp_elements(942);
    -- CP-element group 4 transition  place  bypass 
    -- predecessors 967 
    -- successors 968 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177__exit__
      -- 	branch_block_stmt_377/bb_3_bb_1
      -- 	branch_block_stmt_377/bb_3_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_377/bb_3_bb_1_PhiReq/$exit
      -- 
    cp_elements(4) <= cp_elements(967);
    -- CP-element group 5 fork  transition  bypass 
    -- predecessors 0 
    -- successors 6 8 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/$entry
      -- 
    cp_elements(5) <= cp_elements(0);
    -- CP-element group 6 transition  bypass 
    -- predecessors 5 
    -- successors 7 
    -- members (2) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/assign_stmt_462_trigger_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/assign_stmt_462_active_
      -- 
    cp_elements(6) <= cp_elements(5);
    -- CP-element group 7 join  transition  output  no-bypass 
    -- predecessors 6 11 
    -- successors 12 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_trigger_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/split_req
      -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(6);
      predecessors(1) <= cp_elements(11);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(7)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_459_gather_scatter_req_0); -- 
    -- CP-element group 8 transition  output  bypass 
    -- predecessors 5 
    -- successors 9 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/simple_obj_ref_458_trigger_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/simple_obj_ref_458_active_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/simple_obj_ref_458_completed_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_addr_resize/base_resize_req
      -- 
    cp_elements(8) <= cp_elements(5);
    base_resize_req_2211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => ptr_deref_459_base_resize_req_0); -- 
    -- CP-element group 9 transition  input  output  no-bypass 
    -- predecessors 8 
    -- successors 10 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_base_resize_ack_0, ack => cp_elements(9)); -- 
    sum_rename_req_2216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => ptr_deref_459_root_address_inst_req_0); -- 
    -- CP-element group 10 transition  input  output  no-bypass 
    -- predecessors 9 
    -- successors 11 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2217_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_root_address_inst_ack_0, ack => cp_elements(10)); -- 
    root_register_req_2221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_459_addr_0_req_0); -- 
    -- CP-element group 11 transition  input  no-bypass 
    -- predecessors 10 
    -- successors 7 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_word_addrgen/root_register_ack
      -- 
    root_register_ack_2222_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_addr_0_ack_0, ack => cp_elements(11)); -- 
    -- CP-element group 12 transition  input  output  no-bypass 
    -- predecessors 7 
    -- successors 13 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/word_access_0/rr
      -- 
    split_ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_gather_scatter_ack_0, ack => cp_elements(12)); -- 
    rr_2234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => ptr_deref_459_store_0_req_0); -- 
    -- CP-element group 13 transition  input  output  no-bypass 
    -- predecessors 12 
    -- successors 14 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_active_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/word_access_0/cr
      -- 
    ra_2235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_store_0_ack_0, ack => cp_elements(13)); -- 
    cr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_459_store_0_req_1); -- 
    -- CP-element group 14 transition  place  input  no-bypass 
    -- predecessors 13 
    -- successors 968 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462__exit__
      -- 	branch_block_stmt_377/bb_0_bb_1
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/assign_stmt_462_completed_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_completed_
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_397_to_assign_stmt_462/ptr_deref_459_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/bb_0_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_377/bb_0_bb_1_PhiReq/$exit
      -- 
    ca_2246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_459_store_0_ack_1, ack => cp_elements(14)); -- 
    -- CP-element group 15 fork  transition  bypass 
    -- predecessors 969 
    -- successors 16 24 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/$entry
      -- 
    cp_elements(15) <= cp_elements(969);
    -- CP-element group 16 transition  output  bypass 
    -- predecessors 15 
    -- successors 17 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_466_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_466_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_466_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_addr_resize/base_resize_req
      -- 
    cp_elements(16) <= cp_elements(15);
    base_resize_req_2266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_467_base_resize_req_0); -- 
    -- CP-element group 17 transition  input  output  no-bypass 
    -- predecessors 16 
    -- successors 18 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_base_resize_ack_0, ack => cp_elements(17)); -- 
    sum_rename_req_2271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_467_root_address_inst_req_0); -- 
    -- CP-element group 18 transition  input  output  no-bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_root_address_inst_ack_0, ack => cp_elements(18)); -- 
    root_register_req_2276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_467_addr_0_req_0); -- 
    -- CP-element group 19 transition  input  output  no-bypass 
    -- predecessors 18 
    -- successors 20 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/word_access_0/rr
      -- 
    root_register_ack_2277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_addr_0_ack_0, ack => cp_elements(19)); -- 
    rr_2287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_467_load_0_req_0); -- 
    -- CP-element group 20 transition  input  output  no-bypass 
    -- predecessors 19 
    -- successors 21 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/word_access_0/cr
      -- 
    ra_2288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_0, ack => cp_elements(20)); -- 
    cr_2298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_467_load_0_req_1); -- 
    -- CP-element group 21 transition  input  output  no-bypass 
    -- predecessors 20 
    -- successors 22 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/merge_req
      -- 
    ca_2299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_load_0_ack_1, ack => cp_elements(21)); -- 
    merge_req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_467_gather_scatter_req_0); -- 
    -- CP-element group 22 transition  input  output  no-bypass 
    -- predecessors 21 
    -- successors 23 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_468_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_468_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_468_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/ptr_deref_467_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_470_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_470_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_470_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_complete/req
      -- 
    merge_ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_467_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => type_cast_471_inst_req_0); -- 
    -- CP-element group 23 transition  input  output  no-bypass 
    -- predecessors 22 
    -- successors 28 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_472_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_472_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_472_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_471_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_474_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_474_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/simple_obj_ref_474_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_complete/req
      -- 
    ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_471_inst_ack_0, ack => cp_elements(23)); -- 
    req_2335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => type_cast_475_inst_req_0); -- 
    -- CP-element group 24 transition  bypass 
    -- predecessors 15 
    -- successors 31 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_active_
      -- 
    cp_elements(24) <= cp_elements(15);
    -- CP-element group 25 join  transition  bypass 
    -- predecessors 29 30 
    -- successors 31 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_480_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_480_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/assign_stmt_480_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_completed_
      -- 
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(29);
      predecessors(1) <= cp_elements(30);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(25)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 26 transition  output  bypass 
    -- predecessors 28 
    -- successors 29 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Sample/rr
      -- 
    cp_elements(26) <= cp_elements(28);
    rr_2340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_479_inst_req_0); -- 
    -- CP-element group 27 transition  output  bypass 
    -- predecessors 28 
    -- successors 30 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_update_start_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Update/cr
      -- 
    cp_elements(27) <= cp_elements(28);
    cr_2345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => binary_479_inst_req_1); -- 
    -- CP-element group 28 fork  transition  input  no-bypass 
    -- predecessors 23 
    -- successors 26 27 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_trigger_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_active_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/type_cast_475_complete/ack
      -- 
    ack_2336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_475_inst_ack_0, ack => cp_elements(28)); -- 
    -- CP-element group 29 transition  input  no-bypass 
    -- predecessors 26 
    -- successors 25 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Sample/ra
      -- 
    ra_2341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_479_inst_ack_0, ack => cp_elements(29)); -- 
    -- CP-element group 30 transition  input  no-bypass 
    -- predecessors 27 
    -- successors 25 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/binary_479_Update/ca
      -- 
    ca_2346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_479_inst_ack_1, ack => cp_elements(30)); -- 
    -- CP-element group 31 join  transition  no-bypass 
    -- predecessors 24 25 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480/$exit
      -- 
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(24);
      predecessors(1) <= cp_elements(25);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(31)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 32 transition  bypass 
    -- predecessors 1 
    -- successors 33 
    -- members (1) 
      -- 	branch_block_stmt_377/if_stmt_481_dead_link/$entry
      -- 
    cp_elements(32) <= cp_elements(1);
    -- CP-element group 33 transition  dead  bypass 
    -- predecessors 32 
    -- successors 34 
    -- members (1) 
      -- 	branch_block_stmt_377/if_stmt_481_dead_link/dead_transition
      -- 
    cp_elements(33) <= false;
    -- CP-element group 34 transition  place  bypass 
    -- predecessors 33 
    -- successors 970 
    -- members (4) 
      -- 	branch_block_stmt_377/if_stmt_481__exit__
      -- 	branch_block_stmt_377/merge_stmt_487__entry__
      -- 	branch_block_stmt_377/if_stmt_481_dead_link/$exit
      -- 	branch_block_stmt_377/merge_stmt_487_dead_link/$entry
      -- 
    cp_elements(34) <= cp_elements(33);
    -- CP-element group 35 transition  output  bypass 
    -- predecessors 1 
    -- successors 36 
    -- members (3) 
      -- 	branch_block_stmt_377/if_stmt_481_eval_test/$entry
      -- 	branch_block_stmt_377/if_stmt_481_eval_test/$exit
      -- 	branch_block_stmt_377/if_stmt_481_eval_test/branch_req
      -- 
    cp_elements(35) <= cp_elements(1);
    branch_req_2354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => if_stmt_481_branch_req_0); -- 
    -- CP-element group 36 branch  place  bypass 
    -- predecessors 35 
    -- successors 37 39 
    -- members (1) 
      -- 	branch_block_stmt_377/simple_obj_ref_482_place
      -- 
    cp_elements(36) <= cp_elements(35);
    -- CP-element group 37 transition  bypass 
    -- predecessors 36 
    -- successors 38 
    -- members (1) 
      -- 	branch_block_stmt_377/if_stmt_481_if_link/$entry
      -- 
    cp_elements(37) <= cp_elements(36);
    -- CP-element group 38 transition  place  input  no-bypass 
    -- predecessors 37 
    -- successors 2 
    -- members (9) 
      -- 	branch_block_stmt_377/if_stmt_481_if_link/$exit
      -- 	branch_block_stmt_377/if_stmt_481_if_link/if_choice_transition
      -- 	branch_block_stmt_377/bb_1_bb_2
      -- 	branch_block_stmt_377/merge_stmt_487_PhiReqMerge
      -- 	branch_block_stmt_377/bb_1_bb_2_PhiReq/$entry
      -- 	branch_block_stmt_377/bb_1_bb_2_PhiReq/$exit
      -- 	branch_block_stmt_377/merge_stmt_487_PhiAck/$entry
      -- 	branch_block_stmt_377/merge_stmt_487_PhiAck/$exit
      -- 	branch_block_stmt_377/merge_stmt_487_PhiAck/dummy
      -- 
    if_choice_transition_2359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_481_branch_ack_1, ack => cp_elements(38)); -- 
    -- CP-element group 39 transition  bypass 
    -- predecessors 36 
    -- successors 40 
    -- members (1) 
      -- 	branch_block_stmt_377/if_stmt_481_else_link/$entry
      -- 
    cp_elements(39) <= cp_elements(36);
    -- CP-element group 40 transition  place  input  no-bypass 
    -- predecessors 39 
    -- successors 
    -- members (21) 
      -- 	$exit
      -- 	branch_block_stmt_377/$exit
      -- 	branch_block_stmt_377/branch_block_stmt_377__exit__
      -- 	branch_block_stmt_377/merge_stmt_1179_PhiReqMerge
      -- 	branch_block_stmt_377/merge_stmt_1179__exit__
      -- 	branch_block_stmt_377/return__
      -- 	branch_block_stmt_377/merge_stmt_1181__exit__
      -- 	branch_block_stmt_377/if_stmt_481_else_link/$exit
      -- 	branch_block_stmt_377/if_stmt_481_else_link/else_choice_transition
      -- 	branch_block_stmt_377/bb_1_bb_4
      -- 	branch_block_stmt_377/merge_stmt_1181_PhiReqMerge
      -- 	branch_block_stmt_377/bb_1_bb_4_PhiReq/$entry
      -- 	branch_block_stmt_377/bb_1_bb_4_PhiReq/$exit
      -- 	branch_block_stmt_377/merge_stmt_1179_PhiAck/$entry
      -- 	branch_block_stmt_377/merge_stmt_1179_PhiAck/$exit
      -- 	branch_block_stmt_377/merge_stmt_1179_PhiAck/dummy
      -- 	branch_block_stmt_377/return___PhiReq/$entry
      -- 	branch_block_stmt_377/return___PhiReq/$exit
      -- 	branch_block_stmt_377/merge_stmt_1181_PhiAck/$entry
      -- 	branch_block_stmt_377/merge_stmt_1181_PhiAck/$exit
      -- 	branch_block_stmt_377/merge_stmt_1181_PhiAck/dummy
      -- 
    else_choice_transition_2363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_481_branch_ack_0, ack => cp_elements(40)); -- 
    -- CP-element group 41 fork  transition  bypass 
    -- predecessors 2 
    -- successors 42 50 58 66 74 82 90 98 106 114 122 130 138 146 154 162 170 178 186 194 202 210 218 231 239 253 260 269 277 291 299 313 320 329 337 351 359 373 380 389 397 411 419 433 440 449 457 471 479 493 500 509 517 531 539 553 560 569 577 591 599 613 620 629 637 651 659 673 680 689 696 704 720 728 736 752 760 768 784 792 800 816 824 832 848 856 864 880 888 896 912 920 928 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/$entry
      -- 
    cp_elements(41) <= cp_elements(2);
    -- CP-element group 42 transition  output  bypass 
    -- predecessors 41 
    -- successors 43 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_489_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_489_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_489_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_addr_resize/base_resize_req
      -- 
    cp_elements(42) <= cp_elements(41);
    base_resize_req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_490_base_resize_req_0); -- 
    -- CP-element group 43 transition  input  output  no-bypass 
    -- predecessors 42 
    -- successors 44 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_base_resize_ack_0, ack => cp_elements(43)); -- 
    sum_rename_req_2390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_490_root_address_inst_req_0); -- 
    -- CP-element group 44 transition  input  output  no-bypass 
    -- predecessors 43 
    -- successors 45 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_root_address_inst_ack_0, ack => cp_elements(44)); -- 
    root_register_req_2395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_490_addr_0_req_0); -- 
    -- CP-element group 45 transition  input  output  no-bypass 
    -- predecessors 44 
    -- successors 46 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/word_access_0/rr
      -- 
    root_register_ack_2396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_addr_0_ack_0, ack => cp_elements(45)); -- 
    rr_2406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_490_load_0_req_0); -- 
    -- CP-element group 46 transition  input  output  no-bypass 
    -- predecessors 45 
    -- successors 47 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/word_access_0/cr
      -- 
    ra_2407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_load_0_ack_0, ack => cp_elements(46)); -- 
    cr_2417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_490_load_0_req_1); -- 
    -- CP-element group 47 transition  input  output  no-bypass 
    -- predecessors 46 
    -- successors 48 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/merge_req
      -- 
    ca_2418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_load_0_ack_1, ack => cp_elements(47)); -- 
    merge_req_2419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_490_gather_scatter_req_0); -- 
    -- CP-element group 48 transition  input  output  no-bypass 
    -- predecessors 47 
    -- successors 49 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_491_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_491_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_491_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_490_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_493_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_493_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_493_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_complete/req
      -- 
    merge_ack_2420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_490_gather_scatter_ack_0, ack => cp_elements(48)); -- 
    req_2433_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => type_cast_494_inst_req_0); -- 
    -- CP-element group 49 fork  transition  input  no-bypass 
    -- predecessors 48 
    -- successors 52 53 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_495_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_495_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_495_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_494_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_497_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_497_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_497_completed_
      -- 
    ack_2434_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_494_inst_ack_0, ack => cp_elements(49)); -- 
    -- CP-element group 50 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_active_
      -- 
    cp_elements(50) <= cp_elements(41);
    -- CP-element group 51 join  transition  output  bypass 
    -- predecessors 54 55 
    -- successors 56 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_501_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_501_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_501_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_503_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_503_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_503_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_complete/req
      -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(54);
      predecessors(1) <= cp_elements(55);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(51)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => type_cast_504_inst_req_0); -- 
    -- CP-element group 52 transition  output  bypass 
    -- predecessors 49 
    -- successors 54 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Sample/rr
      -- 
    cp_elements(52) <= cp_elements(49);
    rr_2451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_500_inst_req_0); -- 
    -- CP-element group 53 transition  output  bypass 
    -- predecessors 49 
    -- successors 55 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Update/cr
      -- 
    cp_elements(53) <= cp_elements(49);
    cr_2456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => binary_500_inst_req_1); -- 
    -- CP-element group 54 transition  input  no-bypass 
    -- predecessors 52 
    -- successors 51 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Sample/ra
      -- 
    ra_2452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_500_inst_ack_0, ack => cp_elements(54)); -- 
    -- CP-element group 55 transition  input  no-bypass 
    -- predecessors 53 
    -- successors 51 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_500_Update/ca
      -- 
    ca_2457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_500_inst_ack_1, ack => cp_elements(55)); -- 
    -- CP-element group 56 transition  input  no-bypass 
    -- predecessors 51 
    -- successors 57 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_505_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_505_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_505_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_504_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_509_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_509_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_508_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_508_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_508_completed_
      -- 
    ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_504_inst_ack_0, ack => cp_elements(56)); -- 
    -- CP-element group 57 join  transition  output  bypass 
    -- predecessors 56 61 
    -- successors 62 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/split_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_trigger_
      -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(56);
      predecessors(1) <= cp_elements(61);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(57)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => ptr_deref_507_gather_scatter_req_0); -- 
    -- CP-element group 58 transition  output  bypass 
    -- predecessors 41 
    -- successors 59 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_506_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_506_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_506_active_
      -- 
    cp_elements(58) <= cp_elements(41);
    base_resize_req_2491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_507_base_resize_req_0); -- 
    -- CP-element group 59 transition  input  output  no-bypass 
    -- predecessors 58 
    -- successors 60 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_base_resize_ack_0, ack => cp_elements(59)); -- 
    sum_rename_req_2496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_507_root_address_inst_req_0); -- 
    -- CP-element group 60 transition  input  output  no-bypass 
    -- predecessors 59 
    -- successors 61 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_root_address_inst_ack_0, ack => cp_elements(60)); -- 
    root_register_req_2501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => ptr_deref_507_addr_0_req_0); -- 
    -- CP-element group 61 transition  input  no-bypass 
    -- predecessors 60 
    -- successors 57 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_word_address_calculated
      -- 
    root_register_ack_2502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_addr_0_ack_0, ack => cp_elements(61)); -- 
    -- CP-element group 62 transition  input  output  no-bypass 
    -- predecessors 57 
    -- successors 63 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/word_access_0/rr
      -- 
    split_ack_2507_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_gather_scatter_ack_0, ack => cp_elements(62)); -- 
    rr_2514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_507_store_0_req_0); -- 
    -- CP-element group 63 fork  transition  input  no-bypass 
    -- predecessors 62 
    -- successors 64 268 290 727 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_active_
      -- 
    ra_2515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_store_0_ack_0, ack => cp_elements(63)); -- 
    -- CP-element group 64 transition  output  bypass 
    -- predecessors 63 
    -- successors 65 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/word_access_0/cr
      -- 
    cp_elements(64) <= cp_elements(63);
    cr_2525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_507_store_0_req_1); -- 
    -- CP-element group 65 transition  input  no-bypass 
    -- predecessors 64 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_509_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_507_completed_
      -- 
    ca_2526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_507_store_0_ack_1, ack => cp_elements(65)); -- 
    -- CP-element group 66 transition  output  bypass 
    -- predecessors 41 
    -- successors 67 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_511_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_511_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_511_trigger_
      -- 
    cp_elements(66) <= cp_elements(41);
    base_resize_req_2543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => ptr_deref_512_base_resize_req_0); -- 
    -- CP-element group 67 transition  input  output  no-bypass 
    -- predecessors 66 
    -- successors 68 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_plus_offset/$entry
      -- 
    base_resize_ack_2544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_base_resize_ack_0, ack => cp_elements(67)); -- 
    sum_rename_req_2548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_512_root_address_inst_req_0); -- 
    -- CP-element group 68 transition  input  output  no-bypass 
    -- predecessors 67 
    -- successors 69 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_word_addrgen/$entry
      -- 
    sum_rename_ack_2549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_root_address_inst_ack_0, ack => cp_elements(68)); -- 
    root_register_req_2553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_512_addr_0_req_0); -- 
    -- CP-element group 69 transition  input  output  no-bypass 
    -- predecessors 68 
    -- successors 70 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_trigger_
      -- 
    root_register_ack_2554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_addr_0_ack_0, ack => cp_elements(69)); -- 
    rr_2564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_512_load_0_req_0); -- 
    -- CP-element group 70 transition  input  output  no-bypass 
    -- predecessors 69 
    -- successors 71 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_active_
      -- 
    ra_2565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_load_0_ack_0, ack => cp_elements(70)); -- 
    cr_2575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_512_load_0_req_1); -- 
    -- CP-element group 71 transition  input  output  no-bypass 
    -- predecessors 70 
    -- successors 72 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/merge_req
      -- 
    ca_2576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_load_0_ack_1, ack => cp_elements(71)); -- 
    merge_req_2577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_512_gather_scatter_req_0); -- 
    -- CP-element group 72 transition  input  output  no-bypass 
    -- predecessors 71 
    -- successors 73 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_515_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_515_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_513_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_515_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_513_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_513_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_512_completed_
      -- 
    merge_ack_2578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_512_gather_scatter_ack_0, ack => cp_elements(72)); -- 
    req_2591_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => type_cast_516_inst_req_0); -- 
    -- CP-element group 73 fork  transition  input  no-bypass 
    -- predecessors 72 
    -- successors 76 77 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_519_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_519_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_519_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_517_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_517_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_517_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_516_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_trigger_
      -- 
    ack_2592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_516_inst_ack_0, ack => cp_elements(73)); -- 
    -- CP-element group 74 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_active_
      -- 
    cp_elements(74) <= cp_elements(41);
    -- CP-element group 75 join  transition  output  bypass 
    -- predecessors 78 79 
    -- successors 80 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_525_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_525_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_525_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_523_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_523_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_523_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_completed_
      -- 
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(78);
      predecessors(1) <= cp_elements(79);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(75)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => type_cast_526_inst_req_0); -- 
    -- CP-element group 76 transition  output  bypass 
    -- predecessors 73 
    -- successors 78 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Sample/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_sample_start_
      -- 
    cp_elements(76) <= cp_elements(73);
    rr_2609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => binary_522_inst_req_0); -- 
    -- CP-element group 77 transition  output  bypass 
    -- predecessors 73 
    -- successors 79 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Update/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_update_start_
      -- 
    cp_elements(77) <= cp_elements(73);
    cr_2614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => binary_522_inst_req_1); -- 
    -- CP-element group 78 transition  input  no-bypass 
    -- predecessors 76 
    -- successors 75 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Sample/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_sample_completed_
      -- 
    ra_2610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_522_inst_ack_0, ack => cp_elements(78)); -- 
    -- CP-element group 79 transition  input  no-bypass 
    -- predecessors 77 
    -- successors 75 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Update/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_522_Update/$exit
      -- 
    ca_2615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_522_inst_ack_1, ack => cp_elements(79)); -- 
    -- CP-element group 80 transition  input  no-bypass 
    -- predecessors 75 
    -- successors 81 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_530_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_530_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_527_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_527_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_527_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_531_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_530_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_526_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_531_trigger_
      -- 
    ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_526_inst_ack_0, ack => cp_elements(80)); -- 
    -- CP-element group 81 join  transition  output  bypass 
    -- predecessors 80 85 
    -- successors 86 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/split_req
      -- 
    cpelement_group_81 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(80);
      predecessors(1) <= cp_elements(85);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(81)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(81),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_529_gather_scatter_req_0); -- 
    -- CP-element group 82 transition  output  bypass 
    -- predecessors 41 
    -- successors 83 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_528_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_528_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_528_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_address_calculated
      -- 
    cp_elements(82) <= cp_elements(41);
    base_resize_req_2649_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_529_base_resize_req_0); -- 
    -- CP-element group 83 transition  input  output  no-bypass 
    -- predecessors 82 
    -- successors 84 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_base_resize_ack_0, ack => cp_elements(83)); -- 
    sum_rename_req_2654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_529_root_address_inst_req_0); -- 
    -- CP-element group 84 transition  input  output  no-bypass 
    -- predecessors 83 
    -- successors 85 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_root_address_inst_ack_0, ack => cp_elements(84)); -- 
    root_register_req_2659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_529_addr_0_req_0); -- 
    -- CP-element group 85 transition  input  no-bypass 
    -- predecessors 84 
    -- successors 81 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_word_addrgen/root_register_ack
      -- 
    root_register_ack_2660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_addr_0_ack_0, ack => cp_elements(85)); -- 
    -- CP-element group 86 transition  input  output  no-bypass 
    -- predecessors 81 
    -- successors 87 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/word_access_0/rr
      -- 
    split_ack_2665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_gather_scatter_ack_0, ack => cp_elements(86)); -- 
    rr_2672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_529_store_0_req_0); -- 
    -- CP-element group 87 fork  transition  input  no-bypass 
    -- predecessors 86 
    -- successors 88 328 350 759 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_request/$exit
      -- 
    ra_2673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_store_0_ack_0, ack => cp_elements(87)); -- 
    -- CP-element group 88 transition  output  bypass 
    -- predecessors 87 
    -- successors 89 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/word_access_0/cr
      -- 
    cp_elements(88) <= cp_elements(87);
    cr_2683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_529_store_0_req_1); -- 
    -- CP-element group 89 transition  input  no-bypass 
    -- predecessors 88 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_529_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_531_completed_
      -- 
    ca_2684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_529_store_0_ack_1, ack => cp_elements(89)); -- 
    -- CP-element group 90 transition  output  bypass 
    -- predecessors 41 
    -- successors 91 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_533_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_533_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_533_trigger_
      -- 
    cp_elements(90) <= cp_elements(41);
    base_resize_req_2701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => ptr_deref_534_base_resize_req_0); -- 
    -- CP-element group 91 transition  input  output  no-bypass 
    -- predecessors 90 
    -- successors 92 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_base_resize_ack_0, ack => cp_elements(91)); -- 
    sum_rename_req_2706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => ptr_deref_534_root_address_inst_req_0); -- 
    -- CP-element group 92 transition  input  output  no-bypass 
    -- predecessors 91 
    -- successors 93 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_word_addrgen/$entry
      -- 
    sum_rename_ack_2707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_root_address_inst_ack_0, ack => cp_elements(92)); -- 
    root_register_req_2711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_534_addr_0_req_0); -- 
    -- CP-element group 93 transition  input  output  no-bypass 
    -- predecessors 92 
    -- successors 94 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_word_addrgen/$exit
      -- 
    root_register_ack_2712_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_addr_0_ack_0, ack => cp_elements(93)); -- 
    rr_2722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_534_load_0_req_0); -- 
    -- CP-element group 94 transition  input  output  no-bypass 
    -- predecessors 93 
    -- successors 95 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_request/word_access/word_access_0/ra
      -- 
    ra_2723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_load_0_ack_0, ack => cp_elements(94)); -- 
    cr_2733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_534_load_0_req_1); -- 
    -- CP-element group 95 transition  input  output  no-bypass 
    -- predecessors 94 
    -- successors 96 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/merge_req
      -- 
    ca_2734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_load_0_ack_1, ack => cp_elements(95)); -- 
    merge_req_2735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_534_gather_scatter_req_0); -- 
    -- CP-element group 96 transition  input  output  no-bypass 
    -- predecessors 95 
    -- successors 97 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_537_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_537_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_535_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_535_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_534_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_535_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_537_trigger_
      -- 
    merge_ack_2736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_534_gather_scatter_ack_0, ack => cp_elements(96)); -- 
    req_2749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => type_cast_538_inst_req_0); -- 
    -- CP-element group 97 fork  transition  input  no-bypass 
    -- predecessors 96 
    -- successors 100 101 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_539_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_539_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_539_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_541_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_541_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_538_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_541_completed_
      -- 
    ack_2750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => cp_elements(97)); -- 
    -- CP-element group 98 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_active_
      -- 
    cp_elements(98) <= cp_elements(41);
    -- CP-element group 99 join  transition  output  bypass 
    -- predecessors 102 103 
    -- successors 104 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_545_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_545_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_547_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_547_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_545_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_547_active_
      -- 
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(102);
      predecessors(1) <= cp_elements(103);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(99)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => type_cast_548_inst_req_0); -- 
    -- CP-element group 100 transition  output  bypass 
    -- predecessors 97 
    -- successors 102 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Sample/rr
      -- 
    cp_elements(100) <= cp_elements(97);
    rr_2767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => binary_544_inst_req_0); -- 
    -- CP-element group 101 transition  output  bypass 
    -- predecessors 97 
    -- successors 103 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Update/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Update/$entry
      -- 
    cp_elements(101) <= cp_elements(97);
    cr_2772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => binary_544_inst_req_1); -- 
    -- CP-element group 102 transition  input  no-bypass 
    -- predecessors 100 
    -- successors 99 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Sample/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_sample_completed_
      -- 
    ra_2768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_544_inst_ack_0, ack => cp_elements(102)); -- 
    -- CP-element group 103 transition  input  no-bypass 
    -- predecessors 101 
    -- successors 99 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_544_Update/ca
      -- 
    ca_2773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_544_inst_ack_1, ack => cp_elements(103)); -- 
    -- CP-element group 104 transition  input  no-bypass 
    -- predecessors 99 
    -- successors 105 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_552_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_549_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_549_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_549_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_552_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_552_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_553_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_553_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_548_completed_
      -- 
    ack_2787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_548_inst_ack_0, ack => cp_elements(104)); -- 
    -- CP-element group 105 join  transition  output  bypass 
    -- predecessors 104 109 
    -- successors 110 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/split_req
      -- 
    cpelement_group_105 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(104);
      predecessors(1) <= cp_elements(109);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(105)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(105),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_551_gather_scatter_req_0); -- 
    -- CP-element group 106 transition  output  bypass 
    -- predecessors 41 
    -- successors 107 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_550_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_550_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_550_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_addr_resize/$entry
      -- 
    cp_elements(106) <= cp_elements(41);
    base_resize_req_2807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_551_base_resize_req_0); -- 
    -- CP-element group 107 transition  input  output  no-bypass 
    -- predecessors 106 
    -- successors 108 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_addr_resize/$exit
      -- 
    base_resize_ack_2808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_base_resize_ack_0, ack => cp_elements(107)); -- 
    sum_rename_req_2812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_551_root_address_inst_req_0); -- 
    -- CP-element group 108 transition  input  output  no-bypass 
    -- predecessors 107 
    -- successors 109 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_base_plus_offset/$exit
      -- 
    sum_rename_ack_2813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_root_address_inst_ack_0, ack => cp_elements(108)); -- 
    root_register_req_2817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => ptr_deref_551_addr_0_req_0); -- 
    -- CP-element group 109 transition  input  no-bypass 
    -- predecessors 108 
    -- successors 105 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_word_addrgen/root_register_ack
      -- 
    root_register_ack_2818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_addr_0_ack_0, ack => cp_elements(109)); -- 
    -- CP-element group 110 transition  input  output  no-bypass 
    -- predecessors 105 
    -- successors 111 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/word_access_0/$entry
      -- 
    split_ack_2823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    rr_2830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_551_store_0_req_0); -- 
    -- CP-element group 111 fork  transition  input  no-bypass 
    -- predecessors 110 
    -- successors 112 388 410 791 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_request/word_access/$exit
      -- 
    ra_2831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_store_0_ack_0, ack => cp_elements(111)); -- 
    -- CP-element group 112 transition  output  bypass 
    -- predecessors 111 
    -- successors 113 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/word_access_0/$entry
      -- 
    cp_elements(112) <= cp_elements(111);
    cr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => ptr_deref_551_store_0_req_1); -- 
    -- CP-element group 113 transition  input  no-bypass 
    -- predecessors 112 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_553_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_551_complete/word_access/word_access_0/$exit
      -- 
    ca_2842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_551_store_0_ack_1, ack => cp_elements(113)); -- 
    -- CP-element group 114 transition  output  bypass 
    -- predecessors 41 
    -- successors 115 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_555_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_555_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_555_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_addr_resize/base_resize_req
      -- 
    cp_elements(114) <= cp_elements(41);
    base_resize_req_2859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_556_base_resize_req_0); -- 
    -- CP-element group 115 transition  input  output  no-bypass 
    -- predecessors 114 
    -- successors 116 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_base_resize_ack_0, ack => cp_elements(115)); -- 
    sum_rename_req_2864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_556_root_address_inst_req_0); -- 
    -- CP-element group 116 transition  input  output  no-bypass 
    -- predecessors 115 
    -- successors 117 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_root_address_inst_ack_0, ack => cp_elements(116)); -- 
    root_register_req_2869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => ptr_deref_556_addr_0_req_0); -- 
    -- CP-element group 117 transition  input  output  no-bypass 
    -- predecessors 116 
    -- successors 118 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/word_access_0/rr
      -- 
    root_register_ack_2870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_addr_0_ack_0, ack => cp_elements(117)); -- 
    rr_2880_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_556_load_0_req_0); -- 
    -- CP-element group 118 transition  input  output  no-bypass 
    -- predecessors 117 
    -- successors 119 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/word_access_0/cr
      -- 
    ra_2881_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_load_0_ack_0, ack => cp_elements(118)); -- 
    cr_2891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => ptr_deref_556_load_0_req_1); -- 
    -- CP-element group 119 transition  input  output  no-bypass 
    -- predecessors 118 
    -- successors 120 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/merge_req
      -- 
    ca_2892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_load_0_ack_1, ack => cp_elements(119)); -- 
    merge_req_2893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_556_gather_scatter_req_0); -- 
    -- CP-element group 120 transition  input  output  no-bypass 
    -- predecessors 119 
    -- successors 121 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_557_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_557_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_557_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_556_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_559_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_559_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_559_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_complete/req
      -- 
    merge_ack_2894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_556_gather_scatter_ack_0, ack => cp_elements(120)); -- 
    req_2907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => type_cast_560_inst_req_0); -- 
    -- CP-element group 121 fork  transition  input  no-bypass 
    -- predecessors 120 
    -- successors 124 125 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_561_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_561_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_561_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_560_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_563_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_563_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_563_completed_
      -- 
    ack_2908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_560_inst_ack_0, ack => cp_elements(121)); -- 
    -- CP-element group 122 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_active_
      -- 
    cp_elements(122) <= cp_elements(41);
    -- CP-element group 123 join  transition  output  bypass 
    -- predecessors 126 127 
    -- successors 128 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_567_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_567_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_567_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_569_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_569_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_569_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_complete/req
      -- 
    cpelement_group_123 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(126);
      predecessors(1) <= cp_elements(127);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(123)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(123),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => type_cast_570_inst_req_0); -- 
    -- CP-element group 124 transition  output  bypass 
    -- predecessors 121 
    -- successors 126 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Sample/rr
      -- 
    cp_elements(124) <= cp_elements(121);
    rr_2925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => binary_566_inst_req_0); -- 
    -- CP-element group 125 transition  output  bypass 
    -- predecessors 121 
    -- successors 127 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Update/cr
      -- 
    cp_elements(125) <= cp_elements(121);
    cr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => binary_566_inst_req_1); -- 
    -- CP-element group 126 transition  input  no-bypass 
    -- predecessors 124 
    -- successors 123 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Sample/ra
      -- 
    ra_2926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_566_inst_ack_0, ack => cp_elements(126)); -- 
    -- CP-element group 127 transition  input  no-bypass 
    -- predecessors 125 
    -- successors 123 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_566_Update/ca
      -- 
    ca_2931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_566_inst_ack_1, ack => cp_elements(127)); -- 
    -- CP-element group 128 transition  input  no-bypass 
    -- predecessors 123 
    -- successors 129 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_571_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_571_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_571_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_570_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_575_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_575_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_574_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_574_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_574_completed_
      -- 
    ack_2945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_570_inst_ack_0, ack => cp_elements(128)); -- 
    -- CP-element group 129 join  transition  output  bypass 
    -- predecessors 128 133 
    -- successors 134 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/split_req
      -- 
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(128);
      predecessors(1) <= cp_elements(133);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(129)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_573_gather_scatter_req_0); -- 
    -- CP-element group 130 transition  output  bypass 
    -- predecessors 41 
    -- successors 131 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_572_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_572_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_572_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_addr_resize/base_resize_req
      -- 
    cp_elements(130) <= cp_elements(41);
    base_resize_req_2965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => ptr_deref_573_base_resize_req_0); -- 
    -- CP-element group 131 transition  input  output  no-bypass 
    -- predecessors 130 
    -- successors 132 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_2966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_base_resize_ack_0, ack => cp_elements(131)); -- 
    sum_rename_req_2970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_573_root_address_inst_req_0); -- 
    -- CP-element group 132 transition  input  output  no-bypass 
    -- predecessors 131 
    -- successors 133 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_word_addrgen/root_register_req
      -- 
    sum_rename_ack_2971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_root_address_inst_ack_0, ack => cp_elements(132)); -- 
    root_register_req_2975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_573_addr_0_req_0); -- 
    -- CP-element group 133 transition  input  no-bypass 
    -- predecessors 132 
    -- successors 129 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_word_addrgen/root_register_ack
      -- 
    root_register_ack_2976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_addr_0_ack_0, ack => cp_elements(133)); -- 
    -- CP-element group 134 transition  input  output  no-bypass 
    -- predecessors 129 
    -- successors 135 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/word_access_0/rr
      -- 
    split_ack_2981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_gather_scatter_ack_0, ack => cp_elements(134)); -- 
    rr_2988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_573_store_0_req_0); -- 
    -- CP-element group 135 fork  transition  input  no-bypass 
    -- predecessors 134 
    -- successors 136 448 470 823 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_request/word_access/word_access_0/ra
      -- 
    ra_2989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_store_0_ack_0, ack => cp_elements(135)); -- 
    -- CP-element group 136 transition  output  bypass 
    -- predecessors 135 
    -- successors 137 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/word_access_0/cr
      -- 
    cp_elements(136) <= cp_elements(135);
    cr_2999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => ptr_deref_573_store_0_req_1); -- 
    -- CP-element group 137 transition  input  no-bypass 
    -- predecessors 136 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_575_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_573_complete/word_access/word_access_0/ca
      -- 
    ca_3000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_573_store_0_ack_1, ack => cp_elements(137)); -- 
    -- CP-element group 138 transition  output  bypass 
    -- predecessors 41 
    -- successors 139 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_577_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_577_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_577_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_addr_resize/base_resize_req
      -- 
    cp_elements(138) <= cp_elements(41);
    base_resize_req_3017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_578_base_resize_req_0); -- 
    -- CP-element group 139 transition  input  output  no-bypass 
    -- predecessors 138 
    -- successors 140 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_base_resize_ack_0, ack => cp_elements(139)); -- 
    sum_rename_req_3022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => ptr_deref_578_root_address_inst_req_0); -- 
    -- CP-element group 140 transition  input  output  no-bypass 
    -- predecessors 139 
    -- successors 141 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_root_address_inst_ack_0, ack => cp_elements(140)); -- 
    root_register_req_3027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_578_addr_0_req_0); -- 
    -- CP-element group 141 transition  input  output  no-bypass 
    -- predecessors 140 
    -- successors 142 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_addr_0_ack_0, ack => cp_elements(141)); -- 
    rr_3038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(141), ack => ptr_deref_578_load_0_req_0); -- 
    -- CP-element group 142 transition  input  output  no-bypass 
    -- predecessors 141 
    -- successors 143 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/word_access_0/cr
      -- 
    ra_3039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_load_0_ack_0, ack => cp_elements(142)); -- 
    cr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_578_load_0_req_1); -- 
    -- CP-element group 143 transition  input  output  no-bypass 
    -- predecessors 142 
    -- successors 144 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/merge_req
      -- 
    ca_3050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_load_0_ack_1, ack => cp_elements(143)); -- 
    merge_req_3051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => ptr_deref_578_gather_scatter_req_0); -- 
    -- CP-element group 144 transition  input  output  no-bypass 
    -- predecessors 143 
    -- successors 145 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_579_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_579_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_579_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_578_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_581_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_581_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_581_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_complete/req
      -- 
    merge_ack_3052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_578_gather_scatter_ack_0, ack => cp_elements(144)); -- 
    req_3065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => type_cast_582_inst_req_0); -- 
    -- CP-element group 145 fork  transition  input  no-bypass 
    -- predecessors 144 
    -- successors 148 149 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_583_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_583_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_583_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_582_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_585_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_585_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_585_completed_
      -- 
    ack_3066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_582_inst_ack_0, ack => cp_elements(145)); -- 
    -- CP-element group 146 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_active_
      -- 
    cp_elements(146) <= cp_elements(41);
    -- CP-element group 147 join  transition  output  bypass 
    -- predecessors 150 151 
    -- successors 152 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_589_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_589_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_589_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_591_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_591_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_591_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_complete/req
      -- 
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(150);
      predecessors(1) <= cp_elements(151);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(147)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => type_cast_592_inst_req_0); -- 
    -- CP-element group 148 transition  output  bypass 
    -- predecessors 145 
    -- successors 150 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Sample/rr
      -- 
    cp_elements(148) <= cp_elements(145);
    rr_3083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => binary_588_inst_req_0); -- 
    -- CP-element group 149 transition  output  bypass 
    -- predecessors 145 
    -- successors 151 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Update/cr
      -- 
    cp_elements(149) <= cp_elements(145);
    cr_3088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => binary_588_inst_req_1); -- 
    -- CP-element group 150 transition  input  no-bypass 
    -- predecessors 148 
    -- successors 147 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Sample/ra
      -- 
    ra_3084_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_0, ack => cp_elements(150)); -- 
    -- CP-element group 151 transition  input  no-bypass 
    -- predecessors 149 
    -- successors 147 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_588_Update/ca
      -- 
    ca_3089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_1, ack => cp_elements(151)); -- 
    -- CP-element group 152 transition  input  no-bypass 
    -- predecessors 147 
    -- successors 153 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_593_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_593_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_593_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_592_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_597_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_597_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_596_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_596_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_596_completed_
      -- 
    ack_3103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_592_inst_ack_0, ack => cp_elements(152)); -- 
    -- CP-element group 153 join  transition  output  bypass 
    -- predecessors 152 157 
    -- successors 158 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/split_req
      -- 
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(152);
      predecessors(1) <= cp_elements(157);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(153)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_595_gather_scatter_req_0); -- 
    -- CP-element group 154 transition  output  bypass 
    -- predecessors 41 
    -- successors 155 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_594_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_594_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_594_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_addr_resize/base_resize_req
      -- 
    cp_elements(154) <= cp_elements(41);
    base_resize_req_3123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => ptr_deref_595_base_resize_req_0); -- 
    -- CP-element group 155 transition  input  output  no-bypass 
    -- predecessors 154 
    -- successors 156 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3124_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_base_resize_ack_0, ack => cp_elements(155)); -- 
    sum_rename_req_3128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_595_root_address_inst_req_0); -- 
    -- CP-element group 156 transition  input  output  no-bypass 
    -- predecessors 155 
    -- successors 157 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_root_address_inst_ack_0, ack => cp_elements(156)); -- 
    root_register_req_3133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => ptr_deref_595_addr_0_req_0); -- 
    -- CP-element group 157 transition  input  no-bypass 
    -- predecessors 156 
    -- successors 153 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_word_addrgen/root_register_ack
      -- 
    root_register_ack_3134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_addr_0_ack_0, ack => cp_elements(157)); -- 
    -- CP-element group 158 transition  input  output  no-bypass 
    -- predecessors 153 
    -- successors 159 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/word_access_0/rr
      -- 
    split_ack_3139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_gather_scatter_ack_0, ack => cp_elements(158)); -- 
    rr_3146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => ptr_deref_595_store_0_req_0); -- 
    -- CP-element group 159 fork  transition  input  no-bypass 
    -- predecessors 158 
    -- successors 160 508 530 855 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_request/word_access/word_access_0/ra
      -- 
    ra_3147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_store_0_ack_0, ack => cp_elements(159)); -- 
    -- CP-element group 160 transition  output  bypass 
    -- predecessors 159 
    -- successors 161 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/word_access_0/cr
      -- 
    cp_elements(160) <= cp_elements(159);
    cr_3157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => ptr_deref_595_store_0_req_1); -- 
    -- CP-element group 161 transition  input  no-bypass 
    -- predecessors 160 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_597_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_595_complete/word_access/word_access_0/ca
      -- 
    ca_3158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_595_store_0_ack_1, ack => cp_elements(161)); -- 
    -- CP-element group 162 transition  output  bypass 
    -- predecessors 41 
    -- successors 163 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_599_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_599_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_599_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_addr_resize/base_resize_req
      -- 
    cp_elements(162) <= cp_elements(41);
    base_resize_req_3175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => ptr_deref_600_base_resize_req_0); -- 
    -- CP-element group 163 transition  input  output  no-bypass 
    -- predecessors 162 
    -- successors 164 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_base_resize_ack_0, ack => cp_elements(163)); -- 
    sum_rename_req_3180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => ptr_deref_600_root_address_inst_req_0); -- 
    -- CP-element group 164 transition  input  output  no-bypass 
    -- predecessors 163 
    -- successors 165 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_root_address_inst_ack_0, ack => cp_elements(164)); -- 
    root_register_req_3185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => ptr_deref_600_addr_0_req_0); -- 
    -- CP-element group 165 transition  input  output  no-bypass 
    -- predecessors 164 
    -- successors 166 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_addr_0_ack_0, ack => cp_elements(165)); -- 
    rr_3196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => ptr_deref_600_load_0_req_0); -- 
    -- CP-element group 166 transition  input  output  no-bypass 
    -- predecessors 165 
    -- successors 167 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/word_access_0/cr
      -- 
    ra_3197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_load_0_ack_0, ack => cp_elements(166)); -- 
    cr_3207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => ptr_deref_600_load_0_req_1); -- 
    -- CP-element group 167 transition  input  output  no-bypass 
    -- predecessors 166 
    -- successors 168 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/merge_req
      -- 
    ca_3208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_load_0_ack_1, ack => cp_elements(167)); -- 
    merge_req_3209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => ptr_deref_600_gather_scatter_req_0); -- 
    -- CP-element group 168 transition  input  output  no-bypass 
    -- predecessors 167 
    -- successors 169 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_601_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_601_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_601_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_600_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_603_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_603_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_603_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_complete/req
      -- 
    merge_ack_3210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_600_gather_scatter_ack_0, ack => cp_elements(168)); -- 
    req_3223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => type_cast_604_inst_req_0); -- 
    -- CP-element group 169 fork  transition  input  no-bypass 
    -- predecessors 168 
    -- successors 172 173 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_605_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_605_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_605_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_604_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_607_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_607_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_607_completed_
      -- 
    ack_3224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_604_inst_ack_0, ack => cp_elements(169)); -- 
    -- CP-element group 170 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_active_
      -- 
    cp_elements(170) <= cp_elements(41);
    -- CP-element group 171 join  transition  output  bypass 
    -- predecessors 174 175 
    -- successors 176 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_611_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_611_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_611_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_613_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_613_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_613_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_complete/req
      -- 
    cpelement_group_171 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(174);
      predecessors(1) <= cp_elements(175);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(171)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(171),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => type_cast_614_inst_req_0); -- 
    -- CP-element group 172 transition  output  bypass 
    -- predecessors 169 
    -- successors 174 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Sample/rr
      -- 
    cp_elements(172) <= cp_elements(169);
    rr_3241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(172), ack => binary_610_inst_req_0); -- 
    -- CP-element group 173 transition  output  bypass 
    -- predecessors 169 
    -- successors 175 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Update/cr
      -- 
    cp_elements(173) <= cp_elements(169);
    cr_3246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => binary_610_inst_req_1); -- 
    -- CP-element group 174 transition  input  no-bypass 
    -- predecessors 172 
    -- successors 171 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Sample/ra
      -- 
    ra_3242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_610_inst_ack_0, ack => cp_elements(174)); -- 
    -- CP-element group 175 transition  input  no-bypass 
    -- predecessors 173 
    -- successors 171 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_610_Update/ca
      -- 
    ca_3247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_610_inst_ack_1, ack => cp_elements(175)); -- 
    -- CP-element group 176 transition  input  no-bypass 
    -- predecessors 171 
    -- successors 177 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_615_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_615_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_615_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_614_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_619_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_619_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_618_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_618_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_618_completed_
      -- 
    ack_3261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_614_inst_ack_0, ack => cp_elements(176)); -- 
    -- CP-element group 177 join  transition  output  bypass 
    -- predecessors 176 181 
    -- successors 182 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/split_req
      -- 
    cpelement_group_177 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(176);
      predecessors(1) <= cp_elements(181);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(177)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => ptr_deref_617_gather_scatter_req_0); -- 
    -- CP-element group 178 transition  output  bypass 
    -- predecessors 41 
    -- successors 179 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_616_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_616_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_616_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_addr_resize/base_resize_req
      -- 
    cp_elements(178) <= cp_elements(41);
    base_resize_req_3281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => ptr_deref_617_base_resize_req_0); -- 
    -- CP-element group 179 transition  input  output  no-bypass 
    -- predecessors 178 
    -- successors 180 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_base_resize_ack_0, ack => cp_elements(179)); -- 
    sum_rename_req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => ptr_deref_617_root_address_inst_req_0); -- 
    -- CP-element group 180 transition  input  output  no-bypass 
    -- predecessors 179 
    -- successors 181 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_root_address_inst_ack_0, ack => cp_elements(180)); -- 
    root_register_req_3291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => ptr_deref_617_addr_0_req_0); -- 
    -- CP-element group 181 transition  input  no-bypass 
    -- predecessors 180 
    -- successors 177 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_word_addrgen/root_register_ack
      -- 
    root_register_ack_3292_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_addr_0_ack_0, ack => cp_elements(181)); -- 
    -- CP-element group 182 transition  input  output  no-bypass 
    -- predecessors 177 
    -- successors 183 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/word_access_0/rr
      -- 
    split_ack_3297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_gather_scatter_ack_0, ack => cp_elements(182)); -- 
    rr_3304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(182), ack => ptr_deref_617_store_0_req_0); -- 
    -- CP-element group 183 fork  transition  input  no-bypass 
    -- predecessors 182 
    -- successors 184 568 590 887 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_request/word_access/word_access_0/ra
      -- 
    ra_3305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_store_0_ack_0, ack => cp_elements(183)); -- 
    -- CP-element group 184 transition  output  bypass 
    -- predecessors 183 
    -- successors 185 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/word_access_0/cr
      -- 
    cp_elements(184) <= cp_elements(183);
    cr_3315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(184), ack => ptr_deref_617_store_0_req_1); -- 
    -- CP-element group 185 transition  input  no-bypass 
    -- predecessors 184 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_619_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_617_complete/word_access/word_access_0/ca
      -- 
    ca_3316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_617_store_0_ack_1, ack => cp_elements(185)); -- 
    -- CP-element group 186 transition  output  bypass 
    -- predecessors 41 
    -- successors 187 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_621_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_621_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_621_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_addr_resize/base_resize_req
      -- 
    cp_elements(186) <= cp_elements(41);
    base_resize_req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => ptr_deref_622_base_resize_req_0); -- 
    -- CP-element group 187 transition  input  output  no-bypass 
    -- predecessors 186 
    -- successors 188 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_base_resize_ack_0, ack => cp_elements(187)); -- 
    sum_rename_req_3338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => ptr_deref_622_root_address_inst_req_0); -- 
    -- CP-element group 188 transition  input  output  no-bypass 
    -- predecessors 187 
    -- successors 189 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_root_address_inst_ack_0, ack => cp_elements(188)); -- 
    root_register_req_3343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_622_addr_0_req_0); -- 
    -- CP-element group 189 transition  input  output  no-bypass 
    -- predecessors 188 
    -- successors 190 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_addr_0_ack_0, ack => cp_elements(189)); -- 
    rr_3354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => ptr_deref_622_load_0_req_0); -- 
    -- CP-element group 190 transition  input  output  no-bypass 
    -- predecessors 189 
    -- successors 191 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/word_access_0/cr
      -- 
    ra_3355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_load_0_ack_0, ack => cp_elements(190)); -- 
    cr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_622_load_0_req_1); -- 
    -- CP-element group 191 transition  input  output  no-bypass 
    -- predecessors 190 
    -- successors 192 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/merge_req
      -- 
    ca_3366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_load_0_ack_1, ack => cp_elements(191)); -- 
    merge_req_3367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => ptr_deref_622_gather_scatter_req_0); -- 
    -- CP-element group 192 transition  input  output  no-bypass 
    -- predecessors 191 
    -- successors 193 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_623_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_623_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_623_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_622_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_625_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_625_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_625_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_complete/req
      -- 
    merge_ack_3368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_622_gather_scatter_ack_0, ack => cp_elements(192)); -- 
    req_3381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_626_inst_req_0); -- 
    -- CP-element group 193 fork  transition  input  no-bypass 
    -- predecessors 192 
    -- successors 196 197 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_627_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_627_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_627_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_626_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_629_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_629_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_629_completed_
      -- 
    ack_3382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_626_inst_ack_0, ack => cp_elements(193)); -- 
    -- CP-element group 194 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_active_
      -- 
    cp_elements(194) <= cp_elements(41);
    -- CP-element group 195 join  transition  output  bypass 
    -- predecessors 198 199 
    -- successors 200 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_633_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_633_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_633_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_635_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_635_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_635_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_complete/req
      -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(198);
      predecessors(1) <= cp_elements(199);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(195)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => type_cast_636_inst_req_0); -- 
    -- CP-element group 196 transition  output  bypass 
    -- predecessors 193 
    -- successors 198 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Sample/rr
      -- 
    cp_elements(196) <= cp_elements(193);
    rr_3399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => binary_632_inst_req_0); -- 
    -- CP-element group 197 transition  output  bypass 
    -- predecessors 193 
    -- successors 199 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Update/cr
      -- 
    cp_elements(197) <= cp_elements(193);
    cr_3404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_632_inst_req_1); -- 
    -- CP-element group 198 transition  input  no-bypass 
    -- predecessors 196 
    -- successors 195 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Sample/ra
      -- 
    ra_3400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_632_inst_ack_0, ack => cp_elements(198)); -- 
    -- CP-element group 199 transition  input  no-bypass 
    -- predecessors 197 
    -- successors 195 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_632_Update/ca
      -- 
    ca_3405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_632_inst_ack_1, ack => cp_elements(199)); -- 
    -- CP-element group 200 transition  input  no-bypass 
    -- predecessors 195 
    -- successors 201 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_637_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_637_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_637_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_636_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_641_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_641_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_640_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_640_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_640_completed_
      -- 
    ack_3419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_636_inst_ack_0, ack => cp_elements(200)); -- 
    -- CP-element group 201 join  transition  output  bypass 
    -- predecessors 200 205 
    -- successors 206 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/split_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_trigger_
      -- 
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(200);
      predecessors(1) <= cp_elements(205);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(201)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3454_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => ptr_deref_639_gather_scatter_req_0); -- 
    -- CP-element group 202 transition  output  bypass 
    -- predecessors 41 
    -- successors 203 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_638_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_638_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_638_completed_
      -- 
    cp_elements(202) <= cp_elements(41);
    base_resize_req_3439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(202), ack => ptr_deref_639_base_resize_req_0); -- 
    -- CP-element group 203 transition  input  output  no-bypass 
    -- predecessors 202 
    -- successors 204 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_address_resized
      -- 
    base_resize_ack_3440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_base_resize_ack_0, ack => cp_elements(203)); -- 
    sum_rename_req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => ptr_deref_639_root_address_inst_req_0); -- 
    -- CP-element group 204 transition  input  output  no-bypass 
    -- predecessors 203 
    -- successors 205 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_root_address_calculated
      -- 
    sum_rename_ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_root_address_inst_ack_0, ack => cp_elements(204)); -- 
    root_register_req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_639_addr_0_req_0); -- 
    -- CP-element group 205 transition  input  no-bypass 
    -- predecessors 204 
    -- successors 201 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_word_address_calculated
      -- 
    root_register_ack_3450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_addr_0_ack_0, ack => cp_elements(205)); -- 
    -- CP-element group 206 transition  input  output  no-bypass 
    -- predecessors 201 
    -- successors 207 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/word_access_0/rr
      -- 
    split_ack_3455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_gather_scatter_ack_0, ack => cp_elements(206)); -- 
    rr_3462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_639_store_0_req_0); -- 
    -- CP-element group 207 fork  transition  input  no-bypass 
    -- predecessors 206 
    -- successors 208 628 650 919 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_active_
      -- 
    ra_3463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_store_0_ack_0, ack => cp_elements(207)); -- 
    -- CP-element group 208 transition  output  bypass 
    -- predecessors 207 
    -- successors 209 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/word_access_0/cr
      -- 
    cp_elements(208) <= cp_elements(207);
    cr_3473_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => ptr_deref_639_store_0_req_1); -- 
    -- CP-element group 209 transition  input  no-bypass 
    -- predecessors 208 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_641_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_639_completed_
      -- 
    ca_3474_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_639_store_0_ack_1, ack => cp_elements(209)); -- 
    -- CP-element group 210 transition  output  bypass 
    -- predecessors 41 
    -- successors 211 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_643_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_643_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_643_trigger_
      -- 
    cp_elements(210) <= cp_elements(41);
    base_resize_req_3491_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_644_base_resize_req_0); -- 
    -- CP-element group 211 transition  input  output  no-bypass 
    -- predecessors 210 
    -- successors 212 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_addr_resize/$exit
      -- 
    base_resize_ack_3492_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_base_resize_ack_0, ack => cp_elements(211)); -- 
    sum_rename_req_3496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => ptr_deref_644_root_address_inst_req_0); -- 
    -- CP-element group 212 transition  input  output  no-bypass 
    -- predecessors 211 
    -- successors 213 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_root_address_inst_ack_0, ack => cp_elements(212)); -- 
    root_register_req_3501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_644_addr_0_req_0); -- 
    -- CP-element group 213 transition  input  output  no-bypass 
    -- predecessors 212 
    -- successors 214 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_addr_0_ack_0, ack => cp_elements(213)); -- 
    rr_3512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_644_load_0_req_0); -- 
    -- CP-element group 214 transition  input  output  no-bypass 
    -- predecessors 213 
    -- successors 215 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_request/word_access/word_access_0/ra
      -- 
    ra_3513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_load_0_ack_0, ack => cp_elements(214)); -- 
    cr_3523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => ptr_deref_644_load_0_req_1); -- 
    -- CP-element group 215 transition  input  output  no-bypass 
    -- predecessors 214 
    -- successors 216 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/merge_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/word_access/word_access_0/$exit
      -- 
    ca_3524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_load_0_ack_1, ack => cp_elements(215)); -- 
    merge_req_3525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => ptr_deref_644_gather_scatter_req_0); -- 
    -- CP-element group 216 transition  input  output  no-bypass 
    -- predecessors 215 
    -- successors 217 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_645_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_645_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_645_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_647_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_647_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_647_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_644_complete/merge_ack
      -- 
    merge_ack_3526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_644_gather_scatter_ack_0, ack => cp_elements(216)); -- 
    req_3539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(216), ack => type_cast_648_inst_req_0); -- 
    -- CP-element group 217 transition  input  output  no-bypass 
    -- predecessors 216 
    -- successors 220 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_resize_0/index_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_649_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_649_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_651_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_651_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_649_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_648_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_651_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_resize_0/$entry
      -- 
    ack_3540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_648_inst_ack_0, ack => cp_elements(217)); -- 
    index_resize_req_3558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => array_obj_ref_652_index_0_resize_req_0); -- 
    -- CP-element group 218 transition  bypass 
    -- predecessors 41 
    -- successors 219 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_trigger_
      -- 
    cp_elements(218) <= cp_elements(41);
    -- CP-element group 219 join  transition  output  no-bypass 
    -- predecessors 218 223 
    -- successors 224 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_complete/final_reg_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_complete/$entry
      -- 
    cpelement_group_219 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(218);
      predecessors(1) <= cp_elements(223);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(219)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(219),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => addr_of_653_final_reg_req_0); -- 
    -- CP-element group 220 transition  input  output  no-bypass 
    -- predecessors 217 
    -- successors 221 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_resize_0/$exit
      -- 
    index_resize_ack_3559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_652_index_0_resize_ack_0, ack => cp_elements(220)); -- 
    scale_rename_req_3563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(220), ack => array_obj_ref_652_index_0_rename_req_0); -- 
    -- CP-element group 221 transition  input  output  no-bypass 
    -- predecessors 220 
    -- successors 222 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_add_indices/final_index_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_add_indices/$entry
      -- 
    scale_rename_ack_3564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_652_index_0_rename_ack_0, ack => cp_elements(221)); -- 
    final_index_req_3568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => array_obj_ref_652_offset_inst_req_0); -- 
    -- CP-element group 222 transition  input  output  no-bypass 
    -- predecessors 221 
    -- successors 223 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_add_indices/$exit
      -- 
    final_index_ack_3569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_652_offset_inst_ack_0, ack => cp_elements(222)); -- 
    sum_rename_req_3573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => array_obj_ref_652_root_address_inst_req_0); -- 
    -- CP-element group 223 transition  input  no-bypass 
    -- predecessors 222 
    -- successors 219 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_652_base_plus_offset/$exit
      -- 
    sum_rename_ack_3574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_652_root_address_inst_ack_0, ack => cp_elements(223)); -- 
    -- CP-element group 224 transition  input  output  no-bypass 
    -- predecessors 219 
    -- successors 225 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_654_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_654_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_653_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_654_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_656_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_656_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_656_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_3579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_653_final_reg_ack_0, ack => cp_elements(224)); -- 
    base_resize_req_3596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_657_base_resize_req_0); -- 
    -- CP-element group 225 transition  input  output  no-bypass 
    -- predecessors 224 
    -- successors 226 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_base_resize_ack_0, ack => cp_elements(225)); -- 
    sum_rename_req_3601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => ptr_deref_657_root_address_inst_req_0); -- 
    -- CP-element group 226 transition  input  output  no-bypass 
    -- predecessors 225 
    -- successors 227 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_root_address_inst_ack_0, ack => cp_elements(226)); -- 
    root_register_req_3606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => ptr_deref_657_addr_0_req_0); -- 
    -- CP-element group 227 transition  input  output  no-bypass 
    -- predecessors 226 
    -- successors 228 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_addr_0_ack_0, ack => cp_elements(227)); -- 
    rr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => ptr_deref_657_load_0_req_0); -- 
    -- CP-element group 228 transition  input  output  no-bypass 
    -- predecessors 227 
    -- successors 229 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/word_access_0/cr
      -- 
    ra_3618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_load_0_ack_0, ack => cp_elements(228)); -- 
    cr_3628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => ptr_deref_657_load_0_req_1); -- 
    -- CP-element group 229 transition  input  output  no-bypass 
    -- predecessors 228 
    -- successors 230 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/merge_req
      -- 
    ca_3629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_load_0_ack_1, ack => cp_elements(229)); -- 
    merge_req_3630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => ptr_deref_657_gather_scatter_req_0); -- 
    -- CP-element group 230 transition  input  no-bypass 
    -- predecessors 229 
    -- successors 252 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_658_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_658_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_658_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_657_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_677_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_677_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_677_completed_
      -- 
    merge_ack_3631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_657_gather_scatter_ack_0, ack => cp_elements(230)); -- 
    -- CP-element group 231 transition  output  bypass 
    -- predecessors 41 
    -- successors 232 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_660_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_660_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_660_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_addr_resize/base_resize_req
      -- 
    cp_elements(231) <= cp_elements(41);
    base_resize_req_3648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_661_base_resize_req_0); -- 
    -- CP-element group 232 transition  input  output  no-bypass 
    -- predecessors 231 
    -- successors 233 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_base_resize_ack_0, ack => cp_elements(232)); -- 
    sum_rename_req_3653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(232), ack => ptr_deref_661_root_address_inst_req_0); -- 
    -- CP-element group 233 transition  input  output  no-bypass 
    -- predecessors 232 
    -- successors 234 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_root_address_inst_ack_0, ack => cp_elements(233)); -- 
    root_register_req_3658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_661_addr_0_req_0); -- 
    -- CP-element group 234 transition  input  output  no-bypass 
    -- predecessors 233 
    -- successors 235 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_addr_0_ack_0, ack => cp_elements(234)); -- 
    rr_3669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_661_load_0_req_0); -- 
    -- CP-element group 235 transition  input  output  no-bypass 
    -- predecessors 234 
    -- successors 236 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/word_access_0/cr
      -- 
    ra_3670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_load_0_ack_0, ack => cp_elements(235)); -- 
    cr_3680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => ptr_deref_661_load_0_req_1); -- 
    -- CP-element group 236 transition  input  output  no-bypass 
    -- predecessors 235 
    -- successors 237 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/merge_req
      -- 
    ca_3681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_load_0_ack_1, ack => cp_elements(236)); -- 
    merge_req_3682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_661_gather_scatter_req_0); -- 
    -- CP-element group 237 transition  input  output  no-bypass 
    -- predecessors 236 
    -- successors 238 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_662_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_662_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_662_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_661_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_664_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_664_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_664_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_complete/req
      -- 
    merge_ack_3683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_661_gather_scatter_ack_0, ack => cp_elements(237)); -- 
    req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => type_cast_665_inst_req_0); -- 
    -- CP-element group 238 transition  input  output  no-bypass 
    -- predecessors 237 
    -- successors 241 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_666_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_666_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_666_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_665_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_668_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_668_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_668_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_resize_0/index_resize_req
      -- 
    ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_665_inst_ack_0, ack => cp_elements(238)); -- 
    index_resize_req_3715_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => array_obj_ref_669_index_0_resize_req_0); -- 
    -- CP-element group 239 transition  bypass 
    -- predecessors 41 
    -- successors 240 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_trigger_
      -- 
    cp_elements(239) <= cp_elements(41);
    -- CP-element group 240 join  transition  output  no-bypass 
    -- predecessors 239 244 
    -- successors 245 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_complete/final_reg_req
      -- 
    cpelement_group_240 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(239);
      predecessors(1) <= cp_elements(244);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(240)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(240),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => addr_of_670_final_reg_req_0); -- 
    -- CP-element group 241 transition  input  output  no-bypass 
    -- predecessors 238 
    -- successors 242 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_669_index_0_resize_ack_0, ack => cp_elements(241)); -- 
    scale_rename_req_3720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => array_obj_ref_669_index_0_rename_req_0); -- 
    -- CP-element group 242 transition  input  output  no-bypass 
    -- predecessors 241 
    -- successors 243 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_add_indices/final_index_req
      -- 
    scale_rename_ack_3721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_669_index_0_rename_ack_0, ack => cp_elements(242)); -- 
    final_index_req_3725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => array_obj_ref_669_offset_inst_req_0); -- 
    -- CP-element group 243 transition  input  output  no-bypass 
    -- predecessors 242 
    -- successors 244 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_669_offset_inst_ack_0, ack => cp_elements(243)); -- 
    sum_rename_req_3730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(243), ack => array_obj_ref_669_root_address_inst_req_0); -- 
    -- CP-element group 244 transition  input  no-bypass 
    -- predecessors 243 
    -- successors 240 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_669_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_669_root_address_inst_ack_0, ack => cp_elements(244)); -- 
    -- CP-element group 245 transition  input  output  no-bypass 
    -- predecessors 240 
    -- successors 246 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_671_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_671_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_671_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_670_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_673_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_673_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_673_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_3736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_670_final_reg_ack_0, ack => cp_elements(245)); -- 
    base_resize_req_3753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(245), ack => ptr_deref_674_base_resize_req_0); -- 
    -- CP-element group 246 transition  input  output  no-bypass 
    -- predecessors 245 
    -- successors 247 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_base_resize_ack_0, ack => cp_elements(246)); -- 
    sum_rename_req_3758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_674_root_address_inst_req_0); -- 
    -- CP-element group 247 transition  input  output  no-bypass 
    -- predecessors 246 
    -- successors 248 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_root_address_inst_ack_0, ack => cp_elements(247)); -- 
    root_register_req_3763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => ptr_deref_674_addr_0_req_0); -- 
    -- CP-element group 248 transition  input  output  no-bypass 
    -- predecessors 247 
    -- successors 249 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/word_access_0/rr
      -- 
    root_register_ack_3764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_addr_0_ack_0, ack => cp_elements(248)); -- 
    rr_3774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => ptr_deref_674_load_0_req_0); -- 
    -- CP-element group 249 transition  input  output  no-bypass 
    -- predecessors 248 
    -- successors 250 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/word_access_0/cr
      -- 
    ra_3775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_load_0_ack_0, ack => cp_elements(249)); -- 
    cr_3785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => ptr_deref_674_load_0_req_1); -- 
    -- CP-element group 250 transition  input  output  no-bypass 
    -- predecessors 249 
    -- successors 251 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/merge_req
      -- 
    ca_3786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_load_0_ack_1, ack => cp_elements(250)); -- 
    merge_req_3787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_674_gather_scatter_req_0); -- 
    -- CP-element group 251 transition  input  no-bypass 
    -- predecessors 250 
    -- successors 252 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_675_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_675_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_675_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_674_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_678_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_678_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_678_completed_
      -- 
    merge_ack_3788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_674_gather_scatter_ack_0, ack => cp_elements(251)); -- 
    -- CP-element group 252 join  fork  transition  bypass 
    -- predecessors 230 251 
    -- successors 255 256 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_trigger_
      -- 
    cpelement_group_252 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(230);
      predecessors(1) <= cp_elements(251);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(252)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(252),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 253 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_active_
      -- 
    cp_elements(253) <= cp_elements(41);
    -- CP-element group 254 join  transition  bypass 
    -- predecessors 257 258 
    -- successors 259 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_680_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_680_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_680_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_684_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_684_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_683_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_683_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_683_completed_
      -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(257);
      predecessors(1) <= cp_elements(258);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(254)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 255 transition  output  bypass 
    -- predecessors 252 
    -- successors 257 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Sample/rr
      -- 
    cp_elements(255) <= cp_elements(252);
    rr_3808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => binary_679_inst_req_0); -- 
    -- CP-element group 256 transition  output  bypass 
    -- predecessors 252 
    -- successors 258 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Update/cr
      -- 
    cp_elements(256) <= cp_elements(252);
    cr_3813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => binary_679_inst_req_1); -- 
    -- CP-element group 257 transition  input  no-bypass 
    -- predecessors 255 
    -- successors 254 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Sample/ra
      -- 
    ra_3809_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_679_inst_ack_0, ack => cp_elements(257)); -- 
    -- CP-element group 258 transition  input  no-bypass 
    -- predecessors 256 
    -- successors 254 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_679_Update/ca
      -- 
    ca_3814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_679_inst_ack_1, ack => cp_elements(258)); -- 
    -- CP-element group 259 join  transition  output  bypass 
    -- predecessors 254 263 
    -- successors 264 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/split_req
      -- 
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(254);
      predecessors(1) <= cp_elements(263);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(259)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => ptr_deref_682_gather_scatter_req_0); -- 
    -- CP-element group 260 transition  output  bypass 
    -- predecessors 41 
    -- successors 261 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_681_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_681_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_681_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_addr_resize/base_resize_req
      -- 
    cp_elements(260) <= cp_elements(41);
    base_resize_req_3834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_682_base_resize_req_0); -- 
    -- CP-element group 261 transition  input  output  no-bypass 
    -- predecessors 260 
    -- successors 262 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_base_resize_ack_0, ack => cp_elements(261)); -- 
    sum_rename_req_3839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_682_root_address_inst_req_0); -- 
    -- CP-element group 262 transition  input  output  no-bypass 
    -- predecessors 261 
    -- successors 263 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3840_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_root_address_inst_ack_0, ack => cp_elements(262)); -- 
    root_register_req_3844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(262), ack => ptr_deref_682_addr_0_req_0); -- 
    -- CP-element group 263 transition  input  no-bypass 
    -- predecessors 262 
    -- successors 259 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_word_addrgen/root_register_ack
      -- 
    root_register_ack_3845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_addr_0_ack_0, ack => cp_elements(263)); -- 
    -- CP-element group 264 transition  input  output  no-bypass 
    -- predecessors 259 
    -- successors 265 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/word_access_0/rr
      -- 
    split_ack_3850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_gather_scatter_ack_0, ack => cp_elements(264)); -- 
    rr_3857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_682_store_0_req_0); -- 
    -- CP-element group 265 fork  transition  input  no-bypass 
    -- predecessors 264 
    -- successors 266 688 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_request/word_access/word_access_0/ra
      -- 
    ra_3858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_store_0_ack_0, ack => cp_elements(265)); -- 
    -- CP-element group 266 transition  output  bypass 
    -- predecessors 265 
    -- successors 267 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/word_access_0/cr
      -- 
    cp_elements(266) <= cp_elements(265);
    cr_3868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_682_store_0_req_1); -- 
    -- CP-element group 267 transition  input  no-bypass 
    -- predecessors 266 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_684_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_682_complete/word_access/word_access_0/ca
      -- 
    ca_3869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_682_store_0_ack_1, ack => cp_elements(267)); -- 
    -- CP-element group 268 join  transition  output  bypass 
    -- predecessors 63 272 
    -- successors 273 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/word_access_0/rr
      -- 
    cpelement_group_268 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(63);
      predecessors(1) <= cp_elements(272);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(268)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(268),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_3907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => ptr_deref_687_load_0_req_0); -- 
    -- CP-element group 269 transition  output  bypass 
    -- predecessors 41 
    -- successors 270 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_686_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_686_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_686_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_addr_resize/base_resize_req
      -- 
    cp_elements(269) <= cp_elements(41);
    base_resize_req_3886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_687_base_resize_req_0); -- 
    -- CP-element group 270 transition  input  output  no-bypass 
    -- predecessors 269 
    -- successors 271 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_base_resize_ack_0, ack => cp_elements(270)); -- 
    sum_rename_req_3891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_687_root_address_inst_req_0); -- 
    -- CP-element group 271 transition  input  output  no-bypass 
    -- predecessors 270 
    -- successors 272 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_root_address_inst_ack_0, ack => cp_elements(271)); -- 
    root_register_req_3896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => ptr_deref_687_addr_0_req_0); -- 
    -- CP-element group 272 transition  input  no-bypass 
    -- predecessors 271 
    -- successors 268 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_word_addrgen/root_register_ack
      -- 
    root_register_ack_3897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_addr_0_ack_0, ack => cp_elements(272)); -- 
    -- CP-element group 273 transition  input  output  no-bypass 
    -- predecessors 268 
    -- successors 274 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/word_access_0/cr
      -- 
    ra_3908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_load_0_ack_0, ack => cp_elements(273)); -- 
    cr_3918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_687_load_0_req_1); -- 
    -- CP-element group 274 transition  input  output  no-bypass 
    -- predecessors 273 
    -- successors 275 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/merge_req
      -- 
    ca_3919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_load_0_ack_1, ack => cp_elements(274)); -- 
    merge_req_3920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => ptr_deref_687_gather_scatter_req_0); -- 
    -- CP-element group 275 transition  input  output  no-bypass 
    -- predecessors 274 
    -- successors 276 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_688_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_688_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_688_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_687_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_690_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_690_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_690_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_complete/req
      -- 
    merge_ack_3921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_687_gather_scatter_ack_0, ack => cp_elements(275)); -- 
    req_3934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => type_cast_691_inst_req_0); -- 
    -- CP-element group 276 transition  input  output  no-bypass 
    -- predecessors 275 
    -- successors 279 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_692_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_692_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_692_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_691_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_694_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_694_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_694_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_resize_0/index_resize_req
      -- 
    ack_3935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_691_inst_ack_0, ack => cp_elements(276)); -- 
    index_resize_req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => array_obj_ref_695_index_0_resize_req_0); -- 
    -- CP-element group 277 transition  bypass 
    -- predecessors 41 
    -- successors 278 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_trigger_
      -- 
    cp_elements(277) <= cp_elements(41);
    -- CP-element group 278 join  transition  output  no-bypass 
    -- predecessors 277 282 
    -- successors 283 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_complete/final_reg_req
      -- 
    cpelement_group_278 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(277);
      predecessors(1) <= cp_elements(282);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(278)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(278),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => addr_of_696_final_reg_req_0); -- 
    -- CP-element group 279 transition  input  output  no-bypass 
    -- predecessors 276 
    -- successors 280 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_3954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_695_index_0_resize_ack_0, ack => cp_elements(279)); -- 
    scale_rename_req_3958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => array_obj_ref_695_index_0_rename_req_0); -- 
    -- CP-element group 280 transition  input  output  no-bypass 
    -- predecessors 279 
    -- successors 281 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_add_indices/final_index_req
      -- 
    scale_rename_ack_3959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_695_index_0_rename_ack_0, ack => cp_elements(280)); -- 
    final_index_req_3963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => array_obj_ref_695_offset_inst_req_0); -- 
    -- CP-element group 281 transition  input  output  no-bypass 
    -- predecessors 280 
    -- successors 282 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_3964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_695_offset_inst_ack_0, ack => cp_elements(281)); -- 
    sum_rename_req_3968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => array_obj_ref_695_root_address_inst_req_0); -- 
    -- CP-element group 282 transition  input  no-bypass 
    -- predecessors 281 
    -- successors 278 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_695_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_695_root_address_inst_ack_0, ack => cp_elements(282)); -- 
    -- CP-element group 283 transition  input  output  no-bypass 
    -- predecessors 278 
    -- successors 284 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_697_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_697_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_697_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_696_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_699_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_699_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_699_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_3974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_696_final_reg_ack_0, ack => cp_elements(283)); -- 
    base_resize_req_3991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => ptr_deref_700_base_resize_req_0); -- 
    -- CP-element group 284 transition  input  output  no-bypass 
    -- predecessors 283 
    -- successors 285 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_3992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_base_resize_ack_0, ack => cp_elements(284)); -- 
    sum_rename_req_3996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_700_root_address_inst_req_0); -- 
    -- CP-element group 285 transition  input  output  no-bypass 
    -- predecessors 284 
    -- successors 286 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_word_addrgen/root_register_req
      -- 
    sum_rename_ack_3997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_root_address_inst_ack_0, ack => cp_elements(285)); -- 
    root_register_req_4001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(285), ack => ptr_deref_700_addr_0_req_0); -- 
    -- CP-element group 286 transition  input  output  no-bypass 
    -- predecessors 285 
    -- successors 287 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_addr_0_ack_0, ack => cp_elements(286)); -- 
    rr_4012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_700_load_0_req_0); -- 
    -- CP-element group 287 transition  input  output  no-bypass 
    -- predecessors 286 
    -- successors 288 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/word_access_0/cr
      -- 
    ra_4013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_load_0_ack_0, ack => cp_elements(287)); -- 
    cr_4023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(287), ack => ptr_deref_700_load_0_req_1); -- 
    -- CP-element group 288 transition  input  output  no-bypass 
    -- predecessors 287 
    -- successors 289 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/merge_req
      -- 
    ca_4024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_load_0_ack_1, ack => cp_elements(288)); -- 
    merge_req_4025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_700_gather_scatter_req_0); -- 
    -- CP-element group 289 transition  input  no-bypass 
    -- predecessors 288 
    -- successors 312 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_701_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_701_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_701_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_700_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_720_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_720_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_720_completed_
      -- 
    merge_ack_4026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_700_gather_scatter_ack_0, ack => cp_elements(289)); -- 
    -- CP-element group 290 join  transition  output  bypass 
    -- predecessors 63 294 
    -- successors 295 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/word_access_0/rr
      -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(63);
      predecessors(1) <= cp_elements(294);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(290)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_704_load_0_req_0); -- 
    -- CP-element group 291 transition  output  bypass 
    -- predecessors 41 
    -- successors 292 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_703_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_703_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_703_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_addr_resize/base_resize_req
      -- 
    cp_elements(291) <= cp_elements(41);
    base_resize_req_4043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(291), ack => ptr_deref_704_base_resize_req_0); -- 
    -- CP-element group 292 transition  input  output  no-bypass 
    -- predecessors 291 
    -- successors 293 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_base_resize_ack_0, ack => cp_elements(292)); -- 
    sum_rename_req_4048_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => ptr_deref_704_root_address_inst_req_0); -- 
    -- CP-element group 293 transition  input  output  no-bypass 
    -- predecessors 292 
    -- successors 294 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4049_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_root_address_inst_ack_0, ack => cp_elements(293)); -- 
    root_register_req_4053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => ptr_deref_704_addr_0_req_0); -- 
    -- CP-element group 294 transition  input  no-bypass 
    -- predecessors 293 
    -- successors 290 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_word_addrgen/root_register_ack
      -- 
    root_register_ack_4054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_addr_0_ack_0, ack => cp_elements(294)); -- 
    -- CP-element group 295 transition  input  output  no-bypass 
    -- predecessors 290 
    -- successors 296 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/word_access_0/cr
      -- 
    ra_4065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_load_0_ack_0, ack => cp_elements(295)); -- 
    cr_4075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => ptr_deref_704_load_0_req_1); -- 
    -- CP-element group 296 transition  input  output  no-bypass 
    -- predecessors 295 
    -- successors 297 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/merge_req
      -- 
    ca_4076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_load_0_ack_1, ack => cp_elements(296)); -- 
    merge_req_4077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => ptr_deref_704_gather_scatter_req_0); -- 
    -- CP-element group 297 transition  input  output  no-bypass 
    -- predecessors 296 
    -- successors 298 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_705_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_705_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_705_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_704_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_707_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_707_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_707_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_complete/req
      -- 
    merge_ack_4078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_704_gather_scatter_ack_0, ack => cp_elements(297)); -- 
    req_4091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => type_cast_708_inst_req_0); -- 
    -- CP-element group 298 transition  input  output  no-bypass 
    -- predecessors 297 
    -- successors 301 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_709_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_709_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_709_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_708_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_711_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_711_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_711_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_resize_0/index_resize_req
      -- 
    ack_4092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_708_inst_ack_0, ack => cp_elements(298)); -- 
    index_resize_req_4110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => array_obj_ref_712_index_0_resize_req_0); -- 
    -- CP-element group 299 transition  bypass 
    -- predecessors 41 
    -- successors 300 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_trigger_
      -- 
    cp_elements(299) <= cp_elements(41);
    -- CP-element group 300 join  transition  output  no-bypass 
    -- predecessors 299 304 
    -- successors 305 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_complete/final_reg_req
      -- 
    cpelement_group_300 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(299);
      predecessors(1) <= cp_elements(304);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(300)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(300),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => addr_of_713_final_reg_req_0); -- 
    -- CP-element group 301 transition  input  output  no-bypass 
    -- predecessors 298 
    -- successors 302 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_index_0_resize_ack_0, ack => cp_elements(301)); -- 
    scale_rename_req_4115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => array_obj_ref_712_index_0_rename_req_0); -- 
    -- CP-element group 302 transition  input  output  no-bypass 
    -- predecessors 301 
    -- successors 303 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_add_indices/final_index_req
      -- 
    scale_rename_ack_4116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_index_0_rename_ack_0, ack => cp_elements(302)); -- 
    final_index_req_4120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => array_obj_ref_712_offset_inst_req_0); -- 
    -- CP-element group 303 transition  input  output  no-bypass 
    -- predecessors 302 
    -- successors 304 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_offset_inst_ack_0, ack => cp_elements(303)); -- 
    sum_rename_req_4125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(303), ack => array_obj_ref_712_root_address_inst_req_0); -- 
    -- CP-element group 304 transition  input  no-bypass 
    -- predecessors 303 
    -- successors 300 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_712_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_712_root_address_inst_ack_0, ack => cp_elements(304)); -- 
    -- CP-element group 305 transition  input  output  no-bypass 
    -- predecessors 300 
    -- successors 306 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_714_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_714_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_714_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_713_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_716_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_716_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_716_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_4131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_713_final_reg_ack_0, ack => cp_elements(305)); -- 
    base_resize_req_4148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => ptr_deref_717_base_resize_req_0); -- 
    -- CP-element group 306 transition  input  output  no-bypass 
    -- predecessors 305 
    -- successors 307 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_base_resize_ack_0, ack => cp_elements(306)); -- 
    sum_rename_req_4153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => ptr_deref_717_root_address_inst_req_0); -- 
    -- CP-element group 307 transition  input  output  no-bypass 
    -- predecessors 306 
    -- successors 308 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_root_address_inst_ack_0, ack => cp_elements(307)); -- 
    root_register_req_4158_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(307), ack => ptr_deref_717_addr_0_req_0); -- 
    -- CP-element group 308 transition  input  output  no-bypass 
    -- predecessors 307 
    -- successors 309 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4159_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_addr_0_ack_0, ack => cp_elements(308)); -- 
    rr_4169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => ptr_deref_717_load_0_req_0); -- 
    -- CP-element group 309 transition  input  output  no-bypass 
    -- predecessors 308 
    -- successors 310 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/word_access_0/cr
      -- 
    ra_4170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_load_0_ack_0, ack => cp_elements(309)); -- 
    cr_4180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => ptr_deref_717_load_0_req_1); -- 
    -- CP-element group 310 transition  input  output  no-bypass 
    -- predecessors 309 
    -- successors 311 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/merge_req
      -- 
    ca_4181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_load_0_ack_1, ack => cp_elements(310)); -- 
    merge_req_4182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(310), ack => ptr_deref_717_gather_scatter_req_0); -- 
    -- CP-element group 311 transition  input  no-bypass 
    -- predecessors 310 
    -- successors 312 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_718_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_718_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_718_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_717_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_721_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_721_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_721_completed_
      -- 
    merge_ack_4183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_717_gather_scatter_ack_0, ack => cp_elements(311)); -- 
    -- CP-element group 312 join  fork  transition  bypass 
    -- predecessors 289 311 
    -- successors 315 316 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_trigger_
      -- 
    cpelement_group_312 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(289);
      predecessors(1) <= cp_elements(311);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(312)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(312),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 313 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_active_
      -- 
    cp_elements(313) <= cp_elements(41);
    -- CP-element group 314 join  transition  bypass 
    -- predecessors 317 318 
    -- successors 319 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_723_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_723_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_723_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_727_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_727_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_726_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_726_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_726_completed_
      -- 
    cpelement_group_314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(317);
      predecessors(1) <= cp_elements(318);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(314)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 315 transition  output  bypass 
    -- predecessors 312 
    -- successors 317 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Sample/rr
      -- 
    cp_elements(315) <= cp_elements(312);
    rr_4203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => binary_722_inst_req_0); -- 
    -- CP-element group 316 transition  output  bypass 
    -- predecessors 312 
    -- successors 318 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Update/cr
      -- 
    cp_elements(316) <= cp_elements(312);
    cr_4208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(316), ack => binary_722_inst_req_1); -- 
    -- CP-element group 317 transition  input  no-bypass 
    -- predecessors 315 
    -- successors 314 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Sample/ra
      -- 
    ra_4204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_722_inst_ack_0, ack => cp_elements(317)); -- 
    -- CP-element group 318 transition  input  no-bypass 
    -- predecessors 316 
    -- successors 314 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_722_Update/ca
      -- 
    ca_4209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_722_inst_ack_1, ack => cp_elements(318)); -- 
    -- CP-element group 319 join  transition  output  bypass 
    -- predecessors 314 323 
    -- successors 324 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/split_req
      -- 
    cpelement_group_319 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(314);
      predecessors(1) <= cp_elements(323);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(319)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(319),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_4244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => ptr_deref_725_gather_scatter_req_0); -- 
    -- CP-element group 320 transition  output  bypass 
    -- predecessors 41 
    -- successors 321 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_724_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_724_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_724_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_addr_resize/base_resize_req
      -- 
    cp_elements(320) <= cp_elements(41);
    base_resize_req_4229_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(320), ack => ptr_deref_725_base_resize_req_0); -- 
    -- CP-element group 321 transition  input  output  no-bypass 
    -- predecessors 320 
    -- successors 322 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4230_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_base_resize_ack_0, ack => cp_elements(321)); -- 
    sum_rename_req_4234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => ptr_deref_725_root_address_inst_req_0); -- 
    -- CP-element group 322 transition  input  output  no-bypass 
    -- predecessors 321 
    -- successors 323 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_root_address_inst_ack_0, ack => cp_elements(322)); -- 
    root_register_req_4239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => ptr_deref_725_addr_0_req_0); -- 
    -- CP-element group 323 transition  input  no-bypass 
    -- predecessors 322 
    -- successors 319 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_word_addrgen/root_register_ack
      -- 
    root_register_ack_4240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_addr_0_ack_0, ack => cp_elements(323)); -- 
    -- CP-element group 324 transition  input  output  no-bypass 
    -- predecessors 319 
    -- successors 325 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/word_access_0/rr
      -- 
    split_ack_4245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_gather_scatter_ack_0, ack => cp_elements(324)); -- 
    rr_4252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(324), ack => ptr_deref_725_store_0_req_0); -- 
    -- CP-element group 325 fork  transition  input  no-bypass 
    -- predecessors 324 
    -- successors 326 719 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_request/word_access/word_access_0/ra
      -- 
    ra_4253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_store_0_ack_0, ack => cp_elements(325)); -- 
    -- CP-element group 326 transition  output  bypass 
    -- predecessors 325 
    -- successors 327 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/word_access_0/cr
      -- 
    cp_elements(326) <= cp_elements(325);
    cr_4263_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => ptr_deref_725_store_0_req_1); -- 
    -- CP-element group 327 transition  input  no-bypass 
    -- predecessors 326 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_727_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_725_complete/word_access/word_access_0/ca
      -- 
    ca_4264_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_725_store_0_ack_1, ack => cp_elements(327)); -- 
    -- CP-element group 328 join  transition  output  bypass 
    -- predecessors 87 332 
    -- successors 333 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/word_access_0/rr
      -- 
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(87);
      predecessors(1) <= cp_elements(332);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(328)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => ptr_deref_730_load_0_req_0); -- 
    -- CP-element group 329 transition  output  bypass 
    -- predecessors 41 
    -- successors 330 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_729_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_729_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_729_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_addr_resize/base_resize_req
      -- 
    cp_elements(329) <= cp_elements(41);
    base_resize_req_4281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => ptr_deref_730_base_resize_req_0); -- 
    -- CP-element group 330 transition  input  output  no-bypass 
    -- predecessors 329 
    -- successors 331 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_base_resize_ack_0, ack => cp_elements(330)); -- 
    sum_rename_req_4286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => ptr_deref_730_root_address_inst_req_0); -- 
    -- CP-element group 331 transition  input  output  no-bypass 
    -- predecessors 330 
    -- successors 332 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_root_address_inst_ack_0, ack => cp_elements(331)); -- 
    root_register_req_4291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => ptr_deref_730_addr_0_req_0); -- 
    -- CP-element group 332 transition  input  no-bypass 
    -- predecessors 331 
    -- successors 328 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_word_addrgen/root_register_ack
      -- 
    root_register_ack_4292_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_addr_0_ack_0, ack => cp_elements(332)); -- 
    -- CP-element group 333 transition  input  output  no-bypass 
    -- predecessors 328 
    -- successors 334 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/word_access_0/cr
      -- 
    ra_4303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_load_0_ack_0, ack => cp_elements(333)); -- 
    cr_4313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => ptr_deref_730_load_0_req_1); -- 
    -- CP-element group 334 transition  input  output  no-bypass 
    -- predecessors 333 
    -- successors 335 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/merge_req
      -- 
    ca_4314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_load_0_ack_1, ack => cp_elements(334)); -- 
    merge_req_4315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(334), ack => ptr_deref_730_gather_scatter_req_0); -- 
    -- CP-element group 335 transition  input  output  no-bypass 
    -- predecessors 334 
    -- successors 336 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_731_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_731_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_731_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_730_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_733_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_733_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_733_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_complete/req
      -- 
    merge_ack_4316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_730_gather_scatter_ack_0, ack => cp_elements(335)); -- 
    req_4329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => type_cast_734_inst_req_0); -- 
    -- CP-element group 336 transition  input  output  no-bypass 
    -- predecessors 335 
    -- successors 339 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_735_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_735_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_735_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_734_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_737_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_737_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_737_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_resize_0/index_resize_req
      -- 
    ack_4330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_734_inst_ack_0, ack => cp_elements(336)); -- 
    index_resize_req_4348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => array_obj_ref_738_index_0_resize_req_0); -- 
    -- CP-element group 337 transition  bypass 
    -- predecessors 41 
    -- successors 338 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_trigger_
      -- 
    cp_elements(337) <= cp_elements(41);
    -- CP-element group 338 join  transition  output  no-bypass 
    -- predecessors 337 342 
    -- successors 343 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_complete/final_reg_req
      -- 
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(337);
      predecessors(1) <= cp_elements(342);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(338)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => addr_of_739_final_reg_req_0); -- 
    -- CP-element group 339 transition  input  output  no-bypass 
    -- predecessors 336 
    -- successors 340 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_index_0_resize_ack_0, ack => cp_elements(339)); -- 
    scale_rename_req_4353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => array_obj_ref_738_index_0_rename_req_0); -- 
    -- CP-element group 340 transition  input  output  no-bypass 
    -- predecessors 339 
    -- successors 341 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_add_indices/final_index_req
      -- 
    scale_rename_ack_4354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_index_0_rename_ack_0, ack => cp_elements(340)); -- 
    final_index_req_4358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => array_obj_ref_738_offset_inst_req_0); -- 
    -- CP-element group 341 transition  input  output  no-bypass 
    -- predecessors 340 
    -- successors 342 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_offset_inst_ack_0, ack => cp_elements(341)); -- 
    sum_rename_req_4363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => array_obj_ref_738_root_address_inst_req_0); -- 
    -- CP-element group 342 transition  input  no-bypass 
    -- predecessors 341 
    -- successors 338 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_738_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_738_root_address_inst_ack_0, ack => cp_elements(342)); -- 
    -- CP-element group 343 transition  input  output  no-bypass 
    -- predecessors 338 
    -- successors 344 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_740_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_740_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_740_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_739_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_742_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_742_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_742_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_4369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_739_final_reg_ack_0, ack => cp_elements(343)); -- 
    base_resize_req_4386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(343), ack => ptr_deref_743_base_resize_req_0); -- 
    -- CP-element group 344 transition  input  output  no-bypass 
    -- predecessors 343 
    -- successors 345 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_base_resize_ack_0, ack => cp_elements(344)); -- 
    sum_rename_req_4391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(344), ack => ptr_deref_743_root_address_inst_req_0); -- 
    -- CP-element group 345 transition  input  output  no-bypass 
    -- predecessors 344 
    -- successors 346 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_root_address_inst_ack_0, ack => cp_elements(345)); -- 
    root_register_req_4396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => ptr_deref_743_addr_0_req_0); -- 
    -- CP-element group 346 transition  input  output  no-bypass 
    -- predecessors 345 
    -- successors 347 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_addr_0_ack_0, ack => cp_elements(346)); -- 
    rr_4407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(346), ack => ptr_deref_743_load_0_req_0); -- 
    -- CP-element group 347 transition  input  output  no-bypass 
    -- predecessors 346 
    -- successors 348 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/word_access_0/cr
      -- 
    ra_4408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_load_0_ack_0, ack => cp_elements(347)); -- 
    cr_4418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(347), ack => ptr_deref_743_load_0_req_1); -- 
    -- CP-element group 348 transition  input  output  no-bypass 
    -- predecessors 347 
    -- successors 349 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/merge_req
      -- 
    ca_4419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_load_0_ack_1, ack => cp_elements(348)); -- 
    merge_req_4420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => ptr_deref_743_gather_scatter_req_0); -- 
    -- CP-element group 349 transition  input  no-bypass 
    -- predecessors 348 
    -- successors 372 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_744_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_744_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_744_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_743_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_763_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_763_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_763_completed_
      -- 
    merge_ack_4421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_743_gather_scatter_ack_0, ack => cp_elements(349)); -- 
    -- CP-element group 350 join  transition  output  bypass 
    -- predecessors 87 354 
    -- successors 355 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/word_access_0/rr
      -- 
    cpelement_group_350 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(87);
      predecessors(1) <= cp_elements(354);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(350)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(350),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => ptr_deref_747_load_0_req_0); -- 
    -- CP-element group 351 transition  output  bypass 
    -- predecessors 41 
    -- successors 352 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_746_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_746_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_746_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_addr_resize/base_resize_req
      -- 
    cp_elements(351) <= cp_elements(41);
    base_resize_req_4438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => ptr_deref_747_base_resize_req_0); -- 
    -- CP-element group 352 transition  input  output  no-bypass 
    -- predecessors 351 
    -- successors 353 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_base_resize_ack_0, ack => cp_elements(352)); -- 
    sum_rename_req_4443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(352), ack => ptr_deref_747_root_address_inst_req_0); -- 
    -- CP-element group 353 transition  input  output  no-bypass 
    -- predecessors 352 
    -- successors 354 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_root_address_inst_ack_0, ack => cp_elements(353)); -- 
    root_register_req_4448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => ptr_deref_747_addr_0_req_0); -- 
    -- CP-element group 354 transition  input  no-bypass 
    -- predecessors 353 
    -- successors 350 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_word_addrgen/root_register_ack
      -- 
    root_register_ack_4449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_addr_0_ack_0, ack => cp_elements(354)); -- 
    -- CP-element group 355 transition  input  output  no-bypass 
    -- predecessors 350 
    -- successors 356 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/word_access_0/cr
      -- 
    ra_4460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_load_0_ack_0, ack => cp_elements(355)); -- 
    cr_4470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(355), ack => ptr_deref_747_load_0_req_1); -- 
    -- CP-element group 356 transition  input  output  no-bypass 
    -- predecessors 355 
    -- successors 357 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/merge_req
      -- 
    ca_4471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_load_0_ack_1, ack => cp_elements(356)); -- 
    merge_req_4472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => ptr_deref_747_gather_scatter_req_0); -- 
    -- CP-element group 357 transition  input  output  no-bypass 
    -- predecessors 356 
    -- successors 358 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_748_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_748_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_748_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_747_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_750_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_750_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_750_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_complete/req
      -- 
    merge_ack_4473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_747_gather_scatter_ack_0, ack => cp_elements(357)); -- 
    req_4486_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => type_cast_751_inst_req_0); -- 
    -- CP-element group 358 transition  input  output  no-bypass 
    -- predecessors 357 
    -- successors 361 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_752_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_752_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_752_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_751_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_754_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_754_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_754_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_resize_0/index_resize_req
      -- 
    ack_4487_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_751_inst_ack_0, ack => cp_elements(358)); -- 
    index_resize_req_4505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => array_obj_ref_755_index_0_resize_req_0); -- 
    -- CP-element group 359 transition  bypass 
    -- predecessors 41 
    -- successors 360 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_trigger_
      -- 
    cp_elements(359) <= cp_elements(41);
    -- CP-element group 360 join  transition  output  no-bypass 
    -- predecessors 359 364 
    -- successors 365 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_complete/final_reg_req
      -- 
    cpelement_group_360 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(359);
      predecessors(1) <= cp_elements(364);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(360)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(360),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => addr_of_756_final_reg_req_0); -- 
    -- CP-element group 361 transition  input  output  no-bypass 
    -- predecessors 358 
    -- successors 362 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_755_index_0_resize_ack_0, ack => cp_elements(361)); -- 
    scale_rename_req_4510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(361), ack => array_obj_ref_755_index_0_rename_req_0); -- 
    -- CP-element group 362 transition  input  output  no-bypass 
    -- predecessors 361 
    -- successors 363 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_add_indices/final_index_req
      -- 
    scale_rename_ack_4511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_755_index_0_rename_ack_0, ack => cp_elements(362)); -- 
    final_index_req_4515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => array_obj_ref_755_offset_inst_req_0); -- 
    -- CP-element group 363 transition  input  output  no-bypass 
    -- predecessors 362 
    -- successors 364 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_755_offset_inst_ack_0, ack => cp_elements(363)); -- 
    sum_rename_req_4520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(363), ack => array_obj_ref_755_root_address_inst_req_0); -- 
    -- CP-element group 364 transition  input  no-bypass 
    -- predecessors 363 
    -- successors 360 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_755_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_755_root_address_inst_ack_0, ack => cp_elements(364)); -- 
    -- CP-element group 365 transition  input  output  no-bypass 
    -- predecessors 360 
    -- successors 366 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_757_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_757_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_757_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_756_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_759_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_759_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_759_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_4526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_756_final_reg_ack_0, ack => cp_elements(365)); -- 
    base_resize_req_4543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(365), ack => ptr_deref_760_base_resize_req_0); -- 
    -- CP-element group 366 transition  input  output  no-bypass 
    -- predecessors 365 
    -- successors 367 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_base_resize_ack_0, ack => cp_elements(366)); -- 
    sum_rename_req_4548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(366), ack => ptr_deref_760_root_address_inst_req_0); -- 
    -- CP-element group 367 transition  input  output  no-bypass 
    -- predecessors 366 
    -- successors 368 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_root_address_inst_ack_0, ack => cp_elements(367)); -- 
    root_register_req_4553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(367), ack => ptr_deref_760_addr_0_req_0); -- 
    -- CP-element group 368 transition  input  output  no-bypass 
    -- predecessors 367 
    -- successors 369 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_addr_0_ack_0, ack => cp_elements(368)); -- 
    rr_4564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(368), ack => ptr_deref_760_load_0_req_0); -- 
    -- CP-element group 369 transition  input  output  no-bypass 
    -- predecessors 368 
    -- successors 370 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/word_access_0/cr
      -- 
    ra_4565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_load_0_ack_0, ack => cp_elements(369)); -- 
    cr_4575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(369), ack => ptr_deref_760_load_0_req_1); -- 
    -- CP-element group 370 transition  input  output  no-bypass 
    -- predecessors 369 
    -- successors 371 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/merge_req
      -- 
    ca_4576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_load_0_ack_1, ack => cp_elements(370)); -- 
    merge_req_4577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(370), ack => ptr_deref_760_gather_scatter_req_0); -- 
    -- CP-element group 371 transition  input  no-bypass 
    -- predecessors 370 
    -- successors 372 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_761_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_761_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_761_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_760_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_764_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_764_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_764_completed_
      -- 
    merge_ack_4578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_760_gather_scatter_ack_0, ack => cp_elements(371)); -- 
    -- CP-element group 372 join  fork  transition  bypass 
    -- predecessors 349 371 
    -- successors 375 376 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_trigger_
      -- 
    cpelement_group_372 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(349);
      predecessors(1) <= cp_elements(371);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(372)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(372),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 373 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_active_
      -- 
    cp_elements(373) <= cp_elements(41);
    -- CP-element group 374 join  transition  bypass 
    -- predecessors 377 378 
    -- successors 379 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_766_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_766_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_766_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_770_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_770_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_769_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_769_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_769_completed_
      -- 
    cpelement_group_374 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(377);
      predecessors(1) <= cp_elements(378);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(374)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 375 transition  output  bypass 
    -- predecessors 372 
    -- successors 377 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Sample/rr
      -- 
    cp_elements(375) <= cp_elements(372);
    rr_4598_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(375), ack => binary_765_inst_req_0); -- 
    -- CP-element group 376 transition  output  bypass 
    -- predecessors 372 
    -- successors 378 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Update/cr
      -- 
    cp_elements(376) <= cp_elements(372);
    cr_4603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(376), ack => binary_765_inst_req_1); -- 
    -- CP-element group 377 transition  input  no-bypass 
    -- predecessors 375 
    -- successors 374 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Sample/ra
      -- 
    ra_4599_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_765_inst_ack_0, ack => cp_elements(377)); -- 
    -- CP-element group 378 transition  input  no-bypass 
    -- predecessors 376 
    -- successors 374 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_765_Update/ca
      -- 
    ca_4604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_765_inst_ack_1, ack => cp_elements(378)); -- 
    -- CP-element group 379 join  transition  output  bypass 
    -- predecessors 374 383 
    -- successors 384 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/split_req
      -- 
    cpelement_group_379 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(374);
      predecessors(1) <= cp_elements(383);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(379)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(379),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_4639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => ptr_deref_768_gather_scatter_req_0); -- 
    -- CP-element group 380 transition  output  bypass 
    -- predecessors 41 
    -- successors 381 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_767_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_767_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_767_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_addr_resize/base_resize_req
      -- 
    cp_elements(380) <= cp_elements(41);
    base_resize_req_4624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => ptr_deref_768_base_resize_req_0); -- 
    -- CP-element group 381 transition  input  output  no-bypass 
    -- predecessors 380 
    -- successors 382 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_base_resize_ack_0, ack => cp_elements(381)); -- 
    sum_rename_req_4629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => ptr_deref_768_root_address_inst_req_0); -- 
    -- CP-element group 382 transition  input  output  no-bypass 
    -- predecessors 381 
    -- successors 383 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_root_address_inst_ack_0, ack => cp_elements(382)); -- 
    root_register_req_4634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(382), ack => ptr_deref_768_addr_0_req_0); -- 
    -- CP-element group 383 transition  input  no-bypass 
    -- predecessors 382 
    -- successors 379 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_word_addrgen/root_register_ack
      -- 
    root_register_ack_4635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_addr_0_ack_0, ack => cp_elements(383)); -- 
    -- CP-element group 384 transition  input  output  no-bypass 
    -- predecessors 379 
    -- successors 385 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/word_access_0/rr
      -- 
    split_ack_4640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_gather_scatter_ack_0, ack => cp_elements(384)); -- 
    rr_4647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => ptr_deref_768_store_0_req_0); -- 
    -- CP-element group 385 fork  transition  input  no-bypass 
    -- predecessors 384 
    -- successors 386 751 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_request/word_access/word_access_0/ra
      -- 
    ra_4648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_store_0_ack_0, ack => cp_elements(385)); -- 
    -- CP-element group 386 transition  output  bypass 
    -- predecessors 385 
    -- successors 387 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/word_access_0/cr
      -- 
    cp_elements(386) <= cp_elements(385);
    cr_4658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => ptr_deref_768_store_0_req_1); -- 
    -- CP-element group 387 transition  input  no-bypass 
    -- predecessors 386 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_770_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_768_complete/word_access/word_access_0/ca
      -- 
    ca_4659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_768_store_0_ack_1, ack => cp_elements(387)); -- 
    -- CP-element group 388 join  transition  output  bypass 
    -- predecessors 111 392 
    -- successors 393 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/word_access_0/rr
      -- 
    cpelement_group_388 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(111);
      predecessors(1) <= cp_elements(392);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(388)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(388),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(388), ack => ptr_deref_773_load_0_req_0); -- 
    -- CP-element group 389 transition  output  bypass 
    -- predecessors 41 
    -- successors 390 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_772_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_772_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_772_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_addr_resize/base_resize_req
      -- 
    cp_elements(389) <= cp_elements(41);
    base_resize_req_4676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(389), ack => ptr_deref_773_base_resize_req_0); -- 
    -- CP-element group 390 transition  input  output  no-bypass 
    -- predecessors 389 
    -- successors 391 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_base_resize_ack_0, ack => cp_elements(390)); -- 
    sum_rename_req_4681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(390), ack => ptr_deref_773_root_address_inst_req_0); -- 
    -- CP-element group 391 transition  input  output  no-bypass 
    -- predecessors 390 
    -- successors 392 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4682_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_root_address_inst_ack_0, ack => cp_elements(391)); -- 
    root_register_req_4686_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(391), ack => ptr_deref_773_addr_0_req_0); -- 
    -- CP-element group 392 transition  input  no-bypass 
    -- predecessors 391 
    -- successors 388 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_word_addrgen/root_register_ack
      -- 
    root_register_ack_4687_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_addr_0_ack_0, ack => cp_elements(392)); -- 
    -- CP-element group 393 transition  input  output  no-bypass 
    -- predecessors 388 
    -- successors 394 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/$entry
      -- 
    ra_4698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_load_0_ack_0, ack => cp_elements(393)); -- 
    cr_4708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(393), ack => ptr_deref_773_load_0_req_1); -- 
    -- CP-element group 394 transition  input  output  no-bypass 
    -- predecessors 393 
    -- successors 395 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/merge_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/word_access/$exit
      -- 
    ca_4709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_load_0_ack_1, ack => cp_elements(394)); -- 
    merge_req_4710_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => ptr_deref_773_gather_scatter_req_0); -- 
    -- CP-element group 395 transition  input  output  no-bypass 
    -- predecessors 394 
    -- successors 396 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_774_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_774_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_774_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_773_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_776_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_776_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_776_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_complete/req
      -- 
    merge_ack_4711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_773_gather_scatter_ack_0, ack => cp_elements(395)); -- 
    req_4724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(395), ack => type_cast_777_inst_req_0); -- 
    -- CP-element group 396 transition  input  output  no-bypass 
    -- predecessors 395 
    -- successors 399 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_780_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_780_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_780_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_778_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_778_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_resize_0/index_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_778_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_777_complete/ack
      -- 
    ack_4725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_777_inst_ack_0, ack => cp_elements(396)); -- 
    index_resize_req_4743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(396), ack => array_obj_ref_781_index_0_resize_req_0); -- 
    -- CP-element group 397 transition  bypass 
    -- predecessors 41 
    -- successors 398 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_trigger_
      -- 
    cp_elements(397) <= cp_elements(41);
    -- CP-element group 398 join  transition  output  no-bypass 
    -- predecessors 397 402 
    -- successors 403 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_complete/final_reg_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_complete/$entry
      -- 
    cpelement_group_398 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(397);
      predecessors(1) <= cp_elements(402);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(398)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(398),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(398), ack => addr_of_782_final_reg_req_0); -- 
    -- CP-element group 399 transition  input  output  no-bypass 
    -- predecessors 396 
    -- successors 400 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_index_0_resize_ack_0, ack => cp_elements(399)); -- 
    scale_rename_req_4748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(399), ack => array_obj_ref_781_index_0_rename_req_0); -- 
    -- CP-element group 400 transition  input  output  no-bypass 
    -- predecessors 399 
    -- successors 401 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_add_indices/final_index_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_4749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_index_0_rename_ack_0, ack => cp_elements(400)); -- 
    final_index_req_4753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => array_obj_ref_781_offset_inst_req_0); -- 
    -- CP-element group 401 transition  input  output  no-bypass 
    -- predecessors 400 
    -- successors 402 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_base_plus_offset/$entry
      -- 
    final_index_ack_4754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_offset_inst_ack_0, ack => cp_elements(401)); -- 
    sum_rename_req_4758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(401), ack => array_obj_ref_781_root_address_inst_req_0); -- 
    -- CP-element group 402 transition  input  no-bypass 
    -- predecessors 401 
    -- successors 398 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_781_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_781_root_address_inst_ack_0, ack => cp_elements(402)); -- 
    -- CP-element group 403 transition  input  output  no-bypass 
    -- predecessors 398 
    -- successors 404 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_782_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_785_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_783_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_785_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_783_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_785_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_783_active_
      -- 
    final_reg_ack_4764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_782_final_reg_ack_0, ack => cp_elements(403)); -- 
    base_resize_req_4781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(403), ack => ptr_deref_786_base_resize_req_0); -- 
    -- CP-element group 404 transition  input  output  no-bypass 
    -- predecessors 403 
    -- successors 405 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_4782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_base_resize_ack_0, ack => cp_elements(404)); -- 
    sum_rename_req_4786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(404), ack => ptr_deref_786_root_address_inst_req_0); -- 
    -- CP-element group 405 transition  input  output  no-bypass 
    -- predecessors 404 
    -- successors 406 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_root_address_inst_ack_0, ack => cp_elements(405)); -- 
    root_register_req_4791_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(405), ack => ptr_deref_786_addr_0_req_0); -- 
    -- CP-element group 406 transition  input  output  no-bypass 
    -- predecessors 405 
    -- successors 407 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4792_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_addr_0_ack_0, ack => cp_elements(406)); -- 
    rr_4802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => ptr_deref_786_load_0_req_0); -- 
    -- CP-element group 407 transition  input  output  no-bypass 
    -- predecessors 406 
    -- successors 408 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/word_access_0/cr
      -- 
    ra_4803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_load_0_ack_0, ack => cp_elements(407)); -- 
    cr_4813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(407), ack => ptr_deref_786_load_0_req_1); -- 
    -- CP-element group 408 transition  input  output  no-bypass 
    -- predecessors 407 
    -- successors 409 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/merge_req
      -- 
    ca_4814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_load_0_ack_1, ack => cp_elements(408)); -- 
    merge_req_4815_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(408), ack => ptr_deref_786_gather_scatter_req_0); -- 
    -- CP-element group 409 transition  input  no-bypass 
    -- predecessors 408 
    -- successors 432 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_787_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_787_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_787_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_786_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_806_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_806_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_806_completed_
      -- 
    merge_ack_4816_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_786_gather_scatter_ack_0, ack => cp_elements(409)); -- 
    -- CP-element group 410 join  transition  output  bypass 
    -- predecessors 111 414 
    -- successors 415 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/word_access_0/rr
      -- 
    cpelement_group_410 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(111);
      predecessors(1) <= cp_elements(414);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(410)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(410),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(410), ack => ptr_deref_790_load_0_req_0); -- 
    -- CP-element group 411 transition  output  bypass 
    -- predecessors 41 
    -- successors 412 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_789_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_789_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_789_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_addr_resize/base_resize_req
      -- 
    cp_elements(411) <= cp_elements(41);
    base_resize_req_4833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => ptr_deref_790_base_resize_req_0); -- 
    -- CP-element group 412 transition  input  output  no-bypass 
    -- predecessors 411 
    -- successors 413 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4834_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_base_resize_ack_0, ack => cp_elements(412)); -- 
    sum_rename_req_4838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(412), ack => ptr_deref_790_root_address_inst_req_0); -- 
    -- CP-element group 413 transition  input  output  no-bypass 
    -- predecessors 412 
    -- successors 414 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_root_address_inst_ack_0, ack => cp_elements(413)); -- 
    root_register_req_4843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(413), ack => ptr_deref_790_addr_0_req_0); -- 
    -- CP-element group 414 transition  input  no-bypass 
    -- predecessors 413 
    -- successors 410 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_word_addrgen/root_register_ack
      -- 
    root_register_ack_4844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_addr_0_ack_0, ack => cp_elements(414)); -- 
    -- CP-element group 415 transition  input  output  no-bypass 
    -- predecessors 410 
    -- successors 416 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/word_access_0/cr
      -- 
    ra_4855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_load_0_ack_0, ack => cp_elements(415)); -- 
    cr_4865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(415), ack => ptr_deref_790_load_0_req_1); -- 
    -- CP-element group 416 transition  input  output  no-bypass 
    -- predecessors 415 
    -- successors 417 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/merge_req
      -- 
    ca_4866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_load_0_ack_1, ack => cp_elements(416)); -- 
    merge_req_4867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(416), ack => ptr_deref_790_gather_scatter_req_0); -- 
    -- CP-element group 417 transition  input  output  no-bypass 
    -- predecessors 416 
    -- successors 418 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_791_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_791_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_791_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_790_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_793_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_793_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_793_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_complete/req
      -- 
    merge_ack_4868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_790_gather_scatter_ack_0, ack => cp_elements(417)); -- 
    req_4881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(417), ack => type_cast_794_inst_req_0); -- 
    -- CP-element group 418 transition  input  output  no-bypass 
    -- predecessors 417 
    -- successors 421 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_795_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_795_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_795_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_794_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_797_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_797_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_797_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_resize_0/index_resize_req
      -- 
    ack_4882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_794_inst_ack_0, ack => cp_elements(418)); -- 
    index_resize_req_4900_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(418), ack => array_obj_ref_798_index_0_resize_req_0); -- 
    -- CP-element group 419 transition  bypass 
    -- predecessors 41 
    -- successors 420 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_trigger_
      -- 
    cp_elements(419) <= cp_elements(41);
    -- CP-element group 420 join  transition  output  no-bypass 
    -- predecessors 419 424 
    -- successors 425 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_complete/final_reg_req
      -- 
    cpelement_group_420 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(419);
      predecessors(1) <= cp_elements(424);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(420)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(420),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(420), ack => addr_of_799_final_reg_req_0); -- 
    -- CP-element group 421 transition  input  output  no-bypass 
    -- predecessors 418 
    -- successors 422 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4901_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_index_0_resize_ack_0, ack => cp_elements(421)); -- 
    scale_rename_req_4905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(421), ack => array_obj_ref_798_index_0_rename_req_0); -- 
    -- CP-element group 422 transition  input  output  no-bypass 
    -- predecessors 421 
    -- successors 423 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_add_indices/final_index_req
      -- 
    scale_rename_ack_4906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_index_0_rename_ack_0, ack => cp_elements(422)); -- 
    final_index_req_4910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(422), ack => array_obj_ref_798_offset_inst_req_0); -- 
    -- CP-element group 423 transition  input  output  no-bypass 
    -- predecessors 422 
    -- successors 424 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_offset_inst_ack_0, ack => cp_elements(423)); -- 
    sum_rename_req_4915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(423), ack => array_obj_ref_798_root_address_inst_req_0); -- 
    -- CP-element group 424 transition  input  no-bypass 
    -- predecessors 423 
    -- successors 420 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_798_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_798_root_address_inst_ack_0, ack => cp_elements(424)); -- 
    -- CP-element group 425 transition  input  output  no-bypass 
    -- predecessors 420 
    -- successors 426 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_800_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_800_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_800_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_799_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_802_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_802_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_802_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_4921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_799_final_reg_ack_0, ack => cp_elements(425)); -- 
    base_resize_req_4938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(425), ack => ptr_deref_803_base_resize_req_0); -- 
    -- CP-element group 426 transition  input  output  no-bypass 
    -- predecessors 425 
    -- successors 427 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_base_resize_ack_0, ack => cp_elements(426)); -- 
    sum_rename_req_4943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(426), ack => ptr_deref_803_root_address_inst_req_0); -- 
    -- CP-element group 427 transition  input  output  no-bypass 
    -- predecessors 426 
    -- successors 428 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_root_address_inst_ack_0, ack => cp_elements(427)); -- 
    root_register_req_4948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(427), ack => ptr_deref_803_addr_0_req_0); -- 
    -- CP-element group 428 transition  input  output  no-bypass 
    -- predecessors 427 
    -- successors 429 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/word_access_0/rr
      -- 
    root_register_ack_4949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_addr_0_ack_0, ack => cp_elements(428)); -- 
    rr_4959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(428), ack => ptr_deref_803_load_0_req_0); -- 
    -- CP-element group 429 transition  input  output  no-bypass 
    -- predecessors 428 
    -- successors 430 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/word_access_0/cr
      -- 
    ra_4960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_0_ack_0, ack => cp_elements(429)); -- 
    cr_4970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(429), ack => ptr_deref_803_load_0_req_1); -- 
    -- CP-element group 430 transition  input  output  no-bypass 
    -- predecessors 429 
    -- successors 431 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/merge_req
      -- 
    ca_4971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_0_ack_1, ack => cp_elements(430)); -- 
    merge_req_4972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(430), ack => ptr_deref_803_gather_scatter_req_0); -- 
    -- CP-element group 431 transition  input  no-bypass 
    -- predecessors 430 
    -- successors 432 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_804_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_804_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_804_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_803_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_807_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_807_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_807_completed_
      -- 
    merge_ack_4973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_gather_scatter_ack_0, ack => cp_elements(431)); -- 
    -- CP-element group 432 join  fork  transition  bypass 
    -- predecessors 409 431 
    -- successors 435 436 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_trigger_
      -- 
    cpelement_group_432 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(409);
      predecessors(1) <= cp_elements(431);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(432)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(432),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 433 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_active_
      -- 
    cp_elements(433) <= cp_elements(41);
    -- CP-element group 434 join  transition  bypass 
    -- predecessors 437 438 
    -- successors 439 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_809_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_809_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_809_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_813_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_813_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_812_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_812_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_812_completed_
      -- 
    cpelement_group_434 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(437);
      predecessors(1) <= cp_elements(438);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(434)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(434),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 435 transition  output  bypass 
    -- predecessors 432 
    -- successors 437 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Sample/rr
      -- 
    cp_elements(435) <= cp_elements(432);
    rr_4993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => binary_808_inst_req_0); -- 
    -- CP-element group 436 transition  output  bypass 
    -- predecessors 432 
    -- successors 438 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Update/cr
      -- 
    cp_elements(436) <= cp_elements(432);
    cr_4998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => binary_808_inst_req_1); -- 
    -- CP-element group 437 transition  input  no-bypass 
    -- predecessors 435 
    -- successors 434 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Sample/ra
      -- 
    ra_4994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_808_inst_ack_0, ack => cp_elements(437)); -- 
    -- CP-element group 438 transition  input  no-bypass 
    -- predecessors 436 
    -- successors 434 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_808_Update/ca
      -- 
    ca_4999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_808_inst_ack_1, ack => cp_elements(438)); -- 
    -- CP-element group 439 join  transition  output  bypass 
    -- predecessors 434 443 
    -- successors 444 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/split_req
      -- 
    cpelement_group_439 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(434);
      predecessors(1) <= cp_elements(443);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(439)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(439),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(439), ack => ptr_deref_811_gather_scatter_req_0); -- 
    -- CP-element group 440 transition  output  bypass 
    -- predecessors 41 
    -- successors 441 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_810_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_810_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_810_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_addr_resize/base_resize_req
      -- 
    cp_elements(440) <= cp_elements(41);
    base_resize_req_5019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(440), ack => ptr_deref_811_base_resize_req_0); -- 
    -- CP-element group 441 transition  input  output  no-bypass 
    -- predecessors 440 
    -- successors 442 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_base_resize_ack_0, ack => cp_elements(441)); -- 
    sum_rename_req_5024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => ptr_deref_811_root_address_inst_req_0); -- 
    -- CP-element group 442 transition  input  output  no-bypass 
    -- predecessors 441 
    -- successors 443 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_root_address_inst_ack_0, ack => cp_elements(442)); -- 
    root_register_req_5029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => ptr_deref_811_addr_0_req_0); -- 
    -- CP-element group 443 transition  input  no-bypass 
    -- predecessors 442 
    -- successors 439 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_word_addrgen/root_register_ack
      -- 
    root_register_ack_5030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_addr_0_ack_0, ack => cp_elements(443)); -- 
    -- CP-element group 444 transition  input  output  no-bypass 
    -- predecessors 439 
    -- successors 445 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/word_access_0/rr
      -- 
    split_ack_5035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_gather_scatter_ack_0, ack => cp_elements(444)); -- 
    rr_5042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => ptr_deref_811_store_0_req_0); -- 
    -- CP-element group 445 fork  transition  input  no-bypass 
    -- predecessors 444 
    -- successors 446 783 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_request/word_access/word_access_0/ra
      -- 
    ra_5043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_store_0_ack_0, ack => cp_elements(445)); -- 
    -- CP-element group 446 transition  output  bypass 
    -- predecessors 445 
    -- successors 447 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/word_access_0/cr
      -- 
    cp_elements(446) <= cp_elements(445);
    cr_5053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(446), ack => ptr_deref_811_store_0_req_1); -- 
    -- CP-element group 447 transition  input  no-bypass 
    -- predecessors 446 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_813_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_811_complete/word_access/word_access_0/ca
      -- 
    ca_5054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_811_store_0_ack_1, ack => cp_elements(447)); -- 
    -- CP-element group 448 join  transition  output  bypass 
    -- predecessors 135 452 
    -- successors 453 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/word_access_0/rr
      -- 
    cpelement_group_448 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(135);
      predecessors(1) <= cp_elements(452);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(448)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(448),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(448), ack => ptr_deref_816_load_0_req_0); -- 
    -- CP-element group 449 transition  output  bypass 
    -- predecessors 41 
    -- successors 450 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_815_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_815_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_815_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_addr_resize/base_resize_req
      -- 
    cp_elements(449) <= cp_elements(41);
    base_resize_req_5071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => ptr_deref_816_base_resize_req_0); -- 
    -- CP-element group 450 transition  input  output  no-bypass 
    -- predecessors 449 
    -- successors 451 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_base_resize_ack_0, ack => cp_elements(450)); -- 
    sum_rename_req_5076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(450), ack => ptr_deref_816_root_address_inst_req_0); -- 
    -- CP-element group 451 transition  input  output  no-bypass 
    -- predecessors 450 
    -- successors 452 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_root_address_inst_ack_0, ack => cp_elements(451)); -- 
    root_register_req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(451), ack => ptr_deref_816_addr_0_req_0); -- 
    -- CP-element group 452 transition  input  no-bypass 
    -- predecessors 451 
    -- successors 448 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_word_addrgen/root_register_ack
      -- 
    root_register_ack_5082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_addr_0_ack_0, ack => cp_elements(452)); -- 
    -- CP-element group 453 transition  input  output  no-bypass 
    -- predecessors 448 
    -- successors 454 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/word_access_0/cr
      -- 
    ra_5093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_load_0_ack_0, ack => cp_elements(453)); -- 
    cr_5103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(453), ack => ptr_deref_816_load_0_req_1); -- 
    -- CP-element group 454 transition  input  output  no-bypass 
    -- predecessors 453 
    -- successors 455 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/merge_req
      -- 
    ca_5104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_load_0_ack_1, ack => cp_elements(454)); -- 
    merge_req_5105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(454), ack => ptr_deref_816_gather_scatter_req_0); -- 
    -- CP-element group 455 transition  input  output  no-bypass 
    -- predecessors 454 
    -- successors 456 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_817_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_817_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_817_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_816_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_819_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_819_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_819_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_complete/req
      -- 
    merge_ack_5106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_816_gather_scatter_ack_0, ack => cp_elements(455)); -- 
    req_5119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => type_cast_820_inst_req_0); -- 
    -- CP-element group 456 transition  input  output  no-bypass 
    -- predecessors 455 
    -- successors 459 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_821_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_821_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_821_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_820_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_823_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_823_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_823_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_resize_0/index_resize_req
      -- 
    ack_5120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_820_inst_ack_0, ack => cp_elements(456)); -- 
    index_resize_req_5138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(456), ack => array_obj_ref_824_index_0_resize_req_0); -- 
    -- CP-element group 457 transition  bypass 
    -- predecessors 41 
    -- successors 458 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_trigger_
      -- 
    cp_elements(457) <= cp_elements(41);
    -- CP-element group 458 join  transition  output  no-bypass 
    -- predecessors 457 462 
    -- successors 463 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_complete/final_reg_req
      -- 
    cpelement_group_458 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(457);
      predecessors(1) <= cp_elements(462);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(458)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(458),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5158_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => addr_of_825_final_reg_req_0); -- 
    -- CP-element group 459 transition  input  output  no-bypass 
    -- predecessors 456 
    -- successors 460 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_5139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_824_index_0_resize_ack_0, ack => cp_elements(459)); -- 
    scale_rename_req_5143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(459), ack => array_obj_ref_824_index_0_rename_req_0); -- 
    -- CP-element group 460 transition  input  output  no-bypass 
    -- predecessors 459 
    -- successors 461 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_add_indices/final_index_req
      -- 
    scale_rename_ack_5144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_824_index_0_rename_ack_0, ack => cp_elements(460)); -- 
    final_index_req_5148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => array_obj_ref_824_offset_inst_req_0); -- 
    -- CP-element group 461 transition  input  output  no-bypass 
    -- predecessors 460 
    -- successors 462 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_5149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_824_offset_inst_ack_0, ack => cp_elements(461)); -- 
    sum_rename_req_5153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => array_obj_ref_824_root_address_inst_req_0); -- 
    -- CP-element group 462 transition  input  no-bypass 
    -- predecessors 461 
    -- successors 458 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_824_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_5154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_824_root_address_inst_ack_0, ack => cp_elements(462)); -- 
    -- CP-element group 463 transition  input  output  no-bypass 
    -- predecessors 458 
    -- successors 464 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_826_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_826_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_826_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_825_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_828_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_828_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_828_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_5159_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_825_final_reg_ack_0, ack => cp_elements(463)); -- 
    base_resize_req_5176_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(463), ack => ptr_deref_829_base_resize_req_0); -- 
    -- CP-element group 464 transition  input  output  no-bypass 
    -- predecessors 463 
    -- successors 465 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5177_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_base_resize_ack_0, ack => cp_elements(464)); -- 
    sum_rename_req_5181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(464), ack => ptr_deref_829_root_address_inst_req_0); -- 
    -- CP-element group 465 transition  input  output  no-bypass 
    -- predecessors 464 
    -- successors 466 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_root_address_inst_ack_0, ack => cp_elements(465)); -- 
    root_register_req_5186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(465), ack => ptr_deref_829_addr_0_req_0); -- 
    -- CP-element group 466 transition  input  output  no-bypass 
    -- predecessors 465 
    -- successors 467 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/word_access_0/rr
      -- 
    root_register_ack_5187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_addr_0_ack_0, ack => cp_elements(466)); -- 
    rr_5197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(466), ack => ptr_deref_829_load_0_req_0); -- 
    -- CP-element group 467 transition  input  output  no-bypass 
    -- predecessors 466 
    -- successors 468 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/word_access_0/cr
      -- 
    ra_5198_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_load_0_ack_0, ack => cp_elements(467)); -- 
    cr_5208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => ptr_deref_829_load_0_req_1); -- 
    -- CP-element group 468 transition  input  output  no-bypass 
    -- predecessors 467 
    -- successors 469 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/merge_req
      -- 
    ca_5209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_load_0_ack_1, ack => cp_elements(468)); -- 
    merge_req_5210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(468), ack => ptr_deref_829_gather_scatter_req_0); -- 
    -- CP-element group 469 transition  input  no-bypass 
    -- predecessors 468 
    -- successors 492 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_830_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_830_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_830_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_829_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_849_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_849_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_849_completed_
      -- 
    merge_ack_5211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_829_gather_scatter_ack_0, ack => cp_elements(469)); -- 
    -- CP-element group 470 join  transition  output  bypass 
    -- predecessors 135 474 
    -- successors 475 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/word_access_0/rr
      -- 
    cpelement_group_470 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(135);
      predecessors(1) <= cp_elements(474);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(470)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(470),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(470), ack => ptr_deref_833_load_0_req_0); -- 
    -- CP-element group 471 transition  output  bypass 
    -- predecessors 41 
    -- successors 472 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_832_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_832_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_832_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_addr_resize/base_resize_req
      -- 
    cp_elements(471) <= cp_elements(41);
    base_resize_req_5228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(471), ack => ptr_deref_833_base_resize_req_0); -- 
    -- CP-element group 472 transition  input  output  no-bypass 
    -- predecessors 471 
    -- successors 473 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_base_resize_ack_0, ack => cp_elements(472)); -- 
    sum_rename_req_5233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(472), ack => ptr_deref_833_root_address_inst_req_0); -- 
    -- CP-element group 473 transition  input  output  no-bypass 
    -- predecessors 472 
    -- successors 474 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_root_address_inst_ack_0, ack => cp_elements(473)); -- 
    root_register_req_5238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(473), ack => ptr_deref_833_addr_0_req_0); -- 
    -- CP-element group 474 transition  input  no-bypass 
    -- predecessors 473 
    -- successors 470 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_word_addrgen/root_register_ack
      -- 
    root_register_ack_5239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_addr_0_ack_0, ack => cp_elements(474)); -- 
    -- CP-element group 475 transition  input  output  no-bypass 
    -- predecessors 470 
    -- successors 476 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/word_access_0/cr
      -- 
    ra_5250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_load_0_ack_0, ack => cp_elements(475)); -- 
    cr_5260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(475), ack => ptr_deref_833_load_0_req_1); -- 
    -- CP-element group 476 transition  input  output  no-bypass 
    -- predecessors 475 
    -- successors 477 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/merge_req
      -- 
    ca_5261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_load_0_ack_1, ack => cp_elements(476)); -- 
    merge_req_5262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(476), ack => ptr_deref_833_gather_scatter_req_0); -- 
    -- CP-element group 477 transition  input  output  no-bypass 
    -- predecessors 476 
    -- successors 478 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_834_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_834_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_834_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_833_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_836_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_836_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_836_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_complete/req
      -- 
    merge_ack_5263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_833_gather_scatter_ack_0, ack => cp_elements(477)); -- 
    req_5276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => type_cast_837_inst_req_0); -- 
    -- CP-element group 478 transition  input  output  no-bypass 
    -- predecessors 477 
    -- successors 481 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_838_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_838_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_838_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_837_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_840_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_840_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_840_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_resize_0/index_resize_req
      -- 
    ack_5277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_837_inst_ack_0, ack => cp_elements(478)); -- 
    index_resize_req_5295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(478), ack => array_obj_ref_841_index_0_resize_req_0); -- 
    -- CP-element group 479 transition  bypass 
    -- predecessors 41 
    -- successors 480 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_trigger_
      -- 
    cp_elements(479) <= cp_elements(41);
    -- CP-element group 480 join  transition  output  no-bypass 
    -- predecessors 479 484 
    -- successors 485 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_complete/final_reg_req
      -- 
    cpelement_group_480 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(479);
      predecessors(1) <= cp_elements(484);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(480)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(480),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(480), ack => addr_of_842_final_reg_req_0); -- 
    -- CP-element group 481 transition  input  output  no-bypass 
    -- predecessors 478 
    -- successors 482 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_5296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_index_0_resize_ack_0, ack => cp_elements(481)); -- 
    scale_rename_req_5300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(481), ack => array_obj_ref_841_index_0_rename_req_0); -- 
    -- CP-element group 482 transition  input  output  no-bypass 
    -- predecessors 481 
    -- successors 483 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_add_indices/final_index_req
      -- 
    scale_rename_ack_5301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_index_0_rename_ack_0, ack => cp_elements(482)); -- 
    final_index_req_5305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(482), ack => array_obj_ref_841_offset_inst_req_0); -- 
    -- CP-element group 483 transition  input  output  no-bypass 
    -- predecessors 482 
    -- successors 484 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_5306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_offset_inst_ack_0, ack => cp_elements(483)); -- 
    sum_rename_req_5310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(483), ack => array_obj_ref_841_root_address_inst_req_0); -- 
    -- CP-element group 484 transition  input  no-bypass 
    -- predecessors 483 
    -- successors 480 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_841_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_5311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_841_root_address_inst_ack_0, ack => cp_elements(484)); -- 
    -- CP-element group 485 transition  input  output  no-bypass 
    -- predecessors 480 
    -- successors 486 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_843_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_843_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_843_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_842_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_845_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_845_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_845_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_5316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_842_final_reg_ack_0, ack => cp_elements(485)); -- 
    base_resize_req_5333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(485), ack => ptr_deref_846_base_resize_req_0); -- 
    -- CP-element group 486 transition  input  output  no-bypass 
    -- predecessors 485 
    -- successors 487 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_base_resize_ack_0, ack => cp_elements(486)); -- 
    sum_rename_req_5338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(486), ack => ptr_deref_846_root_address_inst_req_0); -- 
    -- CP-element group 487 transition  input  output  no-bypass 
    -- predecessors 486 
    -- successors 488 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_root_address_inst_ack_0, ack => cp_elements(487)); -- 
    root_register_req_5343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(487), ack => ptr_deref_846_addr_0_req_0); -- 
    -- CP-element group 488 transition  input  output  no-bypass 
    -- predecessors 487 
    -- successors 489 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/word_access_0/rr
      -- 
    root_register_ack_5344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_addr_0_ack_0, ack => cp_elements(488)); -- 
    rr_5354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(488), ack => ptr_deref_846_load_0_req_0); -- 
    -- CP-element group 489 transition  input  output  no-bypass 
    -- predecessors 488 
    -- successors 490 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/word_access_0/cr
      -- 
    ra_5355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_load_0_ack_0, ack => cp_elements(489)); -- 
    cr_5365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(489), ack => ptr_deref_846_load_0_req_1); -- 
    -- CP-element group 490 transition  input  output  no-bypass 
    -- predecessors 489 
    -- successors 491 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/merge_req
      -- 
    ca_5366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_load_0_ack_1, ack => cp_elements(490)); -- 
    merge_req_5367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => ptr_deref_846_gather_scatter_req_0); -- 
    -- CP-element group 491 transition  input  no-bypass 
    -- predecessors 490 
    -- successors 492 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_847_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_847_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_847_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_846_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_850_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_850_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_850_completed_
      -- 
    merge_ack_5368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_846_gather_scatter_ack_0, ack => cp_elements(491)); -- 
    -- CP-element group 492 join  fork  transition  bypass 
    -- predecessors 469 491 
    -- successors 495 496 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_trigger_
      -- 
    cpelement_group_492 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(469);
      predecessors(1) <= cp_elements(491);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(492)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(492),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 493 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_active_
      -- 
    cp_elements(493) <= cp_elements(41);
    -- CP-element group 494 join  transition  bypass 
    -- predecessors 497 498 
    -- successors 499 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_852_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_852_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_852_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_856_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_856_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_855_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_855_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_855_completed_
      -- 
    cpelement_group_494 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(497);
      predecessors(1) <= cp_elements(498);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(494)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(494),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 495 transition  output  bypass 
    -- predecessors 492 
    -- successors 497 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Sample/rr
      -- 
    cp_elements(495) <= cp_elements(492);
    rr_5388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(495), ack => binary_851_inst_req_0); -- 
    -- CP-element group 496 transition  output  bypass 
    -- predecessors 492 
    -- successors 498 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Update/cr
      -- 
    cp_elements(496) <= cp_elements(492);
    cr_5393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => binary_851_inst_req_1); -- 
    -- CP-element group 497 transition  input  no-bypass 
    -- predecessors 495 
    -- successors 494 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Sample/ra
      -- 
    ra_5389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_851_inst_ack_0, ack => cp_elements(497)); -- 
    -- CP-element group 498 transition  input  no-bypass 
    -- predecessors 496 
    -- successors 494 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_851_Update/ca
      -- 
    ca_5394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_851_inst_ack_1, ack => cp_elements(498)); -- 
    -- CP-element group 499 join  transition  output  bypass 
    -- predecessors 494 503 
    -- successors 504 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/split_req
      -- 
    cpelement_group_499 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(494);
      predecessors(1) <= cp_elements(503);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(499)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(499),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => ptr_deref_854_gather_scatter_req_0); -- 
    -- CP-element group 500 transition  output  bypass 
    -- predecessors 41 
    -- successors 501 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_853_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_853_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_853_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_addr_resize/base_resize_req
      -- 
    cp_elements(500) <= cp_elements(41);
    base_resize_req_5414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ptr_deref_854_base_resize_req_0); -- 
    -- CP-element group 501 transition  input  output  no-bypass 
    -- predecessors 500 
    -- successors 502 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_base_resize_ack_0, ack => cp_elements(501)); -- 
    sum_rename_req_5419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => ptr_deref_854_root_address_inst_req_0); -- 
    -- CP-element group 502 transition  input  output  no-bypass 
    -- predecessors 501 
    -- successors 503 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_root_address_inst_ack_0, ack => cp_elements(502)); -- 
    root_register_req_5424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(502), ack => ptr_deref_854_addr_0_req_0); -- 
    -- CP-element group 503 transition  input  no-bypass 
    -- predecessors 502 
    -- successors 499 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_word_addrgen/root_register_ack
      -- 
    root_register_ack_5425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_addr_0_ack_0, ack => cp_elements(503)); -- 
    -- CP-element group 504 transition  input  output  no-bypass 
    -- predecessors 499 
    -- successors 505 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/word_access_0/rr
      -- 
    split_ack_5430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_gather_scatter_ack_0, ack => cp_elements(504)); -- 
    rr_5437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(504), ack => ptr_deref_854_store_0_req_0); -- 
    -- CP-element group 505 fork  transition  input  no-bypass 
    -- predecessors 504 
    -- successors 506 815 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_request/word_access/word_access_0/ra
      -- 
    ra_5438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_store_0_ack_0, ack => cp_elements(505)); -- 
    -- CP-element group 506 transition  output  bypass 
    -- predecessors 505 
    -- successors 507 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/word_access_0/cr
      -- 
    cp_elements(506) <= cp_elements(505);
    cr_5448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_854_store_0_req_1); -- 
    -- CP-element group 507 transition  input  no-bypass 
    -- predecessors 506 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_856_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_854_complete/word_access/word_access_0/ca
      -- 
    ca_5449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_854_store_0_ack_1, ack => cp_elements(507)); -- 
    -- CP-element group 508 join  transition  output  bypass 
    -- predecessors 159 512 
    -- successors 513 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/word_access_0/rr
      -- 
    cpelement_group_508 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(159);
      predecessors(1) <= cp_elements(512);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(508)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(508),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5487_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(508), ack => ptr_deref_859_load_0_req_0); -- 
    -- CP-element group 509 transition  output  bypass 
    -- predecessors 41 
    -- successors 510 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_858_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_858_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_858_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_addr_resize/base_resize_req
      -- 
    cp_elements(509) <= cp_elements(41);
    base_resize_req_5466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ptr_deref_859_base_resize_req_0); -- 
    -- CP-element group 510 transition  input  output  no-bypass 
    -- predecessors 509 
    -- successors 511 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_base_resize_ack_0, ack => cp_elements(510)); -- 
    sum_rename_req_5471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(510), ack => ptr_deref_859_root_address_inst_req_0); -- 
    -- CP-element group 511 transition  input  output  no-bypass 
    -- predecessors 510 
    -- successors 512 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_root_address_inst_ack_0, ack => cp_elements(511)); -- 
    root_register_req_5476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(511), ack => ptr_deref_859_addr_0_req_0); -- 
    -- CP-element group 512 transition  input  no-bypass 
    -- predecessors 511 
    -- successors 508 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_word_addrgen/root_register_ack
      -- 
    root_register_ack_5477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_addr_0_ack_0, ack => cp_elements(512)); -- 
    -- CP-element group 513 transition  input  output  no-bypass 
    -- predecessors 508 
    -- successors 514 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/word_access_0/cr
      -- 
    ra_5488_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_load_0_ack_0, ack => cp_elements(513)); -- 
    cr_5498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(513), ack => ptr_deref_859_load_0_req_1); -- 
    -- CP-element group 514 transition  input  output  no-bypass 
    -- predecessors 513 
    -- successors 515 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/merge_req
      -- 
    ca_5499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_load_0_ack_1, ack => cp_elements(514)); -- 
    merge_req_5500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => ptr_deref_859_gather_scatter_req_0); -- 
    -- CP-element group 515 transition  input  output  no-bypass 
    -- predecessors 514 
    -- successors 516 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_860_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_860_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_860_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_859_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_862_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_862_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_862_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_complete/req
      -- 
    merge_ack_5501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_859_gather_scatter_ack_0, ack => cp_elements(515)); -- 
    req_5514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => type_cast_863_inst_req_0); -- 
    -- CP-element group 516 transition  input  output  no-bypass 
    -- predecessors 515 
    -- successors 519 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_864_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_864_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_864_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_863_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_866_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_866_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_866_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_resize_0/index_resize_req
      -- 
    ack_5515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => cp_elements(516)); -- 
    index_resize_req_5533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(516), ack => array_obj_ref_867_index_0_resize_req_0); -- 
    -- CP-element group 517 transition  bypass 
    -- predecessors 41 
    -- successors 518 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_trigger_
      -- 
    cp_elements(517) <= cp_elements(41);
    -- CP-element group 518 join  transition  output  no-bypass 
    -- predecessors 517 522 
    -- successors 523 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_complete/final_reg_req
      -- 
    cpelement_group_518 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(517);
      predecessors(1) <= cp_elements(522);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(518)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(518), ack => addr_of_868_final_reg_req_0); -- 
    -- CP-element group 519 transition  input  output  no-bypass 
    -- predecessors 516 
    -- successors 520 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_5534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_867_index_0_resize_ack_0, ack => cp_elements(519)); -- 
    scale_rename_req_5538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => array_obj_ref_867_index_0_rename_req_0); -- 
    -- CP-element group 520 transition  input  output  no-bypass 
    -- predecessors 519 
    -- successors 521 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_add_indices/final_index_req
      -- 
    scale_rename_ack_5539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_867_index_0_rename_ack_0, ack => cp_elements(520)); -- 
    final_index_req_5543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(520), ack => array_obj_ref_867_offset_inst_req_0); -- 
    -- CP-element group 521 transition  input  output  no-bypass 
    -- predecessors 520 
    -- successors 522 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_5544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_867_offset_inst_ack_0, ack => cp_elements(521)); -- 
    sum_rename_req_5548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(521), ack => array_obj_ref_867_root_address_inst_req_0); -- 
    -- CP-element group 522 transition  input  no-bypass 
    -- predecessors 521 
    -- successors 518 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_867_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_5549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_867_root_address_inst_ack_0, ack => cp_elements(522)); -- 
    -- CP-element group 523 transition  input  output  no-bypass 
    -- predecessors 518 
    -- successors 524 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_869_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_869_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_869_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_868_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_871_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_871_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_871_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_5554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_868_final_reg_ack_0, ack => cp_elements(523)); -- 
    base_resize_req_5571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => ptr_deref_872_base_resize_req_0); -- 
    -- CP-element group 524 transition  input  output  no-bypass 
    -- predecessors 523 
    -- successors 525 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_base_resize_ack_0, ack => cp_elements(524)); -- 
    sum_rename_req_5576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => ptr_deref_872_root_address_inst_req_0); -- 
    -- CP-element group 525 transition  input  output  no-bypass 
    -- predecessors 524 
    -- successors 526 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_root_address_inst_ack_0, ack => cp_elements(525)); -- 
    root_register_req_5581_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(525), ack => ptr_deref_872_addr_0_req_0); -- 
    -- CP-element group 526 transition  input  output  no-bypass 
    -- predecessors 525 
    -- successors 527 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/word_access_0/rr
      -- 
    root_register_ack_5582_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_addr_0_ack_0, ack => cp_elements(526)); -- 
    rr_5592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(526), ack => ptr_deref_872_load_0_req_0); -- 
    -- CP-element group 527 transition  input  output  no-bypass 
    -- predecessors 526 
    -- successors 528 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/word_access_0/cr
      -- 
    ra_5593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_load_0_ack_0, ack => cp_elements(527)); -- 
    cr_5603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(527), ack => ptr_deref_872_load_0_req_1); -- 
    -- CP-element group 528 transition  input  output  no-bypass 
    -- predecessors 527 
    -- successors 529 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/merge_req
      -- 
    ca_5604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_load_0_ack_1, ack => cp_elements(528)); -- 
    merge_req_5605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => ptr_deref_872_gather_scatter_req_0); -- 
    -- CP-element group 529 transition  input  no-bypass 
    -- predecessors 528 
    -- successors 552 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_873_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_873_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_873_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_872_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_892_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_892_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_892_completed_
      -- 
    merge_ack_5606_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_872_gather_scatter_ack_0, ack => cp_elements(529)); -- 
    -- CP-element group 530 join  transition  output  bypass 
    -- predecessors 159 534 
    -- successors 535 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/word_access_0/rr
      -- 
    cpelement_group_530 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(159);
      predecessors(1) <= cp_elements(534);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(530)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(530),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(530), ack => ptr_deref_876_load_0_req_0); -- 
    -- CP-element group 531 transition  output  bypass 
    -- predecessors 41 
    -- successors 532 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_875_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_875_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_875_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_addr_resize/base_resize_req
      -- 
    cp_elements(531) <= cp_elements(41);
    base_resize_req_5623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(531), ack => ptr_deref_876_base_resize_req_0); -- 
    -- CP-element group 532 transition  input  output  no-bypass 
    -- predecessors 531 
    -- successors 533 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_base_resize_ack_0, ack => cp_elements(532)); -- 
    sum_rename_req_5628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => ptr_deref_876_root_address_inst_req_0); -- 
    -- CP-element group 533 transition  input  output  no-bypass 
    -- predecessors 532 
    -- successors 534 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_root_address_inst_ack_0, ack => cp_elements(533)); -- 
    root_register_req_5633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(533), ack => ptr_deref_876_addr_0_req_0); -- 
    -- CP-element group 534 transition  input  no-bypass 
    -- predecessors 533 
    -- successors 530 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_word_addrgen/root_register_ack
      -- 
    root_register_ack_5634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_addr_0_ack_0, ack => cp_elements(534)); -- 
    -- CP-element group 535 transition  input  output  no-bypass 
    -- predecessors 530 
    -- successors 536 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/word_access_0/cr
      -- 
    ra_5645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_load_0_ack_0, ack => cp_elements(535)); -- 
    cr_5655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => ptr_deref_876_load_0_req_1); -- 
    -- CP-element group 536 transition  input  output  no-bypass 
    -- predecessors 535 
    -- successors 537 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/merge_req
      -- 
    ca_5656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_load_0_ack_1, ack => cp_elements(536)); -- 
    merge_req_5657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(536), ack => ptr_deref_876_gather_scatter_req_0); -- 
    -- CP-element group 537 transition  input  output  no-bypass 
    -- predecessors 536 
    -- successors 538 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_877_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_877_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_877_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_876_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_879_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_879_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_879_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_complete/req
      -- 
    merge_ack_5658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_876_gather_scatter_ack_0, ack => cp_elements(537)); -- 
    req_5671_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(537), ack => type_cast_880_inst_req_0); -- 
    -- CP-element group 538 transition  input  output  no-bypass 
    -- predecessors 537 
    -- successors 541 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_881_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_881_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_881_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_880_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_883_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_883_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_883_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_resize_0/index_resize_req
      -- 
    ack_5672_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_880_inst_ack_0, ack => cp_elements(538)); -- 
    index_resize_req_5690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => array_obj_ref_884_index_0_resize_req_0); -- 
    -- CP-element group 539 transition  bypass 
    -- predecessors 41 
    -- successors 540 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_trigger_
      -- 
    cp_elements(539) <= cp_elements(41);
    -- CP-element group 540 join  transition  output  no-bypass 
    -- predecessors 539 544 
    -- successors 545 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_complete/final_reg_req
      -- 
    cpelement_group_540 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(539);
      predecessors(1) <= cp_elements(544);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(540)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(540),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5710_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(540), ack => addr_of_885_final_reg_req_0); -- 
    -- CP-element group 541 transition  input  output  no-bypass 
    -- predecessors 538 
    -- successors 542 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_5691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_0_resize_ack_0, ack => cp_elements(541)); -- 
    scale_rename_req_5695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => array_obj_ref_884_index_0_rename_req_0); -- 
    -- CP-element group 542 transition  input  output  no-bypass 
    -- predecessors 541 
    -- successors 543 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_add_indices/final_index_req
      -- 
    scale_rename_ack_5696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_index_0_rename_ack_0, ack => cp_elements(542)); -- 
    final_index_req_5700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(542), ack => array_obj_ref_884_offset_inst_req_0); -- 
    -- CP-element group 543 transition  input  output  no-bypass 
    -- predecessors 542 
    -- successors 544 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_5701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_offset_inst_ack_0, ack => cp_elements(543)); -- 
    sum_rename_req_5705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(543), ack => array_obj_ref_884_root_address_inst_req_0); -- 
    -- CP-element group 544 transition  input  no-bypass 
    -- predecessors 543 
    -- successors 540 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_884_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_5706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_884_root_address_inst_ack_0, ack => cp_elements(544)); -- 
    -- CP-element group 545 transition  input  output  no-bypass 
    -- predecessors 540 
    -- successors 546 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_886_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_886_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_886_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_885_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_888_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_888_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_888_completed_
      -- 
    final_reg_ack_5711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_885_final_reg_ack_0, ack => cp_elements(545)); -- 
    base_resize_req_5728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => ptr_deref_889_base_resize_req_0); -- 
    -- CP-element group 546 transition  input  output  no-bypass 
    -- predecessors 545 
    -- successors 547 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_base_resize_ack_0, ack => cp_elements(546)); -- 
    sum_rename_req_5733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(546), ack => ptr_deref_889_root_address_inst_req_0); -- 
    -- CP-element group 547 transition  input  output  no-bypass 
    -- predecessors 546 
    -- successors 548 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_root_address_inst_ack_0, ack => cp_elements(547)); -- 
    root_register_req_5738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => ptr_deref_889_addr_0_req_0); -- 
    -- CP-element group 548 transition  input  output  no-bypass 
    -- predecessors 547 
    -- successors 549 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_word_address_calculated
      -- 
    root_register_ack_5739_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_addr_0_ack_0, ack => cp_elements(548)); -- 
    rr_5749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => ptr_deref_889_load_0_req_0); -- 
    -- CP-element group 549 transition  input  output  no-bypass 
    -- predecessors 548 
    -- successors 550 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_active_
      -- 
    ra_5750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_load_0_ack_0, ack => cp_elements(549)); -- 
    cr_5760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => ptr_deref_889_load_0_req_1); -- 
    -- CP-element group 550 transition  input  output  no-bypass 
    -- predecessors 549 
    -- successors 551 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/merge_req
      -- 
    ca_5761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_load_0_ack_1, ack => cp_elements(550)); -- 
    merge_req_5762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => ptr_deref_889_gather_scatter_req_0); -- 
    -- CP-element group 551 transition  input  no-bypass 
    -- predecessors 550 
    -- successors 552 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_890_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_890_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_890_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_889_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_893_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_893_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_893_completed_
      -- 
    merge_ack_5763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_889_gather_scatter_ack_0, ack => cp_elements(551)); -- 
    -- CP-element group 552 join  fork  transition  bypass 
    -- predecessors 529 551 
    -- successors 555 556 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_trigger_
      -- 
    cpelement_group_552 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(529);
      predecessors(1) <= cp_elements(551);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(552)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(552),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 553 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_active_
      -- 
    cp_elements(553) <= cp_elements(41);
    -- CP-element group 554 join  transition  bypass 
    -- predecessors 557 558 
    -- successors 559 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_895_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_895_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_895_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_899_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_899_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_898_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_898_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_898_completed_
      -- 
    cpelement_group_554 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(557);
      predecessors(1) <= cp_elements(558);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(554)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(554),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 555 transition  output  bypass 
    -- predecessors 552 
    -- successors 557 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Sample/rr
      -- 
    cp_elements(555) <= cp_elements(552);
    rr_5783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(555), ack => binary_894_inst_req_0); -- 
    -- CP-element group 556 transition  output  bypass 
    -- predecessors 552 
    -- successors 558 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Update/cr
      -- 
    cp_elements(556) <= cp_elements(552);
    cr_5788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => binary_894_inst_req_1); -- 
    -- CP-element group 557 transition  input  no-bypass 
    -- predecessors 555 
    -- successors 554 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Sample/ra
      -- 
    ra_5784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_894_inst_ack_0, ack => cp_elements(557)); -- 
    -- CP-element group 558 transition  input  no-bypass 
    -- predecessors 556 
    -- successors 554 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_894_Update/ca
      -- 
    ca_5789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_894_inst_ack_1, ack => cp_elements(558)); -- 
    -- CP-element group 559 join  transition  output  bypass 
    -- predecessors 554 563 
    -- successors 564 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/split_req
      -- 
    cpelement_group_559 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(554);
      predecessors(1) <= cp_elements(563);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(559)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(559),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => ptr_deref_897_gather_scatter_req_0); -- 
    -- CP-element group 560 transition  output  bypass 
    -- predecessors 41 
    -- successors 561 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_896_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_896_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_896_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_addr_resize/base_resize_req
      -- 
    cp_elements(560) <= cp_elements(41);
    base_resize_req_5809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(560), ack => ptr_deref_897_base_resize_req_0); -- 
    -- CP-element group 561 transition  input  output  no-bypass 
    -- predecessors 560 
    -- successors 562 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_base_resize_ack_0, ack => cp_elements(561)); -- 
    sum_rename_req_5814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => ptr_deref_897_root_address_inst_req_0); -- 
    -- CP-element group 562 transition  input  output  no-bypass 
    -- predecessors 561 
    -- successors 563 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_root_address_inst_ack_0, ack => cp_elements(562)); -- 
    root_register_req_5819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(562), ack => ptr_deref_897_addr_0_req_0); -- 
    -- CP-element group 563 transition  input  no-bypass 
    -- predecessors 562 
    -- successors 559 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_word_addrgen/root_register_ack
      -- 
    root_register_ack_5820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_addr_0_ack_0, ack => cp_elements(563)); -- 
    -- CP-element group 564 transition  input  output  no-bypass 
    -- predecessors 559 
    -- successors 565 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/word_access_0/rr
      -- 
    split_ack_5825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_gather_scatter_ack_0, ack => cp_elements(564)); -- 
    rr_5832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => ptr_deref_897_store_0_req_0); -- 
    -- CP-element group 565 fork  transition  input  no-bypass 
    -- predecessors 564 
    -- successors 566 847 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_request/word_access/word_access_0/ra
      -- 
    ra_5833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_store_0_ack_0, ack => cp_elements(565)); -- 
    -- CP-element group 566 transition  output  bypass 
    -- predecessors 565 
    -- successors 567 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/word_access_0/cr
      -- 
    cp_elements(566) <= cp_elements(565);
    cr_5843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => ptr_deref_897_store_0_req_1); -- 
    -- CP-element group 567 transition  input  no-bypass 
    -- predecessors 566 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_899_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_897_complete/word_access/word_access_0/ca
      -- 
    ca_5844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_897_store_0_ack_1, ack => cp_elements(567)); -- 
    -- CP-element group 568 join  transition  output  bypass 
    -- predecessors 183 572 
    -- successors 573 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/word_access_0/rr
      -- 
    cpelement_group_568 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(183);
      predecessors(1) <= cp_elements(572);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(568)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(568),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_902_load_0_req_0); -- 
    -- CP-element group 569 transition  output  bypass 
    -- predecessors 41 
    -- successors 570 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_901_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_901_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_901_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_addr_resize/base_resize_req
      -- 
    cp_elements(569) <= cp_elements(41);
    base_resize_req_5861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => ptr_deref_902_base_resize_req_0); -- 
    -- CP-element group 570 transition  input  output  no-bypass 
    -- predecessors 569 
    -- successors 571 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_base_resize_ack_0, ack => cp_elements(570)); -- 
    sum_rename_req_5866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(570), ack => ptr_deref_902_root_address_inst_req_0); -- 
    -- CP-element group 571 transition  input  output  no-bypass 
    -- predecessors 570 
    -- successors 572 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_root_address_inst_ack_0, ack => cp_elements(571)); -- 
    root_register_req_5871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => ptr_deref_902_addr_0_req_0); -- 
    -- CP-element group 572 transition  input  no-bypass 
    -- predecessors 571 
    -- successors 568 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_word_addrgen/root_register_ack
      -- 
    root_register_ack_5872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_addr_0_ack_0, ack => cp_elements(572)); -- 
    -- CP-element group 573 transition  input  output  no-bypass 
    -- predecessors 568 
    -- successors 574 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/word_access_0/cr
      -- 
    ra_5883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_load_0_ack_0, ack => cp_elements(573)); -- 
    cr_5893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(573), ack => ptr_deref_902_load_0_req_1); -- 
    -- CP-element group 574 transition  input  output  no-bypass 
    -- predecessors 573 
    -- successors 575 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/merge_req
      -- 
    ca_5894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_load_0_ack_1, ack => cp_elements(574)); -- 
    merge_req_5895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => ptr_deref_902_gather_scatter_req_0); -- 
    -- CP-element group 575 transition  input  output  no-bypass 
    -- predecessors 574 
    -- successors 576 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_903_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_903_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_903_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_902_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_905_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_905_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_905_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_complete/req
      -- 
    merge_ack_5896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_902_gather_scatter_ack_0, ack => cp_elements(575)); -- 
    req_5909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => type_cast_906_inst_req_0); -- 
    -- CP-element group 576 transition  input  output  no-bypass 
    -- predecessors 575 
    -- successors 579 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_907_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_907_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_907_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_906_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_909_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_909_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_909_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_resize_0/index_resize_req
      -- 
    ack_5910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_906_inst_ack_0, ack => cp_elements(576)); -- 
    index_resize_req_5928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(576), ack => array_obj_ref_910_index_0_resize_req_0); -- 
    -- CP-element group 577 transition  bypass 
    -- predecessors 41 
    -- successors 578 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_trigger_
      -- 
    cp_elements(577) <= cp_elements(41);
    -- CP-element group 578 join  transition  output  no-bypass 
    -- predecessors 577 582 
    -- successors 583 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_complete/final_reg_req
      -- 
    cpelement_group_578 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(577);
      predecessors(1) <= cp_elements(582);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(578)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(578),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => addr_of_911_final_reg_req_0); -- 
    -- CP-element group 579 transition  input  output  no-bypass 
    -- predecessors 576 
    -- successors 580 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_5929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_910_index_0_resize_ack_0, ack => cp_elements(579)); -- 
    scale_rename_req_5933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(579), ack => array_obj_ref_910_index_0_rename_req_0); -- 
    -- CP-element group 580 transition  input  output  no-bypass 
    -- predecessors 579 
    -- successors 581 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_add_indices/final_index_req
      -- 
    scale_rename_ack_5934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_910_index_0_rename_ack_0, ack => cp_elements(580)); -- 
    final_index_req_5938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(580), ack => array_obj_ref_910_offset_inst_req_0); -- 
    -- CP-element group 581 transition  input  output  no-bypass 
    -- predecessors 580 
    -- successors 582 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_5939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_910_offset_inst_ack_0, ack => cp_elements(581)); -- 
    sum_rename_req_5943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(581), ack => array_obj_ref_910_root_address_inst_req_0); -- 
    -- CP-element group 582 transition  input  no-bypass 
    -- predecessors 581 
    -- successors 578 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_910_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_5944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_910_root_address_inst_ack_0, ack => cp_elements(582)); -- 
    -- CP-element group 583 transition  input  output  no-bypass 
    -- predecessors 578 
    -- successors 584 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_912_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_912_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_912_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_911_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_914_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_914_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_914_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_5949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_911_final_reg_ack_0, ack => cp_elements(583)); -- 
    base_resize_req_5966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(583), ack => ptr_deref_915_base_resize_req_0); -- 
    -- CP-element group 584 transition  input  output  no-bypass 
    -- predecessors 583 
    -- successors 585 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_5967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_base_resize_ack_0, ack => cp_elements(584)); -- 
    sum_rename_req_5971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => ptr_deref_915_root_address_inst_req_0); -- 
    -- CP-element group 585 transition  input  output  no-bypass 
    -- predecessors 584 
    -- successors 586 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_word_addrgen/root_register_req
      -- 
    sum_rename_ack_5972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_root_address_inst_ack_0, ack => cp_elements(585)); -- 
    root_register_req_5976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(585), ack => ptr_deref_915_addr_0_req_0); -- 
    -- CP-element group 586 transition  input  output  no-bypass 
    -- predecessors 585 
    -- successors 587 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/word_access_0/rr
      -- 
    root_register_ack_5977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_addr_0_ack_0, ack => cp_elements(586)); -- 
    rr_5987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ptr_deref_915_load_0_req_0); -- 
    -- CP-element group 587 transition  input  output  no-bypass 
    -- predecessors 586 
    -- successors 588 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/word_access_0/cr
      -- 
    ra_5988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_load_0_ack_0, ack => cp_elements(587)); -- 
    cr_5998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => ptr_deref_915_load_0_req_1); -- 
    -- CP-element group 588 transition  input  output  no-bypass 
    -- predecessors 587 
    -- successors 589 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/merge_req
      -- 
    ca_5999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_load_0_ack_1, ack => cp_elements(588)); -- 
    merge_req_6000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(588), ack => ptr_deref_915_gather_scatter_req_0); -- 
    -- CP-element group 589 transition  input  no-bypass 
    -- predecessors 588 
    -- successors 612 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_916_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_916_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_916_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_915_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_935_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_935_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_935_completed_
      -- 
    merge_ack_6001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_915_gather_scatter_ack_0, ack => cp_elements(589)); -- 
    -- CP-element group 590 join  transition  output  bypass 
    -- predecessors 183 594 
    -- successors 595 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/word_access_0/rr
      -- 
    cpelement_group_590 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(183);
      predecessors(1) <= cp_elements(594);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(590)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(590),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6039_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(590), ack => ptr_deref_919_load_0_req_0); -- 
    -- CP-element group 591 transition  output  bypass 
    -- predecessors 41 
    -- successors 592 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_918_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_918_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_918_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_addr_resize/base_resize_req
      -- 
    cp_elements(591) <= cp_elements(41);
    base_resize_req_6018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => ptr_deref_919_base_resize_req_0); -- 
    -- CP-element group 592 transition  input  output  no-bypass 
    -- predecessors 591 
    -- successors 593 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_base_resize_ack_0, ack => cp_elements(592)); -- 
    sum_rename_req_6023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(592), ack => ptr_deref_919_root_address_inst_req_0); -- 
    -- CP-element group 593 transition  input  output  no-bypass 
    -- predecessors 592 
    -- successors 594 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_root_address_inst_ack_0, ack => cp_elements(593)); -- 
    root_register_req_6028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_919_addr_0_req_0); -- 
    -- CP-element group 594 transition  input  no-bypass 
    -- predecessors 593 
    -- successors 590 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_word_addrgen/root_register_ack
      -- 
    root_register_ack_6029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_addr_0_ack_0, ack => cp_elements(594)); -- 
    -- CP-element group 595 transition  input  output  no-bypass 
    -- predecessors 590 
    -- successors 596 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/word_access_0/cr
      -- 
    ra_6040_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_load_0_ack_0, ack => cp_elements(595)); -- 
    cr_6050_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => ptr_deref_919_load_0_req_1); -- 
    -- CP-element group 596 transition  input  output  no-bypass 
    -- predecessors 595 
    -- successors 597 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/merge_req
      -- 
    ca_6051_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_load_0_ack_1, ack => cp_elements(596)); -- 
    merge_req_6052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(596), ack => ptr_deref_919_gather_scatter_req_0); -- 
    -- CP-element group 597 transition  input  output  no-bypass 
    -- predecessors 596 
    -- successors 598 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_920_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_920_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_920_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_919_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_922_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_922_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_922_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_complete/req
      -- 
    merge_ack_6053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_919_gather_scatter_ack_0, ack => cp_elements(597)); -- 
    req_6066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(597), ack => type_cast_923_inst_req_0); -- 
    -- CP-element group 598 transition  input  output  no-bypass 
    -- predecessors 597 
    -- successors 601 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_924_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_924_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_924_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_923_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_926_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_926_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_926_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_resize_0/index_resize_req
      -- 
    ack_6067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_923_inst_ack_0, ack => cp_elements(598)); -- 
    index_resize_req_6085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(598), ack => array_obj_ref_927_index_0_resize_req_0); -- 
    -- CP-element group 599 transition  bypass 
    -- predecessors 41 
    -- successors 600 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_trigger_
      -- 
    cp_elements(599) <= cp_elements(41);
    -- CP-element group 600 join  transition  output  no-bypass 
    -- predecessors 599 604 
    -- successors 605 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_complete/final_reg_req
      -- 
    cpelement_group_600 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(599);
      predecessors(1) <= cp_elements(604);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(600)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => addr_of_928_final_reg_req_0); -- 
    -- CP-element group 601 transition  input  output  no-bypass 
    -- predecessors 598 
    -- successors 602 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_6086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_927_index_0_resize_ack_0, ack => cp_elements(601)); -- 
    scale_rename_req_6090_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(601), ack => array_obj_ref_927_index_0_rename_req_0); -- 
    -- CP-element group 602 transition  input  output  no-bypass 
    -- predecessors 601 
    -- successors 603 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_add_indices/final_index_req
      -- 
    scale_rename_ack_6091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_927_index_0_rename_ack_0, ack => cp_elements(602)); -- 
    final_index_req_6095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(602), ack => array_obj_ref_927_offset_inst_req_0); -- 
    -- CP-element group 603 transition  input  output  no-bypass 
    -- predecessors 602 
    -- successors 604 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_6096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_927_offset_inst_ack_0, ack => cp_elements(603)); -- 
    sum_rename_req_6100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(603), ack => array_obj_ref_927_root_address_inst_req_0); -- 
    -- CP-element group 604 transition  input  no-bypass 
    -- predecessors 603 
    -- successors 600 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_927_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_6101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_927_root_address_inst_ack_0, ack => cp_elements(604)); -- 
    -- CP-element group 605 transition  input  output  no-bypass 
    -- predecessors 600 
    -- successors 606 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_929_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_929_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_929_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_928_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_931_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_931_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_931_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_6106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_928_final_reg_ack_0, ack => cp_elements(605)); -- 
    base_resize_req_6123_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(605), ack => ptr_deref_932_base_resize_req_0); -- 
    -- CP-element group 606 transition  input  output  no-bypass 
    -- predecessors 605 
    -- successors 607 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6124_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_base_resize_ack_0, ack => cp_elements(606)); -- 
    sum_rename_req_6128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(606), ack => ptr_deref_932_root_address_inst_req_0); -- 
    -- CP-element group 607 transition  input  output  no-bypass 
    -- predecessors 606 
    -- successors 608 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_root_address_inst_ack_0, ack => cp_elements(607)); -- 
    root_register_req_6133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(607), ack => ptr_deref_932_addr_0_req_0); -- 
    -- CP-element group 608 transition  input  output  no-bypass 
    -- predecessors 607 
    -- successors 609 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/word_access_0/rr
      -- 
    root_register_ack_6134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_addr_0_ack_0, ack => cp_elements(608)); -- 
    rr_6144_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(608), ack => ptr_deref_932_load_0_req_0); -- 
    -- CP-element group 609 transition  input  output  no-bypass 
    -- predecessors 608 
    -- successors 610 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/word_access_0/cr
      -- 
    ra_6145_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_load_0_ack_0, ack => cp_elements(609)); -- 
    cr_6155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(609), ack => ptr_deref_932_load_0_req_1); -- 
    -- CP-element group 610 transition  input  output  no-bypass 
    -- predecessors 609 
    -- successors 611 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/merge_req
      -- 
    ca_6156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_load_0_ack_1, ack => cp_elements(610)); -- 
    merge_req_6157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(610), ack => ptr_deref_932_gather_scatter_req_0); -- 
    -- CP-element group 611 transition  input  no-bypass 
    -- predecessors 610 
    -- successors 612 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_933_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_933_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_933_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_932_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_936_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_936_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_936_completed_
      -- 
    merge_ack_6158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_932_gather_scatter_ack_0, ack => cp_elements(611)); -- 
    -- CP-element group 612 join  fork  transition  bypass 
    -- predecessors 589 611 
    -- successors 615 616 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_trigger_
      -- 
    cpelement_group_612 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(589);
      predecessors(1) <= cp_elements(611);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(612)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(612),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 613 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_active_
      -- 
    cp_elements(613) <= cp_elements(41);
    -- CP-element group 614 join  transition  bypass 
    -- predecessors 617 618 
    -- successors 619 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_938_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_938_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_938_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_942_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_942_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_941_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_941_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_941_completed_
      -- 
    cpelement_group_614 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(617);
      predecessors(1) <= cp_elements(618);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(614)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(614),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 615 transition  output  bypass 
    -- predecessors 612 
    -- successors 617 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Sample/rr
      -- 
    cp_elements(615) <= cp_elements(612);
    rr_6178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(615), ack => binary_937_inst_req_0); -- 
    -- CP-element group 616 transition  output  bypass 
    -- predecessors 612 
    -- successors 618 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Update/cr
      -- 
    cp_elements(616) <= cp_elements(612);
    cr_6183_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(616), ack => binary_937_inst_req_1); -- 
    -- CP-element group 617 transition  input  no-bypass 
    -- predecessors 615 
    -- successors 614 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Sample/ra
      -- 
    ra_6179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_937_inst_ack_0, ack => cp_elements(617)); -- 
    -- CP-element group 618 transition  input  no-bypass 
    -- predecessors 616 
    -- successors 614 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_937_Update/ca
      -- 
    ca_6184_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_937_inst_ack_1, ack => cp_elements(618)); -- 
    -- CP-element group 619 join  transition  output  bypass 
    -- predecessors 614 623 
    -- successors 624 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/split_req
      -- 
    cpelement_group_619 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(614);
      predecessors(1) <= cp_elements(623);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(619)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(619),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(619), ack => ptr_deref_940_gather_scatter_req_0); -- 
    -- CP-element group 620 transition  output  bypass 
    -- predecessors 41 
    -- successors 621 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_939_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_939_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_939_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_addr_resize/base_resize_req
      -- 
    cp_elements(620) <= cp_elements(41);
    base_resize_req_6204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(620), ack => ptr_deref_940_base_resize_req_0); -- 
    -- CP-element group 621 transition  input  output  no-bypass 
    -- predecessors 620 
    -- successors 622 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6205_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_base_resize_ack_0, ack => cp_elements(621)); -- 
    sum_rename_req_6209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => ptr_deref_940_root_address_inst_req_0); -- 
    -- CP-element group 622 transition  input  output  no-bypass 
    -- predecessors 621 
    -- successors 623 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_root_address_inst_ack_0, ack => cp_elements(622)); -- 
    root_register_req_6214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(622), ack => ptr_deref_940_addr_0_req_0); -- 
    -- CP-element group 623 transition  input  no-bypass 
    -- predecessors 622 
    -- successors 619 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_word_addrgen/root_register_ack
      -- 
    root_register_ack_6215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_addr_0_ack_0, ack => cp_elements(623)); -- 
    -- CP-element group 624 transition  input  output  no-bypass 
    -- predecessors 619 
    -- successors 625 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/word_access_0/rr
      -- 
    split_ack_6220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_gather_scatter_ack_0, ack => cp_elements(624)); -- 
    rr_6227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(624), ack => ptr_deref_940_store_0_req_0); -- 
    -- CP-element group 625 fork  transition  input  no-bypass 
    -- predecessors 624 
    -- successors 626 879 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_request/word_access/word_access_0/ra
      -- 
    ra_6228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_store_0_ack_0, ack => cp_elements(625)); -- 
    -- CP-element group 626 transition  output  bypass 
    -- predecessors 625 
    -- successors 627 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/word_access_0/cr
      -- 
    cp_elements(626) <= cp_elements(625);
    cr_6238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(626), ack => ptr_deref_940_store_0_req_1); -- 
    -- CP-element group 627 transition  input  no-bypass 
    -- predecessors 626 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_942_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_940_complete/word_access/word_access_0/ca
      -- 
    ca_6239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_940_store_0_ack_1, ack => cp_elements(627)); -- 
    -- CP-element group 628 join  transition  output  bypass 
    -- predecessors 207 632 
    -- successors 633 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/word_access_0/rr
      -- 
    cpelement_group_628 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(207);
      predecessors(1) <= cp_elements(632);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(628)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(628),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(628), ack => ptr_deref_945_load_0_req_0); -- 
    -- CP-element group 629 transition  output  bypass 
    -- predecessors 41 
    -- successors 630 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_944_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_944_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_944_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_addr_resize/base_resize_req
      -- 
    cp_elements(629) <= cp_elements(41);
    base_resize_req_6256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(629), ack => ptr_deref_945_base_resize_req_0); -- 
    -- CP-element group 630 transition  input  output  no-bypass 
    -- predecessors 629 
    -- successors 631 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_base_resize_ack_0, ack => cp_elements(630)); -- 
    sum_rename_req_6261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => ptr_deref_945_root_address_inst_req_0); -- 
    -- CP-element group 631 transition  input  output  no-bypass 
    -- predecessors 630 
    -- successors 632 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_root_address_inst_ack_0, ack => cp_elements(631)); -- 
    root_register_req_6266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(631), ack => ptr_deref_945_addr_0_req_0); -- 
    -- CP-element group 632 transition  input  no-bypass 
    -- predecessors 631 
    -- successors 628 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_word_addrgen/root_register_ack
      -- 
    root_register_ack_6267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_addr_0_ack_0, ack => cp_elements(632)); -- 
    -- CP-element group 633 transition  input  output  no-bypass 
    -- predecessors 628 
    -- successors 634 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/word_access_0/cr
      -- 
    ra_6278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_load_0_ack_0, ack => cp_elements(633)); -- 
    cr_6288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(633), ack => ptr_deref_945_load_0_req_1); -- 
    -- CP-element group 634 transition  input  output  no-bypass 
    -- predecessors 633 
    -- successors 635 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/merge_req
      -- 
    ca_6289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_load_0_ack_1, ack => cp_elements(634)); -- 
    merge_req_6290_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(634), ack => ptr_deref_945_gather_scatter_req_0); -- 
    -- CP-element group 635 transition  input  output  no-bypass 
    -- predecessors 634 
    -- successors 636 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_946_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_946_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_946_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_945_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_948_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_948_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_948_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_complete/req
      -- 
    merge_ack_6291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_945_gather_scatter_ack_0, ack => cp_elements(635)); -- 
    req_6304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(635), ack => type_cast_949_inst_req_0); -- 
    -- CP-element group 636 transition  input  output  no-bypass 
    -- predecessors 635 
    -- successors 639 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_950_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_950_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_950_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_949_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_952_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_952_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_952_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_resize_0/index_resize_req
      -- 
    ack_6305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_949_inst_ack_0, ack => cp_elements(636)); -- 
    index_resize_req_6323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => array_obj_ref_953_index_0_resize_req_0); -- 
    -- CP-element group 637 transition  bypass 
    -- predecessors 41 
    -- successors 638 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_trigger_
      -- 
    cp_elements(637) <= cp_elements(41);
    -- CP-element group 638 join  transition  output  no-bypass 
    -- predecessors 637 642 
    -- successors 643 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_complete/final_reg_req
      -- 
    cpelement_group_638 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(637);
      predecessors(1) <= cp_elements(642);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(638)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(638),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(638), ack => addr_of_954_final_reg_req_0); -- 
    -- CP-element group 639 transition  input  output  no-bypass 
    -- predecessors 636 
    -- successors 640 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_6324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_953_index_0_resize_ack_0, ack => cp_elements(639)); -- 
    scale_rename_req_6328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => array_obj_ref_953_index_0_rename_req_0); -- 
    -- CP-element group 640 transition  input  output  no-bypass 
    -- predecessors 639 
    -- successors 641 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_add_indices/final_index_req
      -- 
    scale_rename_ack_6329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_953_index_0_rename_ack_0, ack => cp_elements(640)); -- 
    final_index_req_6333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => array_obj_ref_953_offset_inst_req_0); -- 
    -- CP-element group 641 transition  input  output  no-bypass 
    -- predecessors 640 
    -- successors 642 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_6334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_953_offset_inst_ack_0, ack => cp_elements(641)); -- 
    sum_rename_req_6338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(641), ack => array_obj_ref_953_root_address_inst_req_0); -- 
    -- CP-element group 642 transition  input  no-bypass 
    -- predecessors 641 
    -- successors 638 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_953_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_6339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_953_root_address_inst_ack_0, ack => cp_elements(642)); -- 
    -- CP-element group 643 transition  input  output  no-bypass 
    -- predecessors 638 
    -- successors 644 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_955_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_955_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_955_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_954_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_957_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_957_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_957_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_6344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_954_final_reg_ack_0, ack => cp_elements(643)); -- 
    base_resize_req_6361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => ptr_deref_958_base_resize_req_0); -- 
    -- CP-element group 644 transition  input  output  no-bypass 
    -- predecessors 643 
    -- successors 645 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_base_resize_ack_0, ack => cp_elements(644)); -- 
    sum_rename_req_6366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(644), ack => ptr_deref_958_root_address_inst_req_0); -- 
    -- CP-element group 645 transition  input  output  no-bypass 
    -- predecessors 644 
    -- successors 646 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_root_address_inst_ack_0, ack => cp_elements(645)); -- 
    root_register_req_6371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => ptr_deref_958_addr_0_req_0); -- 
    -- CP-element group 646 transition  input  output  no-bypass 
    -- predecessors 645 
    -- successors 647 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/word_access_0/rr
      -- 
    root_register_ack_6372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_addr_0_ack_0, ack => cp_elements(646)); -- 
    rr_6382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(646), ack => ptr_deref_958_load_0_req_0); -- 
    -- CP-element group 647 transition  input  output  no-bypass 
    -- predecessors 646 
    -- successors 648 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/word_access_0/cr
      -- 
    ra_6383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_load_0_ack_0, ack => cp_elements(647)); -- 
    cr_6393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(647), ack => ptr_deref_958_load_0_req_1); -- 
    -- CP-element group 648 transition  input  output  no-bypass 
    -- predecessors 647 
    -- successors 649 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/merge_req
      -- 
    ca_6394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_load_0_ack_1, ack => cp_elements(648)); -- 
    merge_req_6395_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(648), ack => ptr_deref_958_gather_scatter_req_0); -- 
    -- CP-element group 649 transition  input  no-bypass 
    -- predecessors 648 
    -- successors 672 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_959_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_959_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_959_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_958_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_978_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_978_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_978_completed_
      -- 
    merge_ack_6396_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_958_gather_scatter_ack_0, ack => cp_elements(649)); -- 
    -- CP-element group 650 join  transition  output  bypass 
    -- predecessors 207 654 
    -- successors 655 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/word_access_0/rr
      -- 
    cpelement_group_650 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(207);
      predecessors(1) <= cp_elements(654);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(650)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(650),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(650), ack => ptr_deref_962_load_0_req_0); -- 
    -- CP-element group 651 transition  output  bypass 
    -- predecessors 41 
    -- successors 652 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_961_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_961_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_961_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_addr_resize/base_resize_req
      -- 
    cp_elements(651) <= cp_elements(41);
    base_resize_req_6413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(651), ack => ptr_deref_962_base_resize_req_0); -- 
    -- CP-element group 652 transition  input  output  no-bypass 
    -- predecessors 651 
    -- successors 653 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_base_resize_ack_0, ack => cp_elements(652)); -- 
    sum_rename_req_6418_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_962_root_address_inst_req_0); -- 
    -- CP-element group 653 transition  input  output  no-bypass 
    -- predecessors 652 
    -- successors 654 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6419_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_root_address_inst_ack_0, ack => cp_elements(653)); -- 
    root_register_req_6423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(653), ack => ptr_deref_962_addr_0_req_0); -- 
    -- CP-element group 654 transition  input  no-bypass 
    -- predecessors 653 
    -- successors 650 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_word_addrgen/root_register_ack
      -- 
    root_register_ack_6424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_addr_0_ack_0, ack => cp_elements(654)); -- 
    -- CP-element group 655 transition  input  output  no-bypass 
    -- predecessors 650 
    -- successors 656 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/word_access_0/cr
      -- 
    ra_6435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_load_0_ack_0, ack => cp_elements(655)); -- 
    cr_6445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => ptr_deref_962_load_0_req_1); -- 
    -- CP-element group 656 transition  input  output  no-bypass 
    -- predecessors 655 
    -- successors 657 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/merge_req
      -- 
    ca_6446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_load_0_ack_1, ack => cp_elements(656)); -- 
    merge_req_6447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => ptr_deref_962_gather_scatter_req_0); -- 
    -- CP-element group 657 transition  input  output  no-bypass 
    -- predecessors 656 
    -- successors 658 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_963_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_963_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_963_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_962_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_965_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_965_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_965_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_complete/req
      -- 
    merge_ack_6448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_962_gather_scatter_ack_0, ack => cp_elements(657)); -- 
    req_6461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(657), ack => type_cast_966_inst_req_0); -- 
    -- CP-element group 658 transition  input  output  no-bypass 
    -- predecessors 657 
    -- successors 661 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_967_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_967_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_967_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_966_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_969_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_969_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_969_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_resize_0/index_resize_req
      -- 
    ack_6462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_966_inst_ack_0, ack => cp_elements(658)); -- 
    index_resize_req_6480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => array_obj_ref_970_index_0_resize_req_0); -- 
    -- CP-element group 659 transition  bypass 
    -- predecessors 41 
    -- successors 660 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_trigger_
      -- 
    cp_elements(659) <= cp_elements(41);
    -- CP-element group 660 join  transition  output  no-bypass 
    -- predecessors 659 664 
    -- successors 665 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_complete/final_reg_req
      -- 
    cpelement_group_660 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(659);
      predecessors(1) <= cp_elements(664);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(660)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(660),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => addr_of_971_final_reg_req_0); -- 
    -- CP-element group 661 transition  input  output  no-bypass 
    -- predecessors 658 
    -- successors 662 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_6481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_970_index_0_resize_ack_0, ack => cp_elements(661)); -- 
    scale_rename_req_6485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(661), ack => array_obj_ref_970_index_0_rename_req_0); -- 
    -- CP-element group 662 transition  input  output  no-bypass 
    -- predecessors 661 
    -- successors 663 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_add_indices/final_index_req
      -- 
    scale_rename_ack_6486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_970_index_0_rename_ack_0, ack => cp_elements(662)); -- 
    final_index_req_6490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(662), ack => array_obj_ref_970_offset_inst_req_0); -- 
    -- CP-element group 663 transition  input  output  no-bypass 
    -- predecessors 662 
    -- successors 664 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_6491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_970_offset_inst_ack_0, ack => cp_elements(663)); -- 
    sum_rename_req_6495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => array_obj_ref_970_root_address_inst_req_0); -- 
    -- CP-element group 664 transition  input  no-bypass 
    -- predecessors 663 
    -- successors 660 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_970_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_6496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_970_root_address_inst_ack_0, ack => cp_elements(664)); -- 
    -- CP-element group 665 transition  input  output  no-bypass 
    -- predecessors 660 
    -- successors 666 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_972_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_972_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_972_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_971_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_974_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_974_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_974_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_6501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_971_final_reg_ack_0, ack => cp_elements(665)); -- 
    base_resize_req_6518_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(665), ack => ptr_deref_975_base_resize_req_0); -- 
    -- CP-element group 666 transition  input  output  no-bypass 
    -- predecessors 665 
    -- successors 667 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6519_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_base_resize_ack_0, ack => cp_elements(666)); -- 
    sum_rename_req_6523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(666), ack => ptr_deref_975_root_address_inst_req_0); -- 
    -- CP-element group 667 transition  input  output  no-bypass 
    -- predecessors 666 
    -- successors 668 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_root_address_inst_ack_0, ack => cp_elements(667)); -- 
    root_register_req_6528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(667), ack => ptr_deref_975_addr_0_req_0); -- 
    -- CP-element group 668 transition  input  output  no-bypass 
    -- predecessors 667 
    -- successors 669 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/word_access_0/rr
      -- 
    root_register_ack_6529_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_addr_0_ack_0, ack => cp_elements(668)); -- 
    rr_6539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => ptr_deref_975_load_0_req_0); -- 
    -- CP-element group 669 transition  input  output  no-bypass 
    -- predecessors 668 
    -- successors 670 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/word_access_0/cr
      -- 
    ra_6540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_load_0_ack_0, ack => cp_elements(669)); -- 
    cr_6550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(669), ack => ptr_deref_975_load_0_req_1); -- 
    -- CP-element group 670 transition  input  output  no-bypass 
    -- predecessors 669 
    -- successors 671 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/merge_req
      -- 
    ca_6551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_load_0_ack_1, ack => cp_elements(670)); -- 
    merge_req_6552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(670), ack => ptr_deref_975_gather_scatter_req_0); -- 
    -- CP-element group 671 transition  input  no-bypass 
    -- predecessors 670 
    -- successors 672 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_976_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_976_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_976_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_975_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_979_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_979_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_979_completed_
      -- 
    merge_ack_6553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_975_gather_scatter_ack_0, ack => cp_elements(671)); -- 
    -- CP-element group 672 join  fork  transition  bypass 
    -- predecessors 649 671 
    -- successors 675 676 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_trigger_
      -- 
    cpelement_group_672 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(649);
      predecessors(1) <= cp_elements(671);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(672)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(672),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 673 transition  bypass 
    -- predecessors 41 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_active_
      -- 
    cp_elements(673) <= cp_elements(41);
    -- CP-element group 674 join  transition  bypass 
    -- predecessors 677 678 
    -- successors 679 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_981_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_981_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_981_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_985_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_985_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_984_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_984_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_984_completed_
      -- 
    cpelement_group_674 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(677);
      predecessors(1) <= cp_elements(678);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(674)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(674),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 675 transition  output  bypass 
    -- predecessors 672 
    -- successors 677 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Sample/rr
      -- 
    cp_elements(675) <= cp_elements(672);
    rr_6573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(675), ack => binary_980_inst_req_0); -- 
    -- CP-element group 676 transition  output  bypass 
    -- predecessors 672 
    -- successors 678 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_update_start_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Update/cr
      -- 
    cp_elements(676) <= cp_elements(672);
    cr_6578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(676), ack => binary_980_inst_req_1); -- 
    -- CP-element group 677 transition  input  no-bypass 
    -- predecessors 675 
    -- successors 674 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Sample/ra
      -- 
    ra_6574_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_980_inst_ack_0, ack => cp_elements(677)); -- 
    -- CP-element group 678 transition  input  no-bypass 
    -- predecessors 676 
    -- successors 674 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/binary_980_Update/ca
      -- 
    ca_6579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_980_inst_ack_1, ack => cp_elements(678)); -- 
    -- CP-element group 679 join  transition  output  bypass 
    -- predecessors 674 683 
    -- successors 684 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/split_req
      -- 
    cpelement_group_679 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(674);
      predecessors(1) <= cp_elements(683);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(679)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(679),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(679), ack => ptr_deref_983_gather_scatter_req_0); -- 
    -- CP-element group 680 transition  output  bypass 
    -- predecessors 41 
    -- successors 681 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_982_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_982_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_982_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_addr_resize/base_resize_req
      -- 
    cp_elements(680) <= cp_elements(41);
    base_resize_req_6599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => ptr_deref_983_base_resize_req_0); -- 
    -- CP-element group 681 transition  input  output  no-bypass 
    -- predecessors 680 
    -- successors 682 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_base_resize_ack_0, ack => cp_elements(681)); -- 
    sum_rename_req_6604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(681), ack => ptr_deref_983_root_address_inst_req_0); -- 
    -- CP-element group 682 transition  input  output  no-bypass 
    -- predecessors 681 
    -- successors 683 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_root_address_inst_ack_0, ack => cp_elements(682)); -- 
    root_register_req_6609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => ptr_deref_983_addr_0_req_0); -- 
    -- CP-element group 683 transition  input  no-bypass 
    -- predecessors 682 
    -- successors 679 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_word_addrgen/root_register_ack
      -- 
    root_register_ack_6610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_addr_0_ack_0, ack => cp_elements(683)); -- 
    -- CP-element group 684 transition  input  output  no-bypass 
    -- predecessors 679 
    -- successors 685 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/word_access_0/rr
      -- 
    split_ack_6615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_gather_scatter_ack_0, ack => cp_elements(684)); -- 
    rr_6622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_983_store_0_req_0); -- 
    -- CP-element group 685 fork  transition  input  no-bypass 
    -- predecessors 684 
    -- successors 686 911 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_request/word_access/word_access_0/ra
      -- 
    ra_6623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_store_0_ack_0, ack => cp_elements(685)); -- 
    -- CP-element group 686 transition  output  bypass 
    -- predecessors 685 
    -- successors 687 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/word_access_0/cr
      -- 
    cp_elements(686) <= cp_elements(685);
    cr_6633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => ptr_deref_983_store_0_req_1); -- 
    -- CP-element group 687 transition  input  no-bypass 
    -- predecessors 686 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_985_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_983_complete/word_access/word_access_0/ca
      -- 
    ca_6634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_983_store_0_ack_1, ack => cp_elements(687)); -- 
    -- CP-element group 688 join  transition  output  bypass 
    -- predecessors 265 692 
    -- successors 693 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/word_access_0/rr
      -- 
    cpelement_group_688 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(265);
      predecessors(1) <= cp_elements(692);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(688)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(688), ack => ptr_deref_988_load_0_req_0); -- 
    -- CP-element group 689 transition  output  bypass 
    -- predecessors 41 
    -- successors 690 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_987_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_987_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_987_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_addr_resize/base_resize_req
      -- 
    cp_elements(689) <= cp_elements(41);
    base_resize_req_6651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(689), ack => ptr_deref_988_base_resize_req_0); -- 
    -- CP-element group 690 transition  input  output  no-bypass 
    -- predecessors 689 
    -- successors 691 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_base_resize_ack_0, ack => cp_elements(690)); -- 
    sum_rename_req_6656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => ptr_deref_988_root_address_inst_req_0); -- 
    -- CP-element group 691 transition  input  output  no-bypass 
    -- predecessors 690 
    -- successors 692 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_root_address_inst_ack_0, ack => cp_elements(691)); -- 
    root_register_req_6661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(691), ack => ptr_deref_988_addr_0_req_0); -- 
    -- CP-element group 692 transition  input  no-bypass 
    -- predecessors 691 
    -- successors 688 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_word_addrgen/root_register_ack
      -- 
    root_register_ack_6662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_addr_0_ack_0, ack => cp_elements(692)); -- 
    -- CP-element group 693 transition  input  output  no-bypass 
    -- predecessors 688 
    -- successors 694 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/$entry
      -- 
    ra_6673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_load_0_ack_0, ack => cp_elements(693)); -- 
    cr_6683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => ptr_deref_988_load_0_req_1); -- 
    -- CP-element group 694 transition  input  output  no-bypass 
    -- predecessors 693 
    -- successors 695 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/merge_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/word_access/$exit
      -- 
    ca_6684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_load_0_ack_1, ack => cp_elements(694)); -- 
    merge_req_6685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => ptr_deref_988_gather_scatter_req_0); -- 
    -- CP-element group 695 transition  input  no-bypass 
    -- predecessors 694 
    -- successors 711 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_989_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_989_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_989_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_988_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1006_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1006_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1005_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1005_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1005_completed_
      -- 
    merge_ack_6686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_988_gather_scatter_ack_0, ack => cp_elements(695)); -- 
    -- CP-element group 696 transition  output  bypass 
    -- predecessors 41 
    -- successors 697 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_991_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_991_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_991_completed_
      -- 
    cp_elements(696) <= cp_elements(41);
    base_resize_req_6703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(696), ack => ptr_deref_992_base_resize_req_0); -- 
    -- CP-element group 697 transition  input  output  no-bypass 
    -- predecessors 696 
    -- successors 698 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_base_resize_ack_0, ack => cp_elements(697)); -- 
    sum_rename_req_6708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => ptr_deref_992_root_address_inst_req_0); -- 
    -- CP-element group 698 transition  input  output  no-bypass 
    -- predecessors 697 
    -- successors 699 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_root_address_inst_ack_0, ack => cp_elements(698)); -- 
    root_register_req_6713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(698), ack => ptr_deref_992_addr_0_req_0); -- 
    -- CP-element group 699 transition  input  output  no-bypass 
    -- predecessors 698 
    -- successors 700 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/word_access_0/rr
      -- 
    root_register_ack_6714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_addr_0_ack_0, ack => cp_elements(699)); -- 
    rr_6724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_992_load_0_req_0); -- 
    -- CP-element group 700 transition  input  output  no-bypass 
    -- predecessors 699 
    -- successors 701 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/word_access_0/cr
      -- 
    ra_6725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_load_0_ack_0, ack => cp_elements(700)); -- 
    cr_6735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(700), ack => ptr_deref_992_load_0_req_1); -- 
    -- CP-element group 701 transition  input  output  no-bypass 
    -- predecessors 700 
    -- successors 702 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/merge_req
      -- 
    ca_6736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_load_0_ack_1, ack => cp_elements(701)); -- 
    merge_req_6737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_992_gather_scatter_req_0); -- 
    -- CP-element group 702 transition  input  output  no-bypass 
    -- predecessors 701 
    -- successors 703 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_993_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_993_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_993_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_992_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_995_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_995_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_995_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_complete/req
      -- 
    merge_ack_6738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_992_gather_scatter_ack_0, ack => cp_elements(702)); -- 
    req_6751_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => type_cast_996_inst_req_0); -- 
    -- CP-element group 703 transition  input  output  no-bypass 
    -- predecessors 702 
    -- successors 706 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_997_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_997_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_997_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_996_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_999_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_999_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_999_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_resize_0/index_resize_req
      -- 
    ack_6752_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_996_inst_ack_0, ack => cp_elements(703)); -- 
    index_resize_req_6770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(703), ack => array_obj_ref_1000_index_0_resize_req_0); -- 
    -- CP-element group 704 transition  bypass 
    -- predecessors 41 
    -- successors 705 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_trigger_
      -- 
    cp_elements(704) <= cp_elements(41);
    -- CP-element group 705 join  transition  output  no-bypass 
    -- predecessors 704 709 
    -- successors 710 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_complete/final_reg_req
      -- 
    cpelement_group_705 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(704);
      predecessors(1) <= cp_elements(709);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(705)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(705),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => addr_of_1001_final_reg_req_0); -- 
    -- CP-element group 706 transition  input  output  no-bypass 
    -- predecessors 703 
    -- successors 707 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_6771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1000_index_0_resize_ack_0, ack => cp_elements(706)); -- 
    scale_rename_req_6775_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(706), ack => array_obj_ref_1000_index_0_rename_req_0); -- 
    -- CP-element group 707 transition  input  output  no-bypass 
    -- predecessors 706 
    -- successors 708 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_add_indices/final_index_req
      -- 
    scale_rename_ack_6776_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1000_index_0_rename_ack_0, ack => cp_elements(707)); -- 
    final_index_req_6780_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => array_obj_ref_1000_offset_inst_req_0); -- 
    -- CP-element group 708 transition  input  output  no-bypass 
    -- predecessors 707 
    -- successors 709 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_6781_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1000_offset_inst_ack_0, ack => cp_elements(708)); -- 
    sum_rename_req_6785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => array_obj_ref_1000_root_address_inst_req_0); -- 
    -- CP-element group 709 transition  input  no-bypass 
    -- predecessors 708 
    -- successors 705 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1000_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_6786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1000_root_address_inst_ack_0, ack => cp_elements(709)); -- 
    -- CP-element group 710 transition  input  output  no-bypass 
    -- predecessors 705 
    -- successors 712 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1002_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1002_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1002_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1001_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1003_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1003_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1003_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_6791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1001_final_reg_ack_0, ack => cp_elements(710)); -- 
    base_resize_req_6811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => ptr_deref_1004_base_resize_req_0); -- 
    -- CP-element group 711 join  transition  output  bypass 
    -- predecessors 695 714 
    -- successors 715 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/split_req
      -- 
    cpelement_group_711 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(695);
      predecessors(1) <= cp_elements(714);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(711)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(711),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => ptr_deref_1004_gather_scatter_req_0); -- 
    -- CP-element group 712 transition  input  output  no-bypass 
    -- predecessors 710 
    -- successors 713 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_base_resize_ack_0, ack => cp_elements(712)); -- 
    sum_rename_req_6816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(712), ack => ptr_deref_1004_root_address_inst_req_0); -- 
    -- CP-element group 713 transition  input  output  no-bypass 
    -- predecessors 712 
    -- successors 714 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_root_address_inst_ack_0, ack => cp_elements(713)); -- 
    root_register_req_6821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(713), ack => ptr_deref_1004_addr_0_req_0); -- 
    -- CP-element group 714 transition  input  no-bypass 
    -- predecessors 713 
    -- successors 711 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_word_addrgen/root_register_ack
      -- 
    root_register_ack_6822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_addr_0_ack_0, ack => cp_elements(714)); -- 
    -- CP-element group 715 transition  input  output  no-bypass 
    -- predecessors 711 
    -- successors 716 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/word_access_0/rr
      -- 
    split_ack_6827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_gather_scatter_ack_0, ack => cp_elements(715)); -- 
    rr_6834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(715), ack => ptr_deref_1004_store_0_req_0); -- 
    -- CP-element group 716 fork  transition  input  no-bypass 
    -- predecessors 715 
    -- successors 717 743 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_request/word_access/word_access_0/ra
      -- 
    ra_6835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_store_0_ack_0, ack => cp_elements(716)); -- 
    -- CP-element group 717 transition  output  bypass 
    -- predecessors 716 
    -- successors 718 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/word_access_0/cr
      -- 
    cp_elements(717) <= cp_elements(716);
    cr_6845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(717), ack => ptr_deref_1004_store_0_req_1); -- 
    -- CP-element group 718 transition  input  no-bypass 
    -- predecessors 717 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1006_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1004_complete/word_access/word_access_0/ca
      -- 
    ca_6846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1004_store_0_ack_1, ack => cp_elements(718)); -- 
    -- CP-element group 719 join  transition  output  bypass 
    -- predecessors 325 723 
    -- successors 724 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/word_access_0/rr
      -- 
    cpelement_group_719 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(325);
      predecessors(1) <= cp_elements(723);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(719)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(719),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(719), ack => ptr_deref_1009_load_0_req_0); -- 
    -- CP-element group 720 transition  output  bypass 
    -- predecessors 41 
    -- successors 721 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1008_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1008_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1008_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_addr_resize/base_resize_req
      -- 
    cp_elements(720) <= cp_elements(41);
    base_resize_req_6863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => ptr_deref_1009_base_resize_req_0); -- 
    -- CP-element group 721 transition  input  output  no-bypass 
    -- predecessors 720 
    -- successors 722 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_base_resize_ack_0, ack => cp_elements(721)); -- 
    sum_rename_req_6868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(721), ack => ptr_deref_1009_root_address_inst_req_0); -- 
    -- CP-element group 722 transition  input  output  no-bypass 
    -- predecessors 721 
    -- successors 723 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_root_address_inst_ack_0, ack => cp_elements(722)); -- 
    root_register_req_6873_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(722), ack => ptr_deref_1009_addr_0_req_0); -- 
    -- CP-element group 723 transition  input  no-bypass 
    -- predecessors 722 
    -- successors 719 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_word_addrgen/root_register_ack
      -- 
    root_register_ack_6874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_addr_0_ack_0, ack => cp_elements(723)); -- 
    -- CP-element group 724 transition  input  output  no-bypass 
    -- predecessors 719 
    -- successors 725 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/word_access_0/cr
      -- 
    ra_6885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_load_0_ack_0, ack => cp_elements(724)); -- 
    cr_6895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(724), ack => ptr_deref_1009_load_0_req_1); -- 
    -- CP-element group 725 transition  input  output  no-bypass 
    -- predecessors 724 
    -- successors 726 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/merge_req
      -- 
    ca_6896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_load_0_ack_1, ack => cp_elements(725)); -- 
    merge_req_6897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => ptr_deref_1009_gather_scatter_req_0); -- 
    -- CP-element group 726 transition  input  no-bypass 
    -- predecessors 725 
    -- successors 743 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1010_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1010_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1010_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1009_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1027_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1027_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1026_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1026_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1026_completed_
      -- 
    merge_ack_6898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1009_gather_scatter_ack_0, ack => cp_elements(726)); -- 
    -- CP-element group 727 join  transition  output  bypass 
    -- predecessors 63 731 
    -- successors 732 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/word_access_0/rr
      -- 
    cpelement_group_727 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(63);
      predecessors(1) <= cp_elements(731);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(727)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(727),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => ptr_deref_1013_load_0_req_0); -- 
    -- CP-element group 728 transition  output  bypass 
    -- predecessors 41 
    -- successors 729 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1012_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1012_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1012_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_addr_resize/base_resize_req
      -- 
    cp_elements(728) <= cp_elements(41);
    base_resize_req_6915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => ptr_deref_1013_base_resize_req_0); -- 
    -- CP-element group 729 transition  input  output  no-bypass 
    -- predecessors 728 
    -- successors 730 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_6916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_base_resize_ack_0, ack => cp_elements(729)); -- 
    sum_rename_req_6920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => ptr_deref_1013_root_address_inst_req_0); -- 
    -- CP-element group 730 transition  input  output  no-bypass 
    -- predecessors 729 
    -- successors 731 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_word_addrgen/root_register_req
      -- 
    sum_rename_ack_6921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_root_address_inst_ack_0, ack => cp_elements(730)); -- 
    root_register_req_6925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(730), ack => ptr_deref_1013_addr_0_req_0); -- 
    -- CP-element group 731 transition  input  no-bypass 
    -- predecessors 730 
    -- successors 727 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_word_addrgen/root_register_ack
      -- 
    root_register_ack_6926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_addr_0_ack_0, ack => cp_elements(731)); -- 
    -- CP-element group 732 transition  input  output  no-bypass 
    -- predecessors 727 
    -- successors 733 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/word_access_0/cr
      -- 
    ra_6937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_load_0_ack_0, ack => cp_elements(732)); -- 
    cr_6947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => ptr_deref_1013_load_0_req_1); -- 
    -- CP-element group 733 transition  input  output  no-bypass 
    -- predecessors 732 
    -- successors 734 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/merge_req
      -- 
    ca_6948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_load_0_ack_1, ack => cp_elements(733)); -- 
    merge_req_6949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(733), ack => ptr_deref_1013_gather_scatter_req_0); -- 
    -- CP-element group 734 transition  input  output  no-bypass 
    -- predecessors 733 
    -- successors 735 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1014_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1014_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1014_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1013_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1016_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1016_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1016_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_complete/req
      -- 
    merge_ack_6950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1013_gather_scatter_ack_0, ack => cp_elements(734)); -- 
    req_6963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => type_cast_1017_inst_req_0); -- 
    -- CP-element group 735 transition  input  output  no-bypass 
    -- predecessors 734 
    -- successors 738 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1018_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1018_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1018_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1017_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1020_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1020_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1020_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_resize_0/index_resize_req
      -- 
    ack_6964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1017_inst_ack_0, ack => cp_elements(735)); -- 
    index_resize_req_6982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => array_obj_ref_1021_index_0_resize_req_0); -- 
    -- CP-element group 736 transition  bypass 
    -- predecessors 41 
    -- successors 737 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_trigger_
      -- 
    cp_elements(736) <= cp_elements(41);
    -- CP-element group 737 join  transition  output  no-bypass 
    -- predecessors 736 741 
    -- successors 742 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_complete/final_reg_req
      -- 
    cpelement_group_737 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(736);
      predecessors(1) <= cp_elements(741);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(737)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(737),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => addr_of_1022_final_reg_req_0); -- 
    -- CP-element group 738 transition  input  output  no-bypass 
    -- predecessors 735 
    -- successors 739 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_6983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_index_0_resize_ack_0, ack => cp_elements(738)); -- 
    scale_rename_req_6987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(738), ack => array_obj_ref_1021_index_0_rename_req_0); -- 
    -- CP-element group 739 transition  input  output  no-bypass 
    -- predecessors 738 
    -- successors 740 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_add_indices/final_index_req
      -- 
    scale_rename_ack_6988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_index_0_rename_ack_0, ack => cp_elements(739)); -- 
    final_index_req_6992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => array_obj_ref_1021_offset_inst_req_0); -- 
    -- CP-element group 740 transition  input  output  no-bypass 
    -- predecessors 739 
    -- successors 741 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_6993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_offset_inst_ack_0, ack => cp_elements(740)); -- 
    sum_rename_req_6997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => array_obj_ref_1021_root_address_inst_req_0); -- 
    -- CP-element group 741 transition  input  no-bypass 
    -- predecessors 740 
    -- successors 737 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1021_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_6998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1021_root_address_inst_ack_0, ack => cp_elements(741)); -- 
    -- CP-element group 742 transition  input  output  no-bypass 
    -- predecessors 737 
    -- successors 744 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1023_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1023_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1023_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1022_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1024_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1024_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1024_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_7003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1022_final_reg_ack_0, ack => cp_elements(742)); -- 
    base_resize_req_7023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => ptr_deref_1025_base_resize_req_0); -- 
    -- CP-element group 743 join  transition  output  bypass 
    -- predecessors 716 726 746 
    -- successors 747 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/split_req
      -- 
    cpelement_group_743 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(716);
      predecessors(1) <= cp_elements(726);
      predecessors(2) <= cp_elements(746);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(743)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(743),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => ptr_deref_1025_gather_scatter_req_0); -- 
    -- CP-element group 744 transition  input  output  no-bypass 
    -- predecessors 742 
    -- successors 745 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_base_resize_ack_0, ack => cp_elements(744)); -- 
    sum_rename_req_7028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => ptr_deref_1025_root_address_inst_req_0); -- 
    -- CP-element group 745 transition  input  output  no-bypass 
    -- predecessors 744 
    -- successors 746 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_root_address_inst_ack_0, ack => cp_elements(745)); -- 
    root_register_req_7033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => ptr_deref_1025_addr_0_req_0); -- 
    -- CP-element group 746 transition  input  no-bypass 
    -- predecessors 745 
    -- successors 743 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_word_addrgen/root_register_ack
      -- 
    root_register_ack_7034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_addr_0_ack_0, ack => cp_elements(746)); -- 
    -- CP-element group 747 transition  input  output  no-bypass 
    -- predecessors 743 
    -- successors 748 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/word_access_0/rr
      -- 
    split_ack_7039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_gather_scatter_ack_0, ack => cp_elements(747)); -- 
    rr_7046_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(747), ack => ptr_deref_1025_store_0_req_0); -- 
    -- CP-element group 748 fork  transition  input  no-bypass 
    -- predecessors 747 
    -- successors 749 775 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_request/word_access/word_access_0/ra
      -- 
    ra_7047_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_store_0_ack_0, ack => cp_elements(748)); -- 
    -- CP-element group 749 transition  output  bypass 
    -- predecessors 748 
    -- successors 750 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/word_access_0/cr
      -- 
    cp_elements(749) <= cp_elements(748);
    cr_7057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => ptr_deref_1025_store_0_req_1); -- 
    -- CP-element group 750 transition  input  no-bypass 
    -- predecessors 749 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1027_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1025_complete/word_access/word_access_0/ca
      -- 
    ca_7058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1025_store_0_ack_1, ack => cp_elements(750)); -- 
    -- CP-element group 751 join  transition  output  bypass 
    -- predecessors 385 755 
    -- successors 756 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_trigger_
      -- 
    cpelement_group_751 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(385);
      predecessors(1) <= cp_elements(755);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(751)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(751),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(751), ack => ptr_deref_1030_load_0_req_0); -- 
    -- CP-element group 752 transition  output  bypass 
    -- predecessors 41 
    -- successors 753 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1029_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1029_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1029_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_address_calculated
      -- 
    cp_elements(752) <= cp_elements(41);
    base_resize_req_7075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(752), ack => ptr_deref_1030_base_resize_req_0); -- 
    -- CP-element group 753 transition  input  output  no-bypass 
    -- predecessors 752 
    -- successors 754 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_address_resized
      -- 
    base_resize_ack_7076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_base_resize_ack_0, ack => cp_elements(753)); -- 
    sum_rename_req_7080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ptr_deref_1030_root_address_inst_req_0); -- 
    -- CP-element group 754 transition  input  output  no-bypass 
    -- predecessors 753 
    -- successors 755 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_root_address_calculated
      -- 
    sum_rename_ack_7081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_root_address_inst_ack_0, ack => cp_elements(754)); -- 
    root_register_req_7085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(754), ack => ptr_deref_1030_addr_0_req_0); -- 
    -- CP-element group 755 transition  input  no-bypass 
    -- predecessors 754 
    -- successors 751 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_word_address_calculated
      -- 
    root_register_ack_7086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_addr_0_ack_0, ack => cp_elements(755)); -- 
    -- CP-element group 756 transition  input  output  no-bypass 
    -- predecessors 751 
    -- successors 757 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_active_
      -- 
    ra_7097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_load_0_ack_0, ack => cp_elements(756)); -- 
    cr_7107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => ptr_deref_1030_load_0_req_1); -- 
    -- CP-element group 757 transition  input  output  no-bypass 
    -- predecessors 756 
    -- successors 758 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/merge_req
      -- 
    ca_7108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_load_0_ack_1, ack => cp_elements(757)); -- 
    merge_req_7109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => ptr_deref_1030_gather_scatter_req_0); -- 
    -- CP-element group 758 transition  input  no-bypass 
    -- predecessors 757 
    -- successors 775 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1047_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1047_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1047_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1048_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1048_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1031_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1031_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1031_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1030_completed_
      -- 
    merge_ack_7110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1030_gather_scatter_ack_0, ack => cp_elements(758)); -- 
    -- CP-element group 759 join  transition  output  bypass 
    -- predecessors 87 763 
    -- successors 764 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/$entry
      -- 
    cpelement_group_759 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(87);
      predecessors(1) <= cp_elements(763);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(759)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(759),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => ptr_deref_1034_load_0_req_0); -- 
    -- CP-element group 760 transition  output  bypass 
    -- predecessors 41 
    -- successors 761 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1033_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1033_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1033_completed_
      -- 
    cp_elements(760) <= cp_elements(41);
    base_resize_req_7127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(760), ack => ptr_deref_1034_base_resize_req_0); -- 
    -- CP-element group 761 transition  input  output  no-bypass 
    -- predecessors 760 
    -- successors 762 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_base_resize_ack_0, ack => cp_elements(761)); -- 
    sum_rename_req_7132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => ptr_deref_1034_root_address_inst_req_0); -- 
    -- CP-element group 762 transition  input  output  no-bypass 
    -- predecessors 761 
    -- successors 763 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_root_address_inst_ack_0, ack => cp_elements(762)); -- 
    root_register_req_7137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(762), ack => ptr_deref_1034_addr_0_req_0); -- 
    -- CP-element group 763 transition  input  no-bypass 
    -- predecessors 762 
    -- successors 759 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_word_addrgen/$exit
      -- 
    root_register_ack_7138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_addr_0_ack_0, ack => cp_elements(763)); -- 
    -- CP-element group 764 transition  input  output  no-bypass 
    -- predecessors 759 
    -- successors 765 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_request/$exit
      -- 
    ra_7149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_load_0_ack_0, ack => cp_elements(764)); -- 
    cr_7159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(764), ack => ptr_deref_1034_load_0_req_1); -- 
    -- CP-element group 765 transition  input  output  no-bypass 
    -- predecessors 764 
    -- successors 766 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/merge_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/word_access/word_access_0/ca
      -- 
    ca_7160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_load_0_ack_1, ack => cp_elements(765)); -- 
    merge_req_7161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => ptr_deref_1034_gather_scatter_req_0); -- 
    -- CP-element group 766 transition  input  output  no-bypass 
    -- predecessors 765 
    -- successors 767 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1037_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1035_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1035_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1035_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1034_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1037_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_complete/req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1037_completed_
      -- 
    merge_ack_7162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1034_gather_scatter_ack_0, ack => cp_elements(766)); -- 
    req_7175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(766), ack => type_cast_1038_inst_req_0); -- 
    -- CP-element group 767 transition  input  output  no-bypass 
    -- predecessors 766 
    -- successors 770 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1041_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1041_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1039_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1039_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1041_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1039_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1038_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_resize_0/index_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_resize_0/$entry
      -- 
    ack_7176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1038_inst_ack_0, ack => cp_elements(767)); -- 
    index_resize_req_7194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => array_obj_ref_1042_index_0_resize_req_0); -- 
    -- CP-element group 768 transition  bypass 
    -- predecessors 41 
    -- successors 769 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_trigger_
      -- 
    cp_elements(768) <= cp_elements(41);
    -- CP-element group 769 join  transition  output  no-bypass 
    -- predecessors 768 773 
    -- successors 774 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_complete/final_reg_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_complete/$entry
      -- 
    cpelement_group_769 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(768);
      predecessors(1) <= cp_elements(773);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(769)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(769),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(769), ack => addr_of_1043_final_reg_req_0); -- 
    -- CP-element group 770 transition  input  output  no-bypass 
    -- predecessors 767 
    -- successors 771 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_resize_0/$exit
      -- 
    index_resize_ack_7195_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1042_index_0_resize_ack_0, ack => cp_elements(770)); -- 
    scale_rename_req_7199_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => array_obj_ref_1042_index_0_rename_req_0); -- 
    -- CP-element group 771 transition  input  output  no-bypass 
    -- predecessors 770 
    -- successors 772 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_add_indices/final_index_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_index_scale_0/$exit
      -- 
    scale_rename_ack_7200_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1042_index_0_rename_ack_0, ack => cp_elements(771)); -- 
    final_index_req_7204_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(771), ack => array_obj_ref_1042_offset_inst_req_0); -- 
    -- CP-element group 772 transition  input  output  no-bypass 
    -- predecessors 771 
    -- successors 773 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_7205_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1042_offset_inst_ack_0, ack => cp_elements(772)); -- 
    sum_rename_req_7209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => array_obj_ref_1042_root_address_inst_req_0); -- 
    -- CP-element group 773 transition  input  no-bypass 
    -- predecessors 772 
    -- successors 769 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1042_root_address_calculated
      -- 
    sum_rename_ack_7210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1042_root_address_inst_ack_0, ack => cp_elements(773)); -- 
    -- CP-element group 774 transition  input  output  no-bypass 
    -- predecessors 769 
    -- successors 776 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1044_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1045_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1045_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1044_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1044_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1045_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1043_complete/$exit
      -- 
    final_reg_ack_7215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1043_final_reg_ack_0, ack => cp_elements(774)); -- 
    base_resize_req_7235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => ptr_deref_1046_base_resize_req_0); -- 
    -- CP-element group 775 join  transition  output  bypass 
    -- predecessors 748 758 778 
    -- successors 779 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/split_req
      -- 
    cpelement_group_775 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(748);
      predecessors(1) <= cp_elements(758);
      predecessors(2) <= cp_elements(778);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(775)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(775),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(775), ack => ptr_deref_1046_gather_scatter_req_0); -- 
    -- CP-element group 776 transition  input  output  no-bypass 
    -- predecessors 774 
    -- successors 777 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_7236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_base_resize_ack_0, ack => cp_elements(776)); -- 
    sum_rename_req_7240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => ptr_deref_1046_root_address_inst_req_0); -- 
    -- CP-element group 777 transition  input  output  no-bypass 
    -- predecessors 776 
    -- successors 778 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_root_address_inst_ack_0, ack => cp_elements(777)); -- 
    root_register_req_7245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(777), ack => ptr_deref_1046_addr_0_req_0); -- 
    -- CP-element group 778 transition  input  no-bypass 
    -- predecessors 777 
    -- successors 775 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_word_addrgen/root_register_ack
      -- 
    root_register_ack_7246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_addr_0_ack_0, ack => cp_elements(778)); -- 
    -- CP-element group 779 transition  input  output  no-bypass 
    -- predecessors 775 
    -- successors 780 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/split_ack
      -- 
    split_ack_7251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_gather_scatter_ack_0, ack => cp_elements(779)); -- 
    rr_7258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(779), ack => ptr_deref_1046_store_0_req_0); -- 
    -- CP-element group 780 fork  transition  input  no-bypass 
    -- predecessors 779 
    -- successors 781 807 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_request/$exit
      -- 
    ra_7259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_store_0_ack_0, ack => cp_elements(780)); -- 
    -- CP-element group 781 transition  output  bypass 
    -- predecessors 780 
    -- successors 782 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/word_access_0/$entry
      -- 
    cp_elements(781) <= cp_elements(780);
    cr_7269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(781), ack => ptr_deref_1046_store_0_req_1); -- 
    -- CP-element group 782 transition  input  no-bypass 
    -- predecessors 781 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1048_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1046_complete/word_access/$exit
      -- 
    ca_7270_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1046_store_0_ack_1, ack => cp_elements(782)); -- 
    -- CP-element group 783 join  transition  output  bypass 
    -- predecessors 445 787 
    -- successors 788 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/$entry
      -- 
    cpelement_group_783 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(445);
      predecessors(1) <= cp_elements(787);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(783)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(783),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => ptr_deref_1051_load_0_req_0); -- 
    -- CP-element group 784 transition  output  bypass 
    -- predecessors 41 
    -- successors 785 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1050_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1050_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1050_active_
      -- 
    cp_elements(784) <= cp_elements(41);
    base_resize_req_7287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => ptr_deref_1051_base_resize_req_0); -- 
    -- CP-element group 785 transition  input  output  no-bypass 
    -- predecessors 784 
    -- successors 786 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_addr_resize/$exit
      -- 
    base_resize_ack_7288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_base_resize_ack_0, ack => cp_elements(785)); -- 
    sum_rename_req_7292_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => ptr_deref_1051_root_address_inst_req_0); -- 
    -- CP-element group 786 transition  input  output  no-bypass 
    -- predecessors 785 
    -- successors 787 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7293_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_root_address_inst_ack_0, ack => cp_elements(786)); -- 
    root_register_req_7297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(786), ack => ptr_deref_1051_addr_0_req_0); -- 
    -- CP-element group 787 transition  input  no-bypass 
    -- predecessors 786 
    -- successors 783 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_word_addrgen/$exit
      -- 
    root_register_ack_7298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_addr_0_ack_0, ack => cp_elements(787)); -- 
    -- CP-element group 788 transition  input  output  no-bypass 
    -- predecessors 783 
    -- successors 789 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_request/$exit
      -- 
    ra_7309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_load_0_ack_0, ack => cp_elements(788)); -- 
    cr_7319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => ptr_deref_1051_load_0_req_1); -- 
    -- CP-element group 789 transition  input  output  no-bypass 
    -- predecessors 788 
    -- successors 790 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/merge_req
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/word_access/word_access_0/ca
      -- 
    ca_7320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_load_0_ack_1, ack => cp_elements(789)); -- 
    merge_req_7321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(789), ack => ptr_deref_1051_gather_scatter_req_0); -- 
    -- CP-element group 790 transition  input  no-bypass 
    -- predecessors 789 
    -- successors 807 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1052_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1052_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1052_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1051_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1069_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1069_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1068_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1068_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1068_completed_
      -- 
    merge_ack_7322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1051_gather_scatter_ack_0, ack => cp_elements(790)); -- 
    -- CP-element group 791 join  transition  output  bypass 
    -- predecessors 111 795 
    -- successors 796 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/word_access_0/rr
      -- 
    cpelement_group_791 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(111);
      predecessors(1) <= cp_elements(795);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(791)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(791),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => ptr_deref_1055_load_0_req_0); -- 
    -- CP-element group 792 transition  output  bypass 
    -- predecessors 41 
    -- successors 793 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1054_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1054_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1054_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_addr_resize/base_resize_req
      -- 
    cp_elements(792) <= cp_elements(41);
    base_resize_req_7339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(792), ack => ptr_deref_1055_base_resize_req_0); -- 
    -- CP-element group 793 transition  input  output  no-bypass 
    -- predecessors 792 
    -- successors 794 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_base_resize_ack_0, ack => cp_elements(793)); -- 
    sum_rename_req_7344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => ptr_deref_1055_root_address_inst_req_0); -- 
    -- CP-element group 794 transition  input  output  no-bypass 
    -- predecessors 793 
    -- successors 795 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_root_address_inst_ack_0, ack => cp_elements(794)); -- 
    root_register_req_7349_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => ptr_deref_1055_addr_0_req_0); -- 
    -- CP-element group 795 transition  input  no-bypass 
    -- predecessors 794 
    -- successors 791 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_word_addrgen/root_register_ack
      -- 
    root_register_ack_7350_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_0_ack_0, ack => cp_elements(795)); -- 
    -- CP-element group 796 transition  input  output  no-bypass 
    -- predecessors 791 
    -- successors 797 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/word_access_0/cr
      -- 
    ra_7361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_load_0_ack_0, ack => cp_elements(796)); -- 
    cr_7371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => ptr_deref_1055_load_0_req_1); -- 
    -- CP-element group 797 transition  input  output  no-bypass 
    -- predecessors 796 
    -- successors 798 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/merge_req
      -- 
    ca_7372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_load_0_ack_1, ack => cp_elements(797)); -- 
    merge_req_7373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => ptr_deref_1055_gather_scatter_req_0); -- 
    -- CP-element group 798 transition  input  output  no-bypass 
    -- predecessors 797 
    -- successors 799 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1056_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1056_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1056_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1055_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1058_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1058_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1058_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_complete/req
      -- 
    merge_ack_7374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_gather_scatter_ack_0, ack => cp_elements(798)); -- 
    req_7387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(798), ack => type_cast_1059_inst_req_0); -- 
    -- CP-element group 799 transition  input  output  no-bypass 
    -- predecessors 798 
    -- successors 802 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1060_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1060_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1060_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1059_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1062_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1062_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1062_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_resize_0/index_resize_req
      -- 
    ack_7388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1059_inst_ack_0, ack => cp_elements(799)); -- 
    index_resize_req_7406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => array_obj_ref_1063_index_0_resize_req_0); -- 
    -- CP-element group 800 transition  bypass 
    -- predecessors 41 
    -- successors 801 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_trigger_
      -- 
    cp_elements(800) <= cp_elements(41);
    -- CP-element group 801 join  transition  output  no-bypass 
    -- predecessors 800 805 
    -- successors 806 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_complete/final_reg_req
      -- 
    cpelement_group_801 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(800);
      predecessors(1) <= cp_elements(805);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(801)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(801),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(801), ack => addr_of_1064_final_reg_req_0); -- 
    -- CP-element group 802 transition  input  output  no-bypass 
    -- predecessors 799 
    -- successors 803 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_7407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_index_0_resize_ack_0, ack => cp_elements(802)); -- 
    scale_rename_req_7411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(802), ack => array_obj_ref_1063_index_0_rename_req_0); -- 
    -- CP-element group 803 transition  input  output  no-bypass 
    -- predecessors 802 
    -- successors 804 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_add_indices/final_index_req
      -- 
    scale_rename_ack_7412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_index_0_rename_ack_0, ack => cp_elements(803)); -- 
    final_index_req_7416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => array_obj_ref_1063_offset_inst_req_0); -- 
    -- CP-element group 804 transition  input  output  no-bypass 
    -- predecessors 803 
    -- successors 805 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_7417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_offset_inst_ack_0, ack => cp_elements(804)); -- 
    sum_rename_req_7421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => array_obj_ref_1063_root_address_inst_req_0); -- 
    -- CP-element group 805 transition  input  no-bypass 
    -- predecessors 804 
    -- successors 801 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1063_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_7422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_root_address_inst_ack_0, ack => cp_elements(805)); -- 
    -- CP-element group 806 transition  input  output  no-bypass 
    -- predecessors 801 
    -- successors 808 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1065_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1065_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1065_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1064_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1066_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1066_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1066_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_7427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1064_final_reg_ack_0, ack => cp_elements(806)); -- 
    base_resize_req_7447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_1067_base_resize_req_0); -- 
    -- CP-element group 807 join  transition  output  bypass 
    -- predecessors 780 790 810 
    -- successors 811 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/split_req
      -- 
    cpelement_group_807 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(780);
      predecessors(1) <= cp_elements(790);
      predecessors(2) <= cp_elements(810);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(807)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(807),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(807), ack => ptr_deref_1067_gather_scatter_req_0); -- 
    -- CP-element group 808 transition  input  output  no-bypass 
    -- predecessors 806 
    -- successors 809 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_base_resize_ack_0, ack => cp_elements(808)); -- 
    sum_rename_req_7452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => ptr_deref_1067_root_address_inst_req_0); -- 
    -- CP-element group 809 transition  input  output  no-bypass 
    -- predecessors 808 
    -- successors 810 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_root_address_inst_ack_0, ack => cp_elements(809)); -- 
    root_register_req_7457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(809), ack => ptr_deref_1067_addr_0_req_0); -- 
    -- CP-element group 810 transition  input  no-bypass 
    -- predecessors 809 
    -- successors 807 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_word_addrgen/root_register_ack
      -- 
    root_register_ack_7458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_addr_0_ack_0, ack => cp_elements(810)); -- 
    -- CP-element group 811 transition  input  output  no-bypass 
    -- predecessors 807 
    -- successors 812 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/word_access_0/rr
      -- 
    split_ack_7463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_gather_scatter_ack_0, ack => cp_elements(811)); -- 
    rr_7470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(811), ack => ptr_deref_1067_store_0_req_0); -- 
    -- CP-element group 812 fork  transition  input  no-bypass 
    -- predecessors 811 
    -- successors 813 839 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_request/word_access/word_access_0/ra
      -- 
    ra_7471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_store_0_ack_0, ack => cp_elements(812)); -- 
    -- CP-element group 813 transition  output  bypass 
    -- predecessors 812 
    -- successors 814 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/word_access_0/cr
      -- 
    cp_elements(813) <= cp_elements(812);
    cr_7481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(813), ack => ptr_deref_1067_store_0_req_1); -- 
    -- CP-element group 814 transition  input  no-bypass 
    -- predecessors 813 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1069_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1067_complete/word_access/word_access_0/ca
      -- 
    ca_7482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1067_store_0_ack_1, ack => cp_elements(814)); -- 
    -- CP-element group 815 join  transition  output  bypass 
    -- predecessors 505 819 
    -- successors 820 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/word_access_0/rr
      -- 
    cpelement_group_815 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(505);
      predecessors(1) <= cp_elements(819);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(815)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(815),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => ptr_deref_1072_load_0_req_0); -- 
    -- CP-element group 816 transition  output  bypass 
    -- predecessors 41 
    -- successors 817 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1071_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1071_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1071_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_addr_resize/base_resize_req
      -- 
    cp_elements(816) <= cp_elements(41);
    base_resize_req_7499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(816), ack => ptr_deref_1072_base_resize_req_0); -- 
    -- CP-element group 817 transition  input  output  no-bypass 
    -- predecessors 816 
    -- successors 818 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_base_resize_ack_0, ack => cp_elements(817)); -- 
    sum_rename_req_7504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(817), ack => ptr_deref_1072_root_address_inst_req_0); -- 
    -- CP-element group 818 transition  input  output  no-bypass 
    -- predecessors 817 
    -- successors 819 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_root_address_inst_ack_0, ack => cp_elements(818)); -- 
    root_register_req_7509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(818), ack => ptr_deref_1072_addr_0_req_0); -- 
    -- CP-element group 819 transition  input  no-bypass 
    -- predecessors 818 
    -- successors 815 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_word_addrgen/root_register_ack
      -- 
    root_register_ack_7510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_addr_0_ack_0, ack => cp_elements(819)); -- 
    -- CP-element group 820 transition  input  output  no-bypass 
    -- predecessors 815 
    -- successors 821 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/word_access_0/cr
      -- 
    ra_7521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_load_0_ack_0, ack => cp_elements(820)); -- 
    cr_7531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(820), ack => ptr_deref_1072_load_0_req_1); -- 
    -- CP-element group 821 transition  input  output  no-bypass 
    -- predecessors 820 
    -- successors 822 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/merge_req
      -- 
    ca_7532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_load_0_ack_1, ack => cp_elements(821)); -- 
    merge_req_7533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => ptr_deref_1072_gather_scatter_req_0); -- 
    -- CP-element group 822 transition  input  no-bypass 
    -- predecessors 821 
    -- successors 839 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1073_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1073_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1073_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1072_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1090_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1090_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1089_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1089_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1089_completed_
      -- 
    merge_ack_7534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1072_gather_scatter_ack_0, ack => cp_elements(822)); -- 
    -- CP-element group 823 join  transition  output  bypass 
    -- predecessors 135 827 
    -- successors 828 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/word_access_0/rr
      -- 
    cpelement_group_823 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(135);
      predecessors(1) <= cp_elements(827);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(823)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(823),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => ptr_deref_1076_load_0_req_0); -- 
    -- CP-element group 824 transition  output  bypass 
    -- predecessors 41 
    -- successors 825 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1075_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1075_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1075_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_addr_resize/base_resize_req
      -- 
    cp_elements(824) <= cp_elements(41);
    base_resize_req_7551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(824), ack => ptr_deref_1076_base_resize_req_0); -- 
    -- CP-element group 825 transition  input  output  no-bypass 
    -- predecessors 824 
    -- successors 826 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_base_resize_ack_0, ack => cp_elements(825)); -- 
    sum_rename_req_7556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(825), ack => ptr_deref_1076_root_address_inst_req_0); -- 
    -- CP-element group 826 transition  input  output  no-bypass 
    -- predecessors 825 
    -- successors 827 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_root_address_inst_ack_0, ack => cp_elements(826)); -- 
    root_register_req_7561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => ptr_deref_1076_addr_0_req_0); -- 
    -- CP-element group 827 transition  input  no-bypass 
    -- predecessors 826 
    -- successors 823 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_word_addrgen/root_register_ack
      -- 
    root_register_ack_7562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_addr_0_ack_0, ack => cp_elements(827)); -- 
    -- CP-element group 828 transition  input  output  no-bypass 
    -- predecessors 823 
    -- successors 829 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/word_access_0/cr
      -- 
    ra_7573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_load_0_ack_0, ack => cp_elements(828)); -- 
    cr_7583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => ptr_deref_1076_load_0_req_1); -- 
    -- CP-element group 829 transition  input  output  no-bypass 
    -- predecessors 828 
    -- successors 830 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/merge_req
      -- 
    ca_7584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_load_0_ack_1, ack => cp_elements(829)); -- 
    merge_req_7585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(829), ack => ptr_deref_1076_gather_scatter_req_0); -- 
    -- CP-element group 830 transition  input  output  no-bypass 
    -- predecessors 829 
    -- successors 831 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1077_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1077_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1077_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1076_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1079_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1079_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1079_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_complete/req
      -- 
    merge_ack_7586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1076_gather_scatter_ack_0, ack => cp_elements(830)); -- 
    req_7599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(830), ack => type_cast_1080_inst_req_0); -- 
    -- CP-element group 831 transition  input  output  no-bypass 
    -- predecessors 830 
    -- successors 834 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1081_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1081_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1081_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1080_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1083_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1083_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1083_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_resize_0/index_resize_req
      -- 
    ack_7600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1080_inst_ack_0, ack => cp_elements(831)); -- 
    index_resize_req_7618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(831), ack => array_obj_ref_1084_index_0_resize_req_0); -- 
    -- CP-element group 832 transition  bypass 
    -- predecessors 41 
    -- successors 833 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_trigger_
      -- 
    cp_elements(832) <= cp_elements(41);
    -- CP-element group 833 join  transition  output  no-bypass 
    -- predecessors 832 837 
    -- successors 838 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_complete/final_reg_req
      -- 
    cpelement_group_833 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(832);
      predecessors(1) <= cp_elements(837);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(833)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(833),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(833), ack => addr_of_1085_final_reg_req_0); -- 
    -- CP-element group 834 transition  input  output  no-bypass 
    -- predecessors 831 
    -- successors 835 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_7619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1084_index_0_resize_ack_0, ack => cp_elements(834)); -- 
    scale_rename_req_7623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(834), ack => array_obj_ref_1084_index_0_rename_req_0); -- 
    -- CP-element group 835 transition  input  output  no-bypass 
    -- predecessors 834 
    -- successors 836 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_add_indices/final_index_req
      -- 
    scale_rename_ack_7624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1084_index_0_rename_ack_0, ack => cp_elements(835)); -- 
    final_index_req_7628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => array_obj_ref_1084_offset_inst_req_0); -- 
    -- CP-element group 836 transition  input  output  no-bypass 
    -- predecessors 835 
    -- successors 837 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_7629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1084_offset_inst_ack_0, ack => cp_elements(836)); -- 
    sum_rename_req_7633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(836), ack => array_obj_ref_1084_root_address_inst_req_0); -- 
    -- CP-element group 837 transition  input  no-bypass 
    -- predecessors 836 
    -- successors 833 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1084_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_7634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1084_root_address_inst_ack_0, ack => cp_elements(837)); -- 
    -- CP-element group 838 transition  input  output  no-bypass 
    -- predecessors 833 
    -- successors 840 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1086_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1086_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1086_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1085_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1087_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1087_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1087_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_7639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1085_final_reg_ack_0, ack => cp_elements(838)); -- 
    base_resize_req_7659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => ptr_deref_1088_base_resize_req_0); -- 
    -- CP-element group 839 join  transition  output  bypass 
    -- predecessors 812 822 842 
    -- successors 843 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/split_req
      -- 
    cpelement_group_839 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(812);
      predecessors(1) <= cp_elements(822);
      predecessors(2) <= cp_elements(842);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(839)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(839),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(839), ack => ptr_deref_1088_gather_scatter_req_0); -- 
    -- CP-element group 840 transition  input  output  no-bypass 
    -- predecessors 838 
    -- successors 841 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_base_resize_ack_0, ack => cp_elements(840)); -- 
    sum_rename_req_7664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => ptr_deref_1088_root_address_inst_req_0); -- 
    -- CP-element group 841 transition  input  output  no-bypass 
    -- predecessors 840 
    -- successors 842 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_root_address_inst_ack_0, ack => cp_elements(841)); -- 
    root_register_req_7669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(841), ack => ptr_deref_1088_addr_0_req_0); -- 
    -- CP-element group 842 transition  input  no-bypass 
    -- predecessors 841 
    -- successors 839 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_word_addrgen/root_register_ack
      -- 
    root_register_ack_7670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_addr_0_ack_0, ack => cp_elements(842)); -- 
    -- CP-element group 843 transition  input  output  no-bypass 
    -- predecessors 839 
    -- successors 844 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/word_access_0/rr
      -- 
    split_ack_7675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_gather_scatter_ack_0, ack => cp_elements(843)); -- 
    rr_7682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => ptr_deref_1088_store_0_req_0); -- 
    -- CP-element group 844 fork  transition  input  no-bypass 
    -- predecessors 843 
    -- successors 845 871 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_request/word_access/word_access_0/ra
      -- 
    ra_7683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_store_0_ack_0, ack => cp_elements(844)); -- 
    -- CP-element group 845 transition  output  bypass 
    -- predecessors 844 
    -- successors 846 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/word_access_0/cr
      -- 
    cp_elements(845) <= cp_elements(844);
    cr_7693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => ptr_deref_1088_store_0_req_1); -- 
    -- CP-element group 846 transition  input  no-bypass 
    -- predecessors 845 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1090_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1088_complete/word_access/word_access_0/ca
      -- 
    ca_7694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1088_store_0_ack_1, ack => cp_elements(846)); -- 
    -- CP-element group 847 join  transition  output  bypass 
    -- predecessors 565 851 
    -- successors 852 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/word_access_0/rr
      -- 
    cpelement_group_847 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(565);
      predecessors(1) <= cp_elements(851);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(847)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(847),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(847), ack => ptr_deref_1093_load_0_req_0); -- 
    -- CP-element group 848 transition  output  bypass 
    -- predecessors 41 
    -- successors 849 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1092_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1092_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1092_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_addr_resize/base_resize_req
      -- 
    cp_elements(848) <= cp_elements(41);
    base_resize_req_7711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => ptr_deref_1093_base_resize_req_0); -- 
    -- CP-element group 849 transition  input  output  no-bypass 
    -- predecessors 848 
    -- successors 850 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7712_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_base_resize_ack_0, ack => cp_elements(849)); -- 
    sum_rename_req_7716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(849), ack => ptr_deref_1093_root_address_inst_req_0); -- 
    -- CP-element group 850 transition  input  output  no-bypass 
    -- predecessors 849 
    -- successors 851 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_root_address_inst_ack_0, ack => cp_elements(850)); -- 
    root_register_req_7721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(850), ack => ptr_deref_1093_addr_0_req_0); -- 
    -- CP-element group 851 transition  input  no-bypass 
    -- predecessors 850 
    -- successors 847 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_word_addrgen/root_register_ack
      -- 
    root_register_ack_7722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_addr_0_ack_0, ack => cp_elements(851)); -- 
    -- CP-element group 852 transition  input  output  no-bypass 
    -- predecessors 847 
    -- successors 853 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/word_access_0/cr
      -- 
    ra_7733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_load_0_ack_0, ack => cp_elements(852)); -- 
    cr_7743_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(852), ack => ptr_deref_1093_load_0_req_1); -- 
    -- CP-element group 853 transition  input  output  no-bypass 
    -- predecessors 852 
    -- successors 854 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/merge_req
      -- 
    ca_7744_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_load_0_ack_1, ack => cp_elements(853)); -- 
    merge_req_7745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => ptr_deref_1093_gather_scatter_req_0); -- 
    -- CP-element group 854 transition  input  no-bypass 
    -- predecessors 853 
    -- successors 871 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1094_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1094_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1094_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1093_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1111_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1111_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1110_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1110_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1110_completed_
      -- 
    merge_ack_7746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1093_gather_scatter_ack_0, ack => cp_elements(854)); -- 
    -- CP-element group 855 join  transition  output  bypass 
    -- predecessors 159 859 
    -- successors 860 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/word_access_0/rr
      -- 
    cpelement_group_855 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(159);
      predecessors(1) <= cp_elements(859);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(855)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(855),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(855), ack => ptr_deref_1097_load_0_req_0); -- 
    -- CP-element group 856 transition  output  bypass 
    -- predecessors 41 
    -- successors 857 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1096_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1096_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1096_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_addr_resize/base_resize_req
      -- 
    cp_elements(856) <= cp_elements(41);
    base_resize_req_7763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(856), ack => ptr_deref_1097_base_resize_req_0); -- 
    -- CP-element group 857 transition  input  output  no-bypass 
    -- predecessors 856 
    -- successors 858 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_base_resize_ack_0, ack => cp_elements(857)); -- 
    sum_rename_req_7768_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => ptr_deref_1097_root_address_inst_req_0); -- 
    -- CP-element group 858 transition  input  output  no-bypass 
    -- predecessors 857 
    -- successors 859 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7769_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_root_address_inst_ack_0, ack => cp_elements(858)); -- 
    root_register_req_7773_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(858), ack => ptr_deref_1097_addr_0_req_0); -- 
    -- CP-element group 859 transition  input  no-bypass 
    -- predecessors 858 
    -- successors 855 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_word_addrgen/root_register_ack
      -- 
    root_register_ack_7774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_addr_0_ack_0, ack => cp_elements(859)); -- 
    -- CP-element group 860 transition  input  output  no-bypass 
    -- predecessors 855 
    -- successors 861 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/word_access_0/cr
      -- 
    ra_7785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_load_0_ack_0, ack => cp_elements(860)); -- 
    cr_7795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(860), ack => ptr_deref_1097_load_0_req_1); -- 
    -- CP-element group 861 transition  input  output  no-bypass 
    -- predecessors 860 
    -- successors 862 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/merge_req
      -- 
    ca_7796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_load_0_ack_1, ack => cp_elements(861)); -- 
    merge_req_7797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(861), ack => ptr_deref_1097_gather_scatter_req_0); -- 
    -- CP-element group 862 transition  input  output  no-bypass 
    -- predecessors 861 
    -- successors 863 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1098_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1098_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1098_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1097_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1100_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1100_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1100_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_complete/req
      -- 
    merge_ack_7798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1097_gather_scatter_ack_0, ack => cp_elements(862)); -- 
    req_7811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(862), ack => type_cast_1101_inst_req_0); -- 
    -- CP-element group 863 transition  input  output  no-bypass 
    -- predecessors 862 
    -- successors 866 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1102_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1102_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1102_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1101_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1104_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1104_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1104_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_resize_0/index_resize_req
      -- 
    ack_7812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1101_inst_ack_0, ack => cp_elements(863)); -- 
    index_resize_req_7830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(863), ack => array_obj_ref_1105_index_0_resize_req_0); -- 
    -- CP-element group 864 transition  bypass 
    -- predecessors 41 
    -- successors 865 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_trigger_
      -- 
    cp_elements(864) <= cp_elements(41);
    -- CP-element group 865 join  transition  output  no-bypass 
    -- predecessors 864 869 
    -- successors 870 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_complete/final_reg_req
      -- 
    cpelement_group_865 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(864);
      predecessors(1) <= cp_elements(869);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(865)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(865),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(865), ack => addr_of_1106_final_reg_req_0); -- 
    -- CP-element group 866 transition  input  output  no-bypass 
    -- predecessors 863 
    -- successors 867 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_7831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_index_0_resize_ack_0, ack => cp_elements(866)); -- 
    scale_rename_req_7835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(866), ack => array_obj_ref_1105_index_0_rename_req_0); -- 
    -- CP-element group 867 transition  input  output  no-bypass 
    -- predecessors 866 
    -- successors 868 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_add_indices/final_index_req
      -- 
    scale_rename_ack_7836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_index_0_rename_ack_0, ack => cp_elements(867)); -- 
    final_index_req_7840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(867), ack => array_obj_ref_1105_offset_inst_req_0); -- 
    -- CP-element group 868 transition  input  output  no-bypass 
    -- predecessors 867 
    -- successors 869 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_7841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_offset_inst_ack_0, ack => cp_elements(868)); -- 
    sum_rename_req_7845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => array_obj_ref_1105_root_address_inst_req_0); -- 
    -- CP-element group 869 transition  input  no-bypass 
    -- predecessors 868 
    -- successors 865 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1105_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_7846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1105_root_address_inst_ack_0, ack => cp_elements(869)); -- 
    -- CP-element group 870 transition  input  output  no-bypass 
    -- predecessors 865 
    -- successors 872 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1107_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1107_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1107_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1106_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1108_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1108_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1108_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_7851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1106_final_reg_ack_0, ack => cp_elements(870)); -- 
    base_resize_req_7871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(870), ack => ptr_deref_1109_base_resize_req_0); -- 
    -- CP-element group 871 join  transition  output  bypass 
    -- predecessors 844 854 874 
    -- successors 875 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/split_req
      -- 
    cpelement_group_871 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(844);
      predecessors(1) <= cp_elements(854);
      predecessors(2) <= cp_elements(874);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(871)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(871),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_7886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => ptr_deref_1109_gather_scatter_req_0); -- 
    -- CP-element group 872 transition  input  output  no-bypass 
    -- predecessors 870 
    -- successors 873 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_base_resize_ack_0, ack => cp_elements(872)); -- 
    sum_rename_req_7876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(872), ack => ptr_deref_1109_root_address_inst_req_0); -- 
    -- CP-element group 873 transition  input  output  no-bypass 
    -- predecessors 872 
    -- successors 874 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_root_address_inst_ack_0, ack => cp_elements(873)); -- 
    root_register_req_7881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(873), ack => ptr_deref_1109_addr_0_req_0); -- 
    -- CP-element group 874 transition  input  no-bypass 
    -- predecessors 873 
    -- successors 871 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_word_addrgen/root_register_ack
      -- 
    root_register_ack_7882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_addr_0_ack_0, ack => cp_elements(874)); -- 
    -- CP-element group 875 transition  input  output  no-bypass 
    -- predecessors 871 
    -- successors 876 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/word_access_0/rr
      -- 
    split_ack_7887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_gather_scatter_ack_0, ack => cp_elements(875)); -- 
    rr_7894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(875), ack => ptr_deref_1109_store_0_req_0); -- 
    -- CP-element group 876 fork  transition  input  no-bypass 
    -- predecessors 875 
    -- successors 877 903 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_request/word_access/word_access_0/ra
      -- 
    ra_7895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_store_0_ack_0, ack => cp_elements(876)); -- 
    -- CP-element group 877 transition  output  bypass 
    -- predecessors 876 
    -- successors 878 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/word_access_0/cr
      -- 
    cp_elements(877) <= cp_elements(876);
    cr_7905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(877), ack => ptr_deref_1109_store_0_req_1); -- 
    -- CP-element group 878 transition  input  no-bypass 
    -- predecessors 877 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1111_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1109_complete/word_access/word_access_0/ca
      -- 
    ca_7906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1109_store_0_ack_1, ack => cp_elements(878)); -- 
    -- CP-element group 879 join  transition  output  bypass 
    -- predecessors 625 883 
    -- successors 884 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/word_access_0/rr
      -- 
    cpelement_group_879 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(625);
      predecessors(1) <= cp_elements(883);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(879)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(879),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7944_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(879), ack => ptr_deref_1114_load_0_req_0); -- 
    -- CP-element group 880 transition  output  bypass 
    -- predecessors 41 
    -- successors 881 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1113_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1113_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1113_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_addr_resize/base_resize_req
      -- 
    cp_elements(880) <= cp_elements(41);
    base_resize_req_7923_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(880), ack => ptr_deref_1114_base_resize_req_0); -- 
    -- CP-element group 881 transition  input  output  no-bypass 
    -- predecessors 880 
    -- successors 882 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7924_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_base_resize_ack_0, ack => cp_elements(881)); -- 
    sum_rename_req_7928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(881), ack => ptr_deref_1114_root_address_inst_req_0); -- 
    -- CP-element group 882 transition  input  output  no-bypass 
    -- predecessors 881 
    -- successors 883 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_root_address_inst_ack_0, ack => cp_elements(882)); -- 
    root_register_req_7933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(882), ack => ptr_deref_1114_addr_0_req_0); -- 
    -- CP-element group 883 transition  input  no-bypass 
    -- predecessors 882 
    -- successors 879 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_word_addrgen/root_register_ack
      -- 
    root_register_ack_7934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_addr_0_ack_0, ack => cp_elements(883)); -- 
    -- CP-element group 884 transition  input  output  no-bypass 
    -- predecessors 879 
    -- successors 885 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/word_access_0/cr
      -- 
    ra_7945_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_load_0_ack_0, ack => cp_elements(884)); -- 
    cr_7955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(884), ack => ptr_deref_1114_load_0_req_1); -- 
    -- CP-element group 885 transition  input  output  no-bypass 
    -- predecessors 884 
    -- successors 886 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/merge_req
      -- 
    ca_7956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_load_0_ack_1, ack => cp_elements(885)); -- 
    merge_req_7957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(885), ack => ptr_deref_1114_gather_scatter_req_0); -- 
    -- CP-element group 886 transition  input  no-bypass 
    -- predecessors 885 
    -- successors 903 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1115_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1115_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1115_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1114_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1132_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1132_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1131_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1131_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1131_completed_
      -- 
    merge_ack_7958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1114_gather_scatter_ack_0, ack => cp_elements(886)); -- 
    -- CP-element group 887 join  transition  output  bypass 
    -- predecessors 183 891 
    -- successors 892 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/word_access_0/rr
      -- 
    cpelement_group_887 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(183);
      predecessors(1) <= cp_elements(891);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(887)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(887),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(887), ack => ptr_deref_1118_load_0_req_0); -- 
    -- CP-element group 888 transition  output  bypass 
    -- predecessors 41 
    -- successors 889 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1117_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1117_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1117_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_addr_resize/base_resize_req
      -- 
    cp_elements(888) <= cp_elements(41);
    base_resize_req_7975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(888), ack => ptr_deref_1118_base_resize_req_0); -- 
    -- CP-element group 889 transition  input  output  no-bypass 
    -- predecessors 888 
    -- successors 890 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_7976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_base_resize_ack_0, ack => cp_elements(889)); -- 
    sum_rename_req_7980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(889), ack => ptr_deref_1118_root_address_inst_req_0); -- 
    -- CP-element group 890 transition  input  output  no-bypass 
    -- predecessors 889 
    -- successors 891 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_word_addrgen/root_register_req
      -- 
    sum_rename_ack_7981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_root_address_inst_ack_0, ack => cp_elements(890)); -- 
    root_register_req_7985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(890), ack => ptr_deref_1118_addr_0_req_0); -- 
    -- CP-element group 891 transition  input  no-bypass 
    -- predecessors 890 
    -- successors 887 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_word_addrgen/root_register_ack
      -- 
    root_register_ack_7986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_addr_0_ack_0, ack => cp_elements(891)); -- 
    -- CP-element group 892 transition  input  output  no-bypass 
    -- predecessors 887 
    -- successors 893 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/word_access_0/cr
      -- 
    ra_7997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_load_0_ack_0, ack => cp_elements(892)); -- 
    cr_8007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(892), ack => ptr_deref_1118_load_0_req_1); -- 
    -- CP-element group 893 transition  input  output  no-bypass 
    -- predecessors 892 
    -- successors 894 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/merge_req
      -- 
    ca_8008_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_load_0_ack_1, ack => cp_elements(893)); -- 
    merge_req_8009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(893), ack => ptr_deref_1118_gather_scatter_req_0); -- 
    -- CP-element group 894 transition  input  output  no-bypass 
    -- predecessors 893 
    -- successors 895 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1119_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1119_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1119_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1118_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1121_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1121_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1121_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_complete/req
      -- 
    merge_ack_8010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1118_gather_scatter_ack_0, ack => cp_elements(894)); -- 
    req_8023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(894), ack => type_cast_1122_inst_req_0); -- 
    -- CP-element group 895 transition  input  output  no-bypass 
    -- predecessors 894 
    -- successors 898 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1123_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1123_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1123_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1122_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1125_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1125_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1125_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_resize_0/index_resize_req
      -- 
    ack_8024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1122_inst_ack_0, ack => cp_elements(895)); -- 
    index_resize_req_8042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(895), ack => array_obj_ref_1126_index_0_resize_req_0); -- 
    -- CP-element group 896 transition  bypass 
    -- predecessors 41 
    -- successors 897 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_trigger_
      -- 
    cp_elements(896) <= cp_elements(41);
    -- CP-element group 897 join  transition  output  no-bypass 
    -- predecessors 896 901 
    -- successors 902 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_complete/final_reg_req
      -- 
    cpelement_group_897 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(896);
      predecessors(1) <= cp_elements(901);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(897)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(897),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8062_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(897), ack => addr_of_1127_final_reg_req_0); -- 
    -- CP-element group 898 transition  input  output  no-bypass 
    -- predecessors 895 
    -- successors 899 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_8043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1126_index_0_resize_ack_0, ack => cp_elements(898)); -- 
    scale_rename_req_8047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(898), ack => array_obj_ref_1126_index_0_rename_req_0); -- 
    -- CP-element group 899 transition  input  output  no-bypass 
    -- predecessors 898 
    -- successors 900 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_add_indices/final_index_req
      -- 
    scale_rename_ack_8048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1126_index_0_rename_ack_0, ack => cp_elements(899)); -- 
    final_index_req_8052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(899), ack => array_obj_ref_1126_offset_inst_req_0); -- 
    -- CP-element group 900 transition  input  output  no-bypass 
    -- predecessors 899 
    -- successors 901 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_8053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1126_offset_inst_ack_0, ack => cp_elements(900)); -- 
    sum_rename_req_8057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(900), ack => array_obj_ref_1126_root_address_inst_req_0); -- 
    -- CP-element group 901 transition  input  no-bypass 
    -- predecessors 900 
    -- successors 897 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1126_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_8058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1126_root_address_inst_ack_0, ack => cp_elements(901)); -- 
    -- CP-element group 902 transition  input  output  no-bypass 
    -- predecessors 897 
    -- successors 904 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1128_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1128_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1128_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1127_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1129_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1129_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1129_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_8063_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1127_final_reg_ack_0, ack => cp_elements(902)); -- 
    base_resize_req_8083_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(902), ack => ptr_deref_1130_base_resize_req_0); -- 
    -- CP-element group 903 join  transition  output  bypass 
    -- predecessors 876 886 906 
    -- successors 907 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/split_req
      -- 
    cpelement_group_903 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(876);
      predecessors(1) <= cp_elements(886);
      predecessors(2) <= cp_elements(906);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(903)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(903),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(903), ack => ptr_deref_1130_gather_scatter_req_0); -- 
    -- CP-element group 904 transition  input  output  no-bypass 
    -- predecessors 902 
    -- successors 905 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8084_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_base_resize_ack_0, ack => cp_elements(904)); -- 
    sum_rename_req_8088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(904), ack => ptr_deref_1130_root_address_inst_req_0); -- 
    -- CP-element group 905 transition  input  output  no-bypass 
    -- predecessors 904 
    -- successors 906 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_root_address_inst_ack_0, ack => cp_elements(905)); -- 
    root_register_req_8093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(905), ack => ptr_deref_1130_addr_0_req_0); -- 
    -- CP-element group 906 transition  input  no-bypass 
    -- predecessors 905 
    -- successors 903 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_word_addrgen/root_register_ack
      -- 
    root_register_ack_8094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_addr_0_ack_0, ack => cp_elements(906)); -- 
    -- CP-element group 907 transition  input  output  no-bypass 
    -- predecessors 903 
    -- successors 908 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/word_access_0/rr
      -- 
    split_ack_8099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_gather_scatter_ack_0, ack => cp_elements(907)); -- 
    rr_8106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(907), ack => ptr_deref_1130_store_0_req_0); -- 
    -- CP-element group 908 fork  transition  input  no-bypass 
    -- predecessors 907 
    -- successors 909 935 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_request/word_access/word_access_0/ra
      -- 
    ra_8107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_store_0_ack_0, ack => cp_elements(908)); -- 
    -- CP-element group 909 transition  output  bypass 
    -- predecessors 908 
    -- successors 910 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/word_access_0/cr
      -- 
    cp_elements(909) <= cp_elements(908);
    cr_8117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => ptr_deref_1130_store_0_req_1); -- 
    -- CP-element group 910 transition  input  no-bypass 
    -- predecessors 909 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1132_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1130_complete/word_access/word_access_0/ca
      -- 
    ca_8118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1130_store_0_ack_1, ack => cp_elements(910)); -- 
    -- CP-element group 911 join  transition  output  bypass 
    -- predecessors 685 915 
    -- successors 916 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/word_access_0/rr
      -- 
    cpelement_group_911 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(685);
      predecessors(1) <= cp_elements(915);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(911)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(911),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => ptr_deref_1135_load_0_req_0); -- 
    -- CP-element group 912 transition  output  bypass 
    -- predecessors 41 
    -- successors 913 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1134_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1134_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1134_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_addr_resize/base_resize_req
      -- 
    cp_elements(912) <= cp_elements(41);
    base_resize_req_8135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(912), ack => ptr_deref_1135_base_resize_req_0); -- 
    -- CP-element group 913 transition  input  output  no-bypass 
    -- predecessors 912 
    -- successors 914 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_base_resize_ack_0, ack => cp_elements(913)); -- 
    sum_rename_req_8140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(913), ack => ptr_deref_1135_root_address_inst_req_0); -- 
    -- CP-element group 914 transition  input  output  no-bypass 
    -- predecessors 913 
    -- successors 915 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8141_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_root_address_inst_ack_0, ack => cp_elements(914)); -- 
    root_register_req_8145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(914), ack => ptr_deref_1135_addr_0_req_0); -- 
    -- CP-element group 915 transition  input  no-bypass 
    -- predecessors 914 
    -- successors 911 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_word_addrgen/root_register_ack
      -- 
    root_register_ack_8146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_addr_0_ack_0, ack => cp_elements(915)); -- 
    -- CP-element group 916 transition  input  output  no-bypass 
    -- predecessors 911 
    -- successors 917 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/word_access_0/cr
      -- 
    ra_8157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_load_0_ack_0, ack => cp_elements(916)); -- 
    cr_8167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(916), ack => ptr_deref_1135_load_0_req_1); -- 
    -- CP-element group 917 transition  input  output  no-bypass 
    -- predecessors 916 
    -- successors 918 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/merge_req
      -- 
    ca_8168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_load_0_ack_1, ack => cp_elements(917)); -- 
    merge_req_8169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(917), ack => ptr_deref_1135_gather_scatter_req_0); -- 
    -- CP-element group 918 transition  input  no-bypass 
    -- predecessors 917 
    -- successors 935 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1136_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1136_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1136_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1135_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1153_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1153_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1152_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1152_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1152_completed_
      -- 
    merge_ack_8170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1135_gather_scatter_ack_0, ack => cp_elements(918)); -- 
    -- CP-element group 919 join  transition  output  bypass 
    -- predecessors 207 923 
    -- successors 924 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/word_access_0/rr
      -- 
    cpelement_group_919 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(207);
      predecessors(1) <= cp_elements(923);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(919)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(919),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(919), ack => ptr_deref_1139_load_0_req_0); -- 
    -- CP-element group 920 transition  output  bypass 
    -- predecessors 41 
    -- successors 921 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1138_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1138_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1138_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_addr_resize/base_resize_req
      -- 
    cp_elements(920) <= cp_elements(41);
    base_resize_req_8187_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(920), ack => ptr_deref_1139_base_resize_req_0); -- 
    -- CP-element group 921 transition  input  output  no-bypass 
    -- predecessors 920 
    -- successors 922 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8188_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_base_resize_ack_0, ack => cp_elements(921)); -- 
    sum_rename_req_8192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(921), ack => ptr_deref_1139_root_address_inst_req_0); -- 
    -- CP-element group 922 transition  input  output  no-bypass 
    -- predecessors 921 
    -- successors 923 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_root_address_inst_ack_0, ack => cp_elements(922)); -- 
    root_register_req_8197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(922), ack => ptr_deref_1139_addr_0_req_0); -- 
    -- CP-element group 923 transition  input  no-bypass 
    -- predecessors 922 
    -- successors 919 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_word_addrgen/root_register_ack
      -- 
    root_register_ack_8198_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_addr_0_ack_0, ack => cp_elements(923)); -- 
    -- CP-element group 924 transition  input  output  no-bypass 
    -- predecessors 919 
    -- successors 925 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/word_access_0/cr
      -- 
    ra_8209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_load_0_ack_0, ack => cp_elements(924)); -- 
    cr_8219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(924), ack => ptr_deref_1139_load_0_req_1); -- 
    -- CP-element group 925 transition  input  output  no-bypass 
    -- predecessors 924 
    -- successors 926 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/merge_req
      -- 
    ca_8220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_load_0_ack_1, ack => cp_elements(925)); -- 
    merge_req_8221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(925), ack => ptr_deref_1139_gather_scatter_req_0); -- 
    -- CP-element group 926 transition  input  output  no-bypass 
    -- predecessors 925 
    -- successors 927 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1140_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1140_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1140_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1139_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1142_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1142_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1142_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_complete/req
      -- 
    merge_ack_8222_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1139_gather_scatter_ack_0, ack => cp_elements(926)); -- 
    req_8235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(926), ack => type_cast_1143_inst_req_0); -- 
    -- CP-element group 927 transition  input  output  no-bypass 
    -- predecessors 926 
    -- successors 930 
    -- members (13) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1144_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1144_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1144_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/type_cast_1143_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_computed_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1146_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1146_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1146_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_resize_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_resize_0/index_resize_req
      -- 
    ack_8236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1143_inst_ack_0, ack => cp_elements(927)); -- 
    index_resize_req_8254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(927), ack => array_obj_ref_1147_index_0_resize_req_0); -- 
    -- CP-element group 928 transition  bypass 
    -- predecessors 41 
    -- successors 929 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_trigger_
      -- 
    cp_elements(928) <= cp_elements(41);
    -- CP-element group 929 join  transition  output  no-bypass 
    -- predecessors 928 933 
    -- successors 934 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_complete/final_reg_req
      -- 
    cpelement_group_929 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(928);
      predecessors(1) <= cp_elements(933);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(929)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(929),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => addr_of_1148_final_reg_req_0); -- 
    -- CP-element group 930 transition  input  output  no-bypass 
    -- predecessors 927 
    -- successors 931 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_resized_0
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_resize_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_scale_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_8255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1147_index_0_resize_ack_0, ack => cp_elements(930)); -- 
    scale_rename_req_8259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(930), ack => array_obj_ref_1147_index_0_rename_req_0); -- 
    -- CP-element group 931 transition  input  output  no-bypass 
    -- predecessors 930 
    -- successors 932 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_indices_scaled
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_scale_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_add_indices/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_add_indices/final_index_req
      -- 
    scale_rename_ack_8260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1147_index_0_rename_ack_0, ack => cp_elements(931)); -- 
    final_index_req_8264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(931), ack => array_obj_ref_1147_offset_inst_req_0); -- 
    -- CP-element group 932 transition  input  output  no-bypass 
    -- predecessors 931 
    -- successors 933 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_offset_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_add_indices/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_add_indices/final_index_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_8265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1147_offset_inst_ack_0, ack => cp_elements(932)); -- 
    sum_rename_req_8269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => array_obj_ref_1147_root_address_inst_req_0); -- 
    -- CP-element group 933 transition  input  no-bypass 
    -- predecessors 932 
    -- successors 929 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/array_obj_ref_1147_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_8270_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1147_root_address_inst_ack_0, ack => cp_elements(933)); -- 
    -- CP-element group 934 transition  input  output  no-bypass 
    -- predecessors 929 
    -- successors 936 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1149_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1149_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1149_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/addr_of_1148_complete/final_reg_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1150_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1150_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/simple_obj_ref_1150_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_addr_resize/base_resize_req
      -- 
    final_reg_ack_8275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1148_final_reg_ack_0, ack => cp_elements(934)); -- 
    base_resize_req_8295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(934), ack => ptr_deref_1151_base_resize_req_0); -- 
    -- CP-element group 935 join  transition  output  bypass 
    -- predecessors 908 918 938 
    -- successors 939 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_trigger_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/split_req
      -- 
    cpelement_group_935 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(908);
      predecessors(1) <= cp_elements(918);
      predecessors(2) <= cp_elements(938);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(935)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(935),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => ptr_deref_1151_gather_scatter_req_0); -- 
    -- CP-element group 936 transition  input  output  no-bypass 
    -- predecessors 934 
    -- successors 937 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_base_resize_ack_0, ack => cp_elements(936)); -- 
    sum_rename_req_8300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(936), ack => ptr_deref_1151_root_address_inst_req_0); -- 
    -- CP-element group 937 transition  input  output  no-bypass 
    -- predecessors 936 
    -- successors 938 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_root_address_inst_ack_0, ack => cp_elements(937)); -- 
    root_register_req_8305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(937), ack => ptr_deref_1151_addr_0_req_0); -- 
    -- CP-element group 938 transition  input  no-bypass 
    -- predecessors 937 
    -- successors 935 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_word_addrgen/root_register_ack
      -- 
    root_register_ack_8306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_addr_0_ack_0, ack => cp_elements(938)); -- 
    -- CP-element group 939 transition  input  output  no-bypass 
    -- predecessors 935 
    -- successors 940 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/word_access_0/rr
      -- 
    split_ack_8311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_gather_scatter_ack_0, ack => cp_elements(939)); -- 
    rr_8318_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => ptr_deref_1151_store_0_req_0); -- 
    -- CP-element group 940 transition  input  output  no-bypass 
    -- predecessors 939 
    -- successors 941 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_active_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/word_access_0/cr
      -- 
    ra_8319_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_store_0_ack_0, ack => cp_elements(940)); -- 
    cr_8329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(940), ack => ptr_deref_1151_store_0_req_1); -- 
    -- CP-element group 941 transition  input  no-bypass 
    -- predecessors 940 
    -- successors 942 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/assign_stmt_1153_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_completed_
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/ptr_deref_1151_complete/word_access/word_access_0/ca
      -- 
    ca_8330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1151_store_0_ack_1, ack => cp_elements(941)); -- 
    -- CP-element group 942 join  transition  no-bypass 
    -- predecessors 50 65 74 89 98 113 122 137 146 161 170 185 194 209 253 267 313 327 373 387 433 447 493 507 553 567 613 627 673 687 718 750 782 814 846 878 910 941 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_491_to_assign_stmt_1153/$exit
      -- 
    cpelement_group_942 : Block -- 
      signal predecessors: BooleanArray(37 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(50);
      predecessors(1) <= cp_elements(65);
      predecessors(2) <= cp_elements(74);
      predecessors(3) <= cp_elements(89);
      predecessors(4) <= cp_elements(98);
      predecessors(5) <= cp_elements(113);
      predecessors(6) <= cp_elements(122);
      predecessors(7) <= cp_elements(137);
      predecessors(8) <= cp_elements(146);
      predecessors(9) <= cp_elements(161);
      predecessors(10) <= cp_elements(170);
      predecessors(11) <= cp_elements(185);
      predecessors(12) <= cp_elements(194);
      predecessors(13) <= cp_elements(209);
      predecessors(14) <= cp_elements(253);
      predecessors(15) <= cp_elements(267);
      predecessors(16) <= cp_elements(313);
      predecessors(17) <= cp_elements(327);
      predecessors(18) <= cp_elements(373);
      predecessors(19) <= cp_elements(387);
      predecessors(20) <= cp_elements(433);
      predecessors(21) <= cp_elements(447);
      predecessors(22) <= cp_elements(493);
      predecessors(23) <= cp_elements(507);
      predecessors(24) <= cp_elements(553);
      predecessors(25) <= cp_elements(567);
      predecessors(26) <= cp_elements(613);
      predecessors(27) <= cp_elements(627);
      predecessors(28) <= cp_elements(673);
      predecessors(29) <= cp_elements(687);
      predecessors(30) <= cp_elements(718);
      predecessors(31) <= cp_elements(750);
      predecessors(32) <= cp_elements(782);
      predecessors(33) <= cp_elements(814);
      predecessors(34) <= cp_elements(846);
      predecessors(35) <= cp_elements(878);
      predecessors(36) <= cp_elements(910);
      predecessors(37) <= cp_elements(941);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(942)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(942),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 943 fork  transition  bypass 
    -- predecessors 3 
    -- successors 944 952 960 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/$entry
      -- 
    cp_elements(943) <= cp_elements(3);
    -- CP-element group 944 transition  output  bypass 
    -- predecessors 943 
    -- successors 945 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1157_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1157_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1157_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_addr_resize/base_resize_req
      -- 
    cp_elements(944) <= cp_elements(943);
    base_resize_req_8350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => ptr_deref_1158_base_resize_req_0); -- 
    -- CP-element group 945 transition  input  output  no-bypass 
    -- predecessors 944 
    -- successors 946 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_addr_resize/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_8351_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_base_resize_ack_0, ack => cp_elements(945)); -- 
    sum_rename_req_8355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(945), ack => ptr_deref_1158_root_address_inst_req_0); -- 
    -- CP-element group 946 transition  input  output  no-bypass 
    -- predecessors 945 
    -- successors 947 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_word_addrgen/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_word_addrgen/root_register_req
      -- 
    sum_rename_ack_8356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_root_address_inst_ack_0, ack => cp_elements(946)); -- 
    root_register_req_8360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(946), ack => ptr_deref_1158_addr_0_req_0); -- 
    -- CP-element group 947 transition  input  output  no-bypass 
    -- predecessors 946 
    -- successors 948 
    -- members (8) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_word_addrgen/root_register_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/word_access_0/rr
      -- 
    root_register_ack_8361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_addr_0_ack_0, ack => cp_elements(947)); -- 
    rr_8371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(947), ack => ptr_deref_1158_load_0_req_0); -- 
    -- CP-element group 948 transition  input  output  no-bypass 
    -- predecessors 947 
    -- successors 949 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/word_access_0/cr
      -- 
    ra_8372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_load_0_ack_0, ack => cp_elements(948)); -- 
    cr_8382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(948), ack => ptr_deref_1158_load_0_req_1); -- 
    -- CP-element group 949 transition  input  output  no-bypass 
    -- predecessors 948 
    -- successors 950 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/merge_req
      -- 
    ca_8383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_load_0_ack_1, ack => cp_elements(949)); -- 
    merge_req_8384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => ptr_deref_1158_gather_scatter_req_0); -- 
    -- CP-element group 950 transition  input  output  no-bypass 
    -- predecessors 949 
    -- successors 951 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1159_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1159_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1159_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1158_complete/merge_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1161_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1161_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1161_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_complete/req
      -- 
    merge_ack_8385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1158_gather_scatter_ack_0, ack => cp_elements(950)); -- 
    req_8398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(950), ack => type_cast_1162_inst_req_0); -- 
    -- CP-element group 951 fork  transition  input  no-bypass 
    -- predecessors 950 
    -- successors 954 955 
    -- members (11) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1163_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1163_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1163_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1162_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1165_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1165_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1165_completed_
      -- 
    ack_8399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1162_inst_ack_0, ack => cp_elements(951)); -- 
    -- CP-element group 952 transition  bypass 
    -- predecessors 943 
    -- successors 967 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_active_
      -- 
    cp_elements(952) <= cp_elements(943);
    -- CP-element group 953 join  transition  output  bypass 
    -- predecessors 956 957 
    -- successors 958 
    -- members (10) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1169_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1169_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1169_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1171_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1171_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1171_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_complete/req
      -- 
    cpelement_group_953 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(956);
      predecessors(1) <= cp_elements(957);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(953)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(953),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(953), ack => type_cast_1172_inst_req_0); -- 
    -- CP-element group 954 transition  output  bypass 
    -- predecessors 951 
    -- successors 956 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_sample_start_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Sample/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Sample/rr
      -- 
    cp_elements(954) <= cp_elements(951);
    rr_8416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(954), ack => binary_1168_inst_req_0); -- 
    -- CP-element group 955 transition  output  bypass 
    -- predecessors 951 
    -- successors 957 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_update_start_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Update/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Update/cr
      -- 
    cp_elements(955) <= cp_elements(951);
    cr_8421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => binary_1168_inst_req_1); -- 
    -- CP-element group 956 transition  input  no-bypass 
    -- predecessors 954 
    -- successors 953 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_sample_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Sample/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Sample/ra
      -- 
    ra_8417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1168_inst_ack_0, ack => cp_elements(956)); -- 
    -- CP-element group 957 transition  input  no-bypass 
    -- predecessors 955 
    -- successors 953 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_update_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Update/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/binary_1168_Update/ca
      -- 
    ca_8422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1168_inst_ack_1, ack => cp_elements(957)); -- 
    -- CP-element group 958 transition  input  no-bypass 
    -- predecessors 953 
    -- successors 959 
    -- members (12) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1173_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1173_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1173_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/type_cast_1172_complete/ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1177_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1177_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1176_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1176_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1176_completed_
      -- 
    ack_8436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1172_inst_ack_0, ack => cp_elements(958)); -- 
    -- CP-element group 959 join  transition  output  bypass 
    -- predecessors 958 963 
    -- successors 964 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/split_req
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_trigger_
      -- 
    cpelement_group_959 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(958);
      predecessors(1) <= cp_elements(963);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(959)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(959),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(959), ack => ptr_deref_1175_gather_scatter_req_0); -- 
    -- CP-element group 960 transition  output  bypass 
    -- predecessors 943 
    -- successors 961 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1174_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_addr_resize/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1174_trigger_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/simple_obj_ref_1174_active_
      -- 
    cp_elements(960) <= cp_elements(943);
    base_resize_req_8456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(960), ack => ptr_deref_1175_base_resize_req_0); -- 
    -- CP-element group 961 transition  input  output  no-bypass 
    -- predecessors 960 
    -- successors 962 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_plus_offset/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_address_resized
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_addr_resize/$exit
      -- 
    base_resize_ack_8457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_base_resize_ack_0, ack => cp_elements(961)); -- 
    sum_rename_req_8461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => ptr_deref_1175_root_address_inst_req_0); -- 
    -- CP-element group 962 transition  input  output  no-bypass 
    -- predecessors 961 
    -- successors 963 
    -- members (5) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_root_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_word_addrgen/root_register_req
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_plus_offset/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_word_addrgen/$entry
      -- 
    sum_rename_ack_8462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_root_address_inst_ack_0, ack => cp_elements(962)); -- 
    root_register_req_8466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => ptr_deref_1175_addr_0_req_0); -- 
    -- CP-element group 963 transition  input  no-bypass 
    -- predecessors 962 
    -- successors 959 
    -- members (3) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_word_address_calculated
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_word_addrgen/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_word_addrgen/root_register_ack
      -- 
    root_register_ack_8467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_addr_0_ack_0, ack => cp_elements(963)); -- 
    -- CP-element group 964 transition  input  output  no-bypass 
    -- predecessors 959 
    -- successors 965 
    -- members (4) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/split_ack
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/word_access_0/rr
      -- 
    split_ack_8472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_gather_scatter_ack_0, ack => cp_elements(964)); -- 
    rr_8479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(964), ack => ptr_deref_1175_store_0_req_0); -- 
    -- CP-element group 965 transition  input  output  no-bypass 
    -- predecessors 964 
    -- successors 966 
    -- members (9) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_active_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/word_access_0/cr
      -- 
    ra_8480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_store_0_ack_0, ack => cp_elements(965)); -- 
    cr_8490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(965), ack => ptr_deref_1175_store_0_req_1); -- 
    -- CP-element group 966 transition  input  no-bypass 
    -- predecessors 965 
    -- successors 967 
    -- members (6) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/assign_stmt_1177_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_completed_
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/ptr_deref_1175_complete/word_access/word_access_0/ca
      -- 
    ca_8491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1175_store_0_ack_1, ack => cp_elements(966)); -- 
    -- CP-element group 967 join  transition  no-bypass 
    -- predecessors 952 966 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_377/assign_stmt_1159_to_assign_stmt_1177/$exit
      -- 
    cpelement_group_967 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(952);
      predecessors(1) <= cp_elements(966);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => false,
        name => " cp_elements(967)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(967),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 968 merge  place  bypass 
    -- predecessors 4 14 
    -- successors 969 
    -- members (1) 
      -- 	branch_block_stmt_377/merge_stmt_464_PhiReqMerge
      -- 
    cp_elements(968) <= OrReduce(cp_elements(4) & cp_elements(14));
    -- CP-element group 969 transition  place  bypass 
    -- predecessors 968 
    -- successors 15 
    -- members (5) 
      -- 	branch_block_stmt_377/merge_stmt_464__exit__
      -- 	branch_block_stmt_377/assign_stmt_468_to_assign_stmt_480__entry__
      -- 	branch_block_stmt_377/merge_stmt_464_PhiAck/$entry
      -- 	branch_block_stmt_377/merge_stmt_464_PhiAck/$exit
      -- 	branch_block_stmt_377/merge_stmt_464_PhiAck/dummy
      -- 
    cp_elements(969) <= cp_elements(968);
    -- CP-element group 970 transition  dead  bypass 
    -- predecessors 34 
    -- successors 971 
    -- members (1) 
      -- 	branch_block_stmt_377/merge_stmt_487_dead_link/dead_transition
      -- 
    cp_elements(970) <= false;
    -- CP-element group 971 transition  bypass 
    -- predecessors 970 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_377/merge_stmt_487_dead_link/$exit
      -- 
    cp_elements(971) <= cp_elements(970);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I1_401 : std_logic_vector(31 downto 0);
    signal I2_405 : std_logic_vector(31 downto 0);
    signal I3_409 : std_logic_vector(31 downto 0);
    signal I4_413 : std_logic_vector(31 downto 0);
    signal I5_417 : std_logic_vector(31 downto 0);
    signal I6_421 : std_logic_vector(31 downto 0);
    signal I7_425 : std_logic_vector(31 downto 0);
    signal I_397 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1000_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1000_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1000_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1000_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1021_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1021_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1021_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1021_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1042_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1042_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1042_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1042_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1063_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1063_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1063_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1063_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1084_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1084_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1084_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1084_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1105_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1105_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1105_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1105_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1126_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1126_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1126_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1126_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1147_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_1147_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_1147_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_1147_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_652_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_652_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_652_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_652_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_669_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_669_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_669_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_669_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_695_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_695_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_695_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_695_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_712_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_712_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_712_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_712_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_738_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_738_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_738_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_738_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_755_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_755_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_755_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_755_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_781_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_781_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_781_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_781_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_798_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_798_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_798_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_798_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_824_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_824_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_824_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_824_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_841_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_841_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_841_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_841_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_867_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_867_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_867_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_867_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_884_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_884_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_884_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_884_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_910_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_910_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_910_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_910_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_927_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_927_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_927_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_927_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_953_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_953_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_953_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_953_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_970_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_970_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_970_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_970_root_address : std_logic_vector(6 downto 0);
    signal c0_429 : std_logic_vector(31 downto 0);
    signal c1_433 : std_logic_vector(31 downto 0);
    signal c2_437 : std_logic_vector(31 downto 0);
    signal c3_441 : std_logic_vector(31 downto 0);
    signal c4_445 : std_logic_vector(31 downto 0);
    signal c5_449 : std_logic_vector(31 downto 0);
    signal c6_453 : std_logic_vector(31 downto 0);
    signal c7_457 : std_logic_vector(31 downto 0);
    signal iNsTr_100_895 : std_logic_vector(31 downto 0);
    signal iNsTr_102_903 : std_logic_vector(7 downto 0);
    signal iNsTr_103_907 : std_logic_vector(31 downto 0);
    signal iNsTr_104_912 : std_logic_vector(31 downto 0);
    signal iNsTr_105_916 : std_logic_vector(31 downto 0);
    signal iNsTr_106_920 : std_logic_vector(7 downto 0);
    signal iNsTr_107_924 : std_logic_vector(31 downto 0);
    signal iNsTr_108_929 : std_logic_vector(31 downto 0);
    signal iNsTr_109_933 : std_logic_vector(31 downto 0);
    signal iNsTr_10_505 : std_logic_vector(7 downto 0);
    signal iNsTr_110_938 : std_logic_vector(31 downto 0);
    signal iNsTr_112_946 : std_logic_vector(7 downto 0);
    signal iNsTr_113_950 : std_logic_vector(31 downto 0);
    signal iNsTr_114_955 : std_logic_vector(31 downto 0);
    signal iNsTr_115_959 : std_logic_vector(31 downto 0);
    signal iNsTr_116_963 : std_logic_vector(7 downto 0);
    signal iNsTr_117_967 : std_logic_vector(31 downto 0);
    signal iNsTr_118_972 : std_logic_vector(31 downto 0);
    signal iNsTr_119_976 : std_logic_vector(31 downto 0);
    signal iNsTr_120_981 : std_logic_vector(31 downto 0);
    signal iNsTr_122_989 : std_logic_vector(31 downto 0);
    signal iNsTr_123_993 : std_logic_vector(7 downto 0);
    signal iNsTr_124_997 : std_logic_vector(31 downto 0);
    signal iNsTr_125_1002 : std_logic_vector(31 downto 0);
    signal iNsTr_127_1010 : std_logic_vector(31 downto 0);
    signal iNsTr_128_1014 : std_logic_vector(7 downto 0);
    signal iNsTr_129_1018 : std_logic_vector(31 downto 0);
    signal iNsTr_12_513 : std_logic_vector(7 downto 0);
    signal iNsTr_130_1023 : std_logic_vector(31 downto 0);
    signal iNsTr_132_1031 : std_logic_vector(31 downto 0);
    signal iNsTr_133_1035 : std_logic_vector(7 downto 0);
    signal iNsTr_134_1039 : std_logic_vector(31 downto 0);
    signal iNsTr_135_1044 : std_logic_vector(31 downto 0);
    signal iNsTr_137_1052 : std_logic_vector(31 downto 0);
    signal iNsTr_138_1056 : std_logic_vector(7 downto 0);
    signal iNsTr_139_1060 : std_logic_vector(31 downto 0);
    signal iNsTr_13_517 : std_logic_vector(31 downto 0);
    signal iNsTr_140_1065 : std_logic_vector(31 downto 0);
    signal iNsTr_142_1073 : std_logic_vector(31 downto 0);
    signal iNsTr_143_1077 : std_logic_vector(7 downto 0);
    signal iNsTr_144_1081 : std_logic_vector(31 downto 0);
    signal iNsTr_145_1086 : std_logic_vector(31 downto 0);
    signal iNsTr_147_1094 : std_logic_vector(31 downto 0);
    signal iNsTr_148_1098 : std_logic_vector(7 downto 0);
    signal iNsTr_149_1102 : std_logic_vector(31 downto 0);
    signal iNsTr_14_523 : std_logic_vector(31 downto 0);
    signal iNsTr_150_1107 : std_logic_vector(31 downto 0);
    signal iNsTr_152_1115 : std_logic_vector(31 downto 0);
    signal iNsTr_153_1119 : std_logic_vector(7 downto 0);
    signal iNsTr_154_1123 : std_logic_vector(31 downto 0);
    signal iNsTr_155_1128 : std_logic_vector(31 downto 0);
    signal iNsTr_157_1136 : std_logic_vector(31 downto 0);
    signal iNsTr_158_1140 : std_logic_vector(7 downto 0);
    signal iNsTr_159_1144 : std_logic_vector(31 downto 0);
    signal iNsTr_15_527 : std_logic_vector(7 downto 0);
    signal iNsTr_160_1149 : std_logic_vector(31 downto 0);
    signal iNsTr_164_1159 : std_logic_vector(7 downto 0);
    signal iNsTr_165_1163 : std_logic_vector(31 downto 0);
    signal iNsTr_166_1169 : std_logic_vector(31 downto 0);
    signal iNsTr_167_1173 : std_logic_vector(7 downto 0);
    signal iNsTr_17_535 : std_logic_vector(7 downto 0);
    signal iNsTr_18_539 : std_logic_vector(31 downto 0);
    signal iNsTr_19_545 : std_logic_vector(31 downto 0);
    signal iNsTr_20_549 : std_logic_vector(7 downto 0);
    signal iNsTr_22_557 : std_logic_vector(7 downto 0);
    signal iNsTr_23_561 : std_logic_vector(31 downto 0);
    signal iNsTr_24_567 : std_logic_vector(31 downto 0);
    signal iNsTr_25_571 : std_logic_vector(7 downto 0);
    signal iNsTr_27_579 : std_logic_vector(7 downto 0);
    signal iNsTr_28_583 : std_logic_vector(31 downto 0);
    signal iNsTr_29_589 : std_logic_vector(31 downto 0);
    signal iNsTr_2_468 : std_logic_vector(7 downto 0);
    signal iNsTr_30_593 : std_logic_vector(7 downto 0);
    signal iNsTr_32_601 : std_logic_vector(7 downto 0);
    signal iNsTr_33_605 : std_logic_vector(31 downto 0);
    signal iNsTr_34_611 : std_logic_vector(31 downto 0);
    signal iNsTr_35_615 : std_logic_vector(7 downto 0);
    signal iNsTr_37_623 : std_logic_vector(7 downto 0);
    signal iNsTr_38_627 : std_logic_vector(31 downto 0);
    signal iNsTr_39_633 : std_logic_vector(31 downto 0);
    signal iNsTr_3_472 : std_logic_vector(31 downto 0);
    signal iNsTr_40_637 : std_logic_vector(7 downto 0);
    signal iNsTr_42_645 : std_logic_vector(7 downto 0);
    signal iNsTr_43_649 : std_logic_vector(31 downto 0);
    signal iNsTr_44_654 : std_logic_vector(31 downto 0);
    signal iNsTr_45_658 : std_logic_vector(31 downto 0);
    signal iNsTr_46_662 : std_logic_vector(7 downto 0);
    signal iNsTr_47_666 : std_logic_vector(31 downto 0);
    signal iNsTr_48_671 : std_logic_vector(31 downto 0);
    signal iNsTr_49_675 : std_logic_vector(31 downto 0);
    signal iNsTr_4_480 : std_logic_vector(0 downto 0);
    signal iNsTr_50_680 : std_logic_vector(31 downto 0);
    signal iNsTr_52_688 : std_logic_vector(7 downto 0);
    signal iNsTr_53_692 : std_logic_vector(31 downto 0);
    signal iNsTr_54_697 : std_logic_vector(31 downto 0);
    signal iNsTr_55_701 : std_logic_vector(31 downto 0);
    signal iNsTr_56_705 : std_logic_vector(7 downto 0);
    signal iNsTr_57_709 : std_logic_vector(31 downto 0);
    signal iNsTr_58_714 : std_logic_vector(31 downto 0);
    signal iNsTr_59_718 : std_logic_vector(31 downto 0);
    signal iNsTr_60_723 : std_logic_vector(31 downto 0);
    signal iNsTr_62_731 : std_logic_vector(7 downto 0);
    signal iNsTr_63_735 : std_logic_vector(31 downto 0);
    signal iNsTr_64_740 : std_logic_vector(31 downto 0);
    signal iNsTr_65_744 : std_logic_vector(31 downto 0);
    signal iNsTr_66_748 : std_logic_vector(7 downto 0);
    signal iNsTr_67_752 : std_logic_vector(31 downto 0);
    signal iNsTr_68_757 : std_logic_vector(31 downto 0);
    signal iNsTr_69_761 : std_logic_vector(31 downto 0);
    signal iNsTr_70_766 : std_logic_vector(31 downto 0);
    signal iNsTr_72_774 : std_logic_vector(7 downto 0);
    signal iNsTr_73_778 : std_logic_vector(31 downto 0);
    signal iNsTr_74_783 : std_logic_vector(31 downto 0);
    signal iNsTr_75_787 : std_logic_vector(31 downto 0);
    signal iNsTr_76_791 : std_logic_vector(7 downto 0);
    signal iNsTr_77_795 : std_logic_vector(31 downto 0);
    signal iNsTr_78_800 : std_logic_vector(31 downto 0);
    signal iNsTr_79_804 : std_logic_vector(31 downto 0);
    signal iNsTr_7_491 : std_logic_vector(7 downto 0);
    signal iNsTr_80_809 : std_logic_vector(31 downto 0);
    signal iNsTr_82_817 : std_logic_vector(7 downto 0);
    signal iNsTr_83_821 : std_logic_vector(31 downto 0);
    signal iNsTr_84_826 : std_logic_vector(31 downto 0);
    signal iNsTr_85_830 : std_logic_vector(31 downto 0);
    signal iNsTr_86_834 : std_logic_vector(7 downto 0);
    signal iNsTr_87_838 : std_logic_vector(31 downto 0);
    signal iNsTr_88_843 : std_logic_vector(31 downto 0);
    signal iNsTr_89_847 : std_logic_vector(31 downto 0);
    signal iNsTr_8_495 : std_logic_vector(31 downto 0);
    signal iNsTr_90_852 : std_logic_vector(31 downto 0);
    signal iNsTr_92_860 : std_logic_vector(7 downto 0);
    signal iNsTr_93_864 : std_logic_vector(31 downto 0);
    signal iNsTr_94_869 : std_logic_vector(31 downto 0);
    signal iNsTr_95_873 : std_logic_vector(31 downto 0);
    signal iNsTr_96_877 : std_logic_vector(7 downto 0);
    signal iNsTr_97_881 : std_logic_vector(31 downto 0);
    signal iNsTr_98_886 : std_logic_vector(31 downto 0);
    signal iNsTr_99_890 : std_logic_vector(31 downto 0);
    signal iNsTr_9_501 : std_logic_vector(31 downto 0);
    signal ptr_deref_1004_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1004_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1004_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1004_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1004_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1004_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1009_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1009_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1009_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1009_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1009_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1013_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1013_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1013_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1013_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1013_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1025_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1025_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1025_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1025_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1025_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1025_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1030_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1030_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1030_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1030_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1030_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1034_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1034_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1034_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1034_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1034_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1046_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1046_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1046_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1046_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1046_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1046_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1051_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1051_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1051_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1051_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1051_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1055_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1055_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1055_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1055_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1055_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1067_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1067_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1067_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1067_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1067_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1067_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1072_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1072_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1072_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1072_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1072_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1076_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1076_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1076_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1076_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1076_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1088_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1088_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1088_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1088_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1088_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1088_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1093_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1093_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1093_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1093_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1093_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1097_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1097_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1097_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1097_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1097_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1109_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1109_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1109_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1109_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1114_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1114_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1114_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1114_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1114_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1118_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1118_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1118_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1118_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1118_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1130_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1130_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1130_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1130_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1130_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1130_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1135_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1135_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1135_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1135_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1135_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1139_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1139_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1139_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1139_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1139_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1151_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1151_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1151_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_1151_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1151_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1151_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_1158_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1158_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1158_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1158_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1158_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1175_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1175_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1175_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_1175_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1175_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_1175_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_459_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_459_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_459_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_459_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_459_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_459_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_467_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_467_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_467_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_467_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_467_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_490_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_490_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_490_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_490_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_490_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_507_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_507_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_507_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_507_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_507_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_507_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_512_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_512_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_512_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_512_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_512_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_529_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_529_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_529_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_529_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_529_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_529_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_534_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_534_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_534_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_534_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_534_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_551_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_551_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_551_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_551_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_551_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_551_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_556_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_556_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_556_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_556_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_556_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_573_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_573_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_573_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_573_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_573_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_573_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_578_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_578_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_578_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_578_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_578_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_595_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_595_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_595_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_595_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_595_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_595_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_600_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_600_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_600_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_600_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_600_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_617_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_617_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_617_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_617_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_617_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_617_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_622_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_622_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_622_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_622_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_622_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_639_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_639_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_639_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_639_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_639_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_639_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_644_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_644_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_644_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_644_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_644_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_657_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_657_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_657_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_657_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_657_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_661_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_661_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_661_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_661_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_661_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_674_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_674_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_674_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_674_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_674_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_682_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_682_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_682_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_682_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_682_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_682_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_687_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_687_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_687_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_687_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_687_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_700_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_700_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_700_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_700_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_700_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_704_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_704_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_704_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_704_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_704_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_717_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_717_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_717_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_717_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_717_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_725_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_725_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_725_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_725_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_725_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_725_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_730_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_730_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_730_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_730_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_730_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_743_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_743_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_743_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_743_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_743_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_747_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_747_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_747_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_747_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_747_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_760_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_760_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_760_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_760_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_760_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_768_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_768_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_768_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_768_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_768_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_768_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_773_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_773_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_773_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_773_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_773_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_786_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_786_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_786_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_786_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_786_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_790_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_790_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_790_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_790_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_790_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_803_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_803_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_803_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_803_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_803_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_811_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_811_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_811_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_811_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_811_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_811_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_816_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_816_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_816_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_816_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_816_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_829_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_829_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_829_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_829_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_829_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_833_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_833_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_833_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_833_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_833_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_846_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_846_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_846_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_846_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_846_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_854_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_854_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_854_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_854_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_854_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_854_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_859_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_859_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_859_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_859_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_859_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_872_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_872_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_872_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_872_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_872_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_876_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_876_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_876_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_876_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_876_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_889_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_889_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_889_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_889_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_889_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_897_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_897_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_897_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_897_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_897_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_897_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_902_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_902_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_902_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_902_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_902_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_915_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_915_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_915_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_915_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_915_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_919_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_919_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_919_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_919_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_919_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_932_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_932_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_932_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_932_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_932_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_940_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_940_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_940_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_940_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_940_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_940_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_945_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_945_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_945_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_945_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_945_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_958_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_958_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_958_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_958_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_958_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_962_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_962_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_962_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_962_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_962_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_975_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_975_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_975_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_975_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_975_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_983_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_983_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_983_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_983_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_983_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_983_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_988_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_988_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_988_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_988_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_988_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_992_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_992_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_992_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_992_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_992_word_offset_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1020_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1020_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1041_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1041_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1062_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1062_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1083_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1083_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1104_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1104_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1125_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1125_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1146_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_1146_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_651_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_651_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_668_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_668_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_694_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_694_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_711_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_711_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_737_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_737_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_754_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_754_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_780_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_780_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_797_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_797_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_823_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_823_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_840_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_840_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_866_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_866_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_883_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_883_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_909_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_909_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_926_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_926_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_952_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_952_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_969_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_969_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_999_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_999_scaled : std_logic_vector(6 downto 0);
    signal type_cast_1167_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_461_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_475_wire : std_logic_vector(31 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_521_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_543_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_565_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_609_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_631_wire_constant : std_logic_vector(31 downto 0);
    signal xxx_vectorSum_xxbodyxxI1_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI2_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI3_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI4_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI5_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI6_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI7_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxI_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc0_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc1_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc2_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc3_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc4_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc5_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc6_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxx_vectorSum_xxbodyxxc7_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    I1_401 <= "00000000000000000000000000000000";
    I2_405 <= "00000000000000000000000000000000";
    I3_409 <= "00000000000000000000000000000000";
    I4_413 <= "00000000000000000000000000000000";
    I5_417 <= "00000000000000000000000000000000";
    I6_421 <= "00000000000000000000000000000000";
    I7_425 <= "00000000000000000000000000000000";
    I_397 <= "00000000000000000000000000000000";
    array_obj_ref_1000_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1000_resized_base_address <= "0000000";
    array_obj_ref_1021_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1021_resized_base_address <= "0000000";
    array_obj_ref_1042_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1042_resized_base_address <= "0000000";
    array_obj_ref_1063_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1063_resized_base_address <= "0000000";
    array_obj_ref_1084_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1084_resized_base_address <= "0000000";
    array_obj_ref_1105_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1105_resized_base_address <= "0000000";
    array_obj_ref_1126_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1126_resized_base_address <= "0000000";
    array_obj_ref_1147_offset_scale_factor_0 <= "0000001";
    array_obj_ref_1147_resized_base_address <= "0000000";
    array_obj_ref_652_offset_scale_factor_0 <= "0000001";
    array_obj_ref_652_resized_base_address <= "0000000";
    array_obj_ref_669_offset_scale_factor_0 <= "0000001";
    array_obj_ref_669_resized_base_address <= "0000000";
    array_obj_ref_695_offset_scale_factor_0 <= "0000001";
    array_obj_ref_695_resized_base_address <= "0000000";
    array_obj_ref_712_offset_scale_factor_0 <= "0000001";
    array_obj_ref_712_resized_base_address <= "0000000";
    array_obj_ref_738_offset_scale_factor_0 <= "0000001";
    array_obj_ref_738_resized_base_address <= "0000000";
    array_obj_ref_755_offset_scale_factor_0 <= "0000001";
    array_obj_ref_755_resized_base_address <= "0000000";
    array_obj_ref_781_offset_scale_factor_0 <= "0000001";
    array_obj_ref_781_resized_base_address <= "0000000";
    array_obj_ref_798_offset_scale_factor_0 <= "0000001";
    array_obj_ref_798_resized_base_address <= "0000000";
    array_obj_ref_824_offset_scale_factor_0 <= "0000001";
    array_obj_ref_824_resized_base_address <= "0000000";
    array_obj_ref_841_offset_scale_factor_0 <= "0000001";
    array_obj_ref_841_resized_base_address <= "0000000";
    array_obj_ref_867_offset_scale_factor_0 <= "0000001";
    array_obj_ref_867_resized_base_address <= "0000000";
    array_obj_ref_884_offset_scale_factor_0 <= "0000001";
    array_obj_ref_884_resized_base_address <= "0000000";
    array_obj_ref_910_offset_scale_factor_0 <= "0000001";
    array_obj_ref_910_resized_base_address <= "0000000";
    array_obj_ref_927_offset_scale_factor_0 <= "0000001";
    array_obj_ref_927_resized_base_address <= "0000000";
    array_obj_ref_953_offset_scale_factor_0 <= "0000001";
    array_obj_ref_953_resized_base_address <= "0000000";
    array_obj_ref_970_offset_scale_factor_0 <= "0000001";
    array_obj_ref_970_resized_base_address <= "0000000";
    c0_429 <= "00000000000000000000000000000000";
    c1_433 <= "00000000000000000000000000000000";
    c2_437 <= "00000000000000000000000000000000";
    c3_441 <= "00000000000000000000000000000000";
    c4_445 <= "00000000000000000000000000000000";
    c5_449 <= "00000000000000000000000000000000";
    c6_453 <= "00000000000000000000000000000000";
    c7_457 <= "00000000000000000000000000000000";
    ptr_deref_1004_word_offset_0 <= "0000000";
    ptr_deref_1009_word_offset_0 <= "0";
    ptr_deref_1013_word_offset_0 <= "0";
    ptr_deref_1025_word_offset_0 <= "0000000";
    ptr_deref_1030_word_offset_0 <= "0";
    ptr_deref_1034_word_offset_0 <= "0";
    ptr_deref_1046_word_offset_0 <= "0000000";
    ptr_deref_1051_word_offset_0 <= "0";
    ptr_deref_1055_word_offset_0 <= "0";
    ptr_deref_1067_word_offset_0 <= "0000000";
    ptr_deref_1072_word_offset_0 <= "0";
    ptr_deref_1076_word_offset_0 <= "0";
    ptr_deref_1088_word_offset_0 <= "0000000";
    ptr_deref_1093_word_offset_0 <= "0";
    ptr_deref_1097_word_offset_0 <= "0";
    ptr_deref_1109_word_offset_0 <= "0000000";
    ptr_deref_1114_word_offset_0 <= "0";
    ptr_deref_1118_word_offset_0 <= "0";
    ptr_deref_1130_word_offset_0 <= "0000000";
    ptr_deref_1135_word_offset_0 <= "0";
    ptr_deref_1139_word_offset_0 <= "0";
    ptr_deref_1151_word_offset_0 <= "0000000";
    ptr_deref_1158_word_offset_0 <= "0";
    ptr_deref_1175_word_offset_0 <= "0";
    ptr_deref_459_word_offset_0 <= "0";
    ptr_deref_467_word_offset_0 <= "0";
    ptr_deref_490_word_offset_0 <= "0";
    ptr_deref_507_word_offset_0 <= "0";
    ptr_deref_512_word_offset_0 <= "0";
    ptr_deref_529_word_offset_0 <= "0";
    ptr_deref_534_word_offset_0 <= "0";
    ptr_deref_551_word_offset_0 <= "0";
    ptr_deref_556_word_offset_0 <= "0";
    ptr_deref_573_word_offset_0 <= "0";
    ptr_deref_578_word_offset_0 <= "0";
    ptr_deref_595_word_offset_0 <= "0";
    ptr_deref_600_word_offset_0 <= "0";
    ptr_deref_617_word_offset_0 <= "0";
    ptr_deref_622_word_offset_0 <= "0";
    ptr_deref_639_word_offset_0 <= "0";
    ptr_deref_644_word_offset_0 <= "0";
    ptr_deref_657_word_offset_0 <= "0000000";
    ptr_deref_661_word_offset_0 <= "0";
    ptr_deref_674_word_offset_0 <= "0000000";
    ptr_deref_682_word_offset_0 <= "0";
    ptr_deref_687_word_offset_0 <= "0";
    ptr_deref_700_word_offset_0 <= "0000000";
    ptr_deref_704_word_offset_0 <= "0";
    ptr_deref_717_word_offset_0 <= "0000000";
    ptr_deref_725_word_offset_0 <= "0";
    ptr_deref_730_word_offset_0 <= "0";
    ptr_deref_743_word_offset_0 <= "0000000";
    ptr_deref_747_word_offset_0 <= "0";
    ptr_deref_760_word_offset_0 <= "0000000";
    ptr_deref_768_word_offset_0 <= "0";
    ptr_deref_773_word_offset_0 <= "0";
    ptr_deref_786_word_offset_0 <= "0000000";
    ptr_deref_790_word_offset_0 <= "0";
    ptr_deref_803_word_offset_0 <= "0000000";
    ptr_deref_811_word_offset_0 <= "0";
    ptr_deref_816_word_offset_0 <= "0";
    ptr_deref_829_word_offset_0 <= "0000000";
    ptr_deref_833_word_offset_0 <= "0";
    ptr_deref_846_word_offset_0 <= "0000000";
    ptr_deref_854_word_offset_0 <= "0";
    ptr_deref_859_word_offset_0 <= "0";
    ptr_deref_872_word_offset_0 <= "0000000";
    ptr_deref_876_word_offset_0 <= "0";
    ptr_deref_889_word_offset_0 <= "0000000";
    ptr_deref_897_word_offset_0 <= "0";
    ptr_deref_902_word_offset_0 <= "0";
    ptr_deref_915_word_offset_0 <= "0000000";
    ptr_deref_919_word_offset_0 <= "0";
    ptr_deref_932_word_offset_0 <= "0000000";
    ptr_deref_940_word_offset_0 <= "0";
    ptr_deref_945_word_offset_0 <= "0";
    ptr_deref_958_word_offset_0 <= "0000000";
    ptr_deref_962_word_offset_0 <= "0";
    ptr_deref_975_word_offset_0 <= "0000000";
    ptr_deref_983_word_offset_0 <= "0";
    ptr_deref_988_word_offset_0 <= "0";
    ptr_deref_992_word_offset_0 <= "0";
    type_cast_1167_wire_constant <= "00000000000000000000000000001000";
    type_cast_461_wire_constant <= "00000000";
    type_cast_478_wire_constant <= "00000000000000000000000001000000";
    type_cast_499_wire_constant <= "00000000000000000000000000000001";
    type_cast_521_wire_constant <= "00000000000000000000000000000010";
    type_cast_543_wire_constant <= "00000000000000000000000000000011";
    type_cast_565_wire_constant <= "00000000000000000000000000000100";
    type_cast_587_wire_constant <= "00000000000000000000000000000101";
    type_cast_609_wire_constant <= "00000000000000000000000000000110";
    type_cast_631_wire_constant <= "00000000000000000000000000000111";
    xxx_vectorSum_xxbodyxxI1_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI2_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI3_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI4_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI5_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI6_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI7_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxI_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc0_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc1_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc2_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc3_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc4_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc5_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc6_alloc_base_address <= "0";
    xxx_vectorSum_xxbodyxxc7_alloc_base_address <= "0";
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1001_final_reg_req_0,addr_of_1001_final_reg_ack_0,sl_one,"addr_of_1001_final_reg ",false,array_obj_ref_1000_root_address,
    false,iNsTr_125_1002);
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1001_final_reg_req_0;
      addr_of_1001_final_reg_ack_0 <= ack; 
      addr_of_1001_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1000_root_address, dout => iNsTr_125_1002, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1022_final_reg_req_0,addr_of_1022_final_reg_ack_0,sl_one,"addr_of_1022_final_reg ",false,array_obj_ref_1021_root_address,
    false,iNsTr_130_1023);
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1022_final_reg_req_0;
      addr_of_1022_final_reg_ack_0 <= ack; 
      addr_of_1022_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1021_root_address, dout => iNsTr_130_1023, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1043_final_reg_req_0,addr_of_1043_final_reg_ack_0,sl_one,"addr_of_1043_final_reg ",false,array_obj_ref_1042_root_address,
    false,iNsTr_135_1044);
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1043_final_reg_req_0;
      addr_of_1043_final_reg_ack_0 <= ack; 
      addr_of_1043_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1042_root_address, dout => iNsTr_135_1044, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1064_final_reg_req_0,addr_of_1064_final_reg_ack_0,sl_one,"addr_of_1064_final_reg ",false,array_obj_ref_1063_root_address,
    false,iNsTr_140_1065);
    register_block_3 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1064_final_reg_req_0;
      addr_of_1064_final_reg_ack_0 <= ack; 
      addr_of_1064_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1063_root_address, dout => iNsTr_140_1065, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1085_final_reg_req_0,addr_of_1085_final_reg_ack_0,sl_one,"addr_of_1085_final_reg ",false,array_obj_ref_1084_root_address,
    false,iNsTr_145_1086);
    register_block_4 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1085_final_reg_req_0;
      addr_of_1085_final_reg_ack_0 <= ack; 
      addr_of_1085_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1084_root_address, dout => iNsTr_145_1086, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1106_final_reg_req_0,addr_of_1106_final_reg_ack_0,sl_one,"addr_of_1106_final_reg ",false,array_obj_ref_1105_root_address,
    false,iNsTr_150_1107);
    register_block_5 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1106_final_reg_req_0;
      addr_of_1106_final_reg_ack_0 <= ack; 
      addr_of_1106_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1105_root_address, dout => iNsTr_150_1107, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1127_final_reg_req_0,addr_of_1127_final_reg_ack_0,sl_one,"addr_of_1127_final_reg ",false,array_obj_ref_1126_root_address,
    false,iNsTr_155_1128);
    register_block_6 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1127_final_reg_req_0;
      addr_of_1127_final_reg_ack_0 <= ack; 
      addr_of_1127_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1126_root_address, dout => iNsTr_155_1128, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_1148_final_reg_req_0,addr_of_1148_final_reg_ack_0,sl_one,"addr_of_1148_final_reg ",false,array_obj_ref_1147_root_address,
    false,iNsTr_160_1149);
    register_block_7 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_1148_final_reg_req_0;
      addr_of_1148_final_reg_ack_0 <= ack; 
      addr_of_1148_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_1147_root_address, dout => iNsTr_160_1149, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_653_final_reg_req_0,addr_of_653_final_reg_ack_0,sl_one,"addr_of_653_final_reg ",false,array_obj_ref_652_root_address,
    false,iNsTr_44_654);
    register_block_8 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_653_final_reg_req_0;
      addr_of_653_final_reg_ack_0 <= ack; 
      addr_of_653_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_652_root_address, dout => iNsTr_44_654, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_670_final_reg_req_0,addr_of_670_final_reg_ack_0,sl_one,"addr_of_670_final_reg ",false,array_obj_ref_669_root_address,
    false,iNsTr_48_671);
    register_block_9 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_670_final_reg_req_0;
      addr_of_670_final_reg_ack_0 <= ack; 
      addr_of_670_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_669_root_address, dout => iNsTr_48_671, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_696_final_reg_req_0,addr_of_696_final_reg_ack_0,sl_one,"addr_of_696_final_reg ",false,array_obj_ref_695_root_address,
    false,iNsTr_54_697);
    register_block_10 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_696_final_reg_req_0;
      addr_of_696_final_reg_ack_0 <= ack; 
      addr_of_696_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_695_root_address, dout => iNsTr_54_697, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_713_final_reg_req_0,addr_of_713_final_reg_ack_0,sl_one,"addr_of_713_final_reg ",false,array_obj_ref_712_root_address,
    false,iNsTr_58_714);
    register_block_11 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_713_final_reg_req_0;
      addr_of_713_final_reg_ack_0 <= ack; 
      addr_of_713_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_712_root_address, dout => iNsTr_58_714, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_739_final_reg_req_0,addr_of_739_final_reg_ack_0,sl_one,"addr_of_739_final_reg ",false,array_obj_ref_738_root_address,
    false,iNsTr_64_740);
    register_block_12 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_739_final_reg_req_0;
      addr_of_739_final_reg_ack_0 <= ack; 
      addr_of_739_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_738_root_address, dout => iNsTr_64_740, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_756_final_reg_req_0,addr_of_756_final_reg_ack_0,sl_one,"addr_of_756_final_reg ",false,array_obj_ref_755_root_address,
    false,iNsTr_68_757);
    register_block_13 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_756_final_reg_req_0;
      addr_of_756_final_reg_ack_0 <= ack; 
      addr_of_756_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_755_root_address, dout => iNsTr_68_757, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_782_final_reg_req_0,addr_of_782_final_reg_ack_0,sl_one,"addr_of_782_final_reg ",false,array_obj_ref_781_root_address,
    false,iNsTr_74_783);
    register_block_14 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_782_final_reg_req_0;
      addr_of_782_final_reg_ack_0 <= ack; 
      addr_of_782_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_781_root_address, dout => iNsTr_74_783, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_799_final_reg_req_0,addr_of_799_final_reg_ack_0,sl_one,"addr_of_799_final_reg ",false,array_obj_ref_798_root_address,
    false,iNsTr_78_800);
    register_block_15 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_799_final_reg_req_0;
      addr_of_799_final_reg_ack_0 <= ack; 
      addr_of_799_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_798_root_address, dout => iNsTr_78_800, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_825_final_reg_req_0,addr_of_825_final_reg_ack_0,sl_one,"addr_of_825_final_reg ",false,array_obj_ref_824_root_address,
    false,iNsTr_84_826);
    register_block_16 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_825_final_reg_req_0;
      addr_of_825_final_reg_ack_0 <= ack; 
      addr_of_825_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_824_root_address, dout => iNsTr_84_826, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_842_final_reg_req_0,addr_of_842_final_reg_ack_0,sl_one,"addr_of_842_final_reg ",false,array_obj_ref_841_root_address,
    false,iNsTr_88_843);
    register_block_17 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_842_final_reg_req_0;
      addr_of_842_final_reg_ack_0 <= ack; 
      addr_of_842_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_841_root_address, dout => iNsTr_88_843, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_868_final_reg_req_0,addr_of_868_final_reg_ack_0,sl_one,"addr_of_868_final_reg ",false,array_obj_ref_867_root_address,
    false,iNsTr_94_869);
    register_block_18 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_868_final_reg_req_0;
      addr_of_868_final_reg_ack_0 <= ack; 
      addr_of_868_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_867_root_address, dout => iNsTr_94_869, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_885_final_reg_req_0,addr_of_885_final_reg_ack_0,sl_one,"addr_of_885_final_reg ",false,array_obj_ref_884_root_address,
    false,iNsTr_98_886);
    register_block_19 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_885_final_reg_req_0;
      addr_of_885_final_reg_ack_0 <= ack; 
      addr_of_885_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_884_root_address, dout => iNsTr_98_886, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_911_final_reg_req_0,addr_of_911_final_reg_ack_0,sl_one,"addr_of_911_final_reg ",false,array_obj_ref_910_root_address,
    false,iNsTr_104_912);
    register_block_20 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_911_final_reg_req_0;
      addr_of_911_final_reg_ack_0 <= ack; 
      addr_of_911_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_910_root_address, dout => iNsTr_104_912, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_928_final_reg_req_0,addr_of_928_final_reg_ack_0,sl_one,"addr_of_928_final_reg ",false,array_obj_ref_927_root_address,
    false,iNsTr_108_929);
    register_block_21 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_928_final_reg_req_0;
      addr_of_928_final_reg_ack_0 <= ack; 
      addr_of_928_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_927_root_address, dout => iNsTr_108_929, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_954_final_reg_req_0,addr_of_954_final_reg_ack_0,sl_one,"addr_of_954_final_reg ",false,array_obj_ref_953_root_address,
    false,iNsTr_114_955);
    register_block_22 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_954_final_reg_req_0;
      addr_of_954_final_reg_ack_0 <= ack; 
      addr_of_954_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_953_root_address, dout => iNsTr_114_955, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_971_final_reg_req_0,addr_of_971_final_reg_ack_0,sl_one,"addr_of_971_final_reg ",false,array_obj_ref_970_root_address,
    false,iNsTr_118_972);
    register_block_23 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_971_final_reg_req_0;
      addr_of_971_final_reg_ack_0 <= ack; 
      addr_of_971_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_970_root_address, dout => iNsTr_118_972, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1017_inst_req_0,type_cast_1017_inst_ack_0,sl_one,"type_cast_1017_inst ",false,iNsTr_128_1014,
    false,iNsTr_129_1018);
    register_block_24 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1017_inst_req_0;
      type_cast_1017_inst_ack_0 <= ack; 
      type_cast_1017_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_128_1014, dout => iNsTr_129_1018, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1038_inst_req_0,type_cast_1038_inst_ack_0,sl_one,"type_cast_1038_inst ",false,iNsTr_133_1035,
    false,iNsTr_134_1039);
    register_block_25 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1038_inst_req_0;
      type_cast_1038_inst_ack_0 <= ack; 
      type_cast_1038_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_133_1035, dout => iNsTr_134_1039, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1059_inst_req_0,type_cast_1059_inst_ack_0,sl_one,"type_cast_1059_inst ",false,iNsTr_138_1056,
    false,iNsTr_139_1060);
    register_block_26 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1059_inst_req_0;
      type_cast_1059_inst_ack_0 <= ack; 
      type_cast_1059_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_138_1056, dout => iNsTr_139_1060, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1080_inst_req_0,type_cast_1080_inst_ack_0,sl_one,"type_cast_1080_inst ",false,iNsTr_143_1077,
    false,iNsTr_144_1081);
    register_block_27 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1080_inst_req_0;
      type_cast_1080_inst_ack_0 <= ack; 
      type_cast_1080_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_143_1077, dout => iNsTr_144_1081, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1101_inst_req_0,type_cast_1101_inst_ack_0,sl_one,"type_cast_1101_inst ",false,iNsTr_148_1098,
    false,iNsTr_149_1102);
    register_block_28 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1101_inst_req_0;
      type_cast_1101_inst_ack_0 <= ack; 
      type_cast_1101_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_148_1098, dout => iNsTr_149_1102, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1122_inst_req_0,type_cast_1122_inst_ack_0,sl_one,"type_cast_1122_inst ",false,iNsTr_153_1119,
    false,iNsTr_154_1123);
    register_block_29 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1122_inst_req_0;
      type_cast_1122_inst_ack_0 <= ack; 
      type_cast_1122_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_153_1119, dout => iNsTr_154_1123, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1143_inst_req_0,type_cast_1143_inst_ack_0,sl_one,"type_cast_1143_inst ",false,iNsTr_158_1140,
    false,iNsTr_159_1144);
    register_block_30 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1143_inst_req_0;
      type_cast_1143_inst_ack_0 <= ack; 
      type_cast_1143_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_158_1140, dout => iNsTr_159_1144, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1162_inst_req_0,type_cast_1162_inst_ack_0,sl_one,"type_cast_1162_inst ",false,iNsTr_164_1159,
    false,iNsTr_165_1163);
    register_block_31 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1162_inst_req_0;
      type_cast_1162_inst_ack_0 <= ack; 
      type_cast_1162_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_164_1159, dout => iNsTr_165_1163, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_1172_inst_req_0,type_cast_1172_inst_ack_0,sl_one,"type_cast_1172_inst ",false,iNsTr_166_1169,
    false,iNsTr_167_1173);
    register_block_32 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_1172_inst_req_0;
      type_cast_1172_inst_ack_0 <= ack; 
      type_cast_1172_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_166_1169, dout => iNsTr_167_1173, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_471_inst_req_0,type_cast_471_inst_ack_0,sl_one,"type_cast_471_inst ",false,iNsTr_2_468,
    false,iNsTr_3_472);
    register_block_33 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_471_inst_req_0;
      type_cast_471_inst_ack_0 <= ack; 
      type_cast_471_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_2_468, dout => iNsTr_3_472, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_475_inst_req_0,type_cast_475_inst_ack_0,sl_one,"type_cast_475_inst ",false,iNsTr_3_472,
    false,type_cast_475_wire);
    register_block_34 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_475_inst_req_0;
      type_cast_475_inst_ack_0 <= ack; 
      type_cast_475_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_3_472, dout => type_cast_475_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_494_inst_req_0,type_cast_494_inst_ack_0,sl_one,"type_cast_494_inst ",false,iNsTr_7_491,
    false,iNsTr_8_495);
    register_block_35 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_494_inst_req_0;
      type_cast_494_inst_ack_0 <= ack; 
      type_cast_494_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_7_491, dout => iNsTr_8_495, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_504_inst_req_0,type_cast_504_inst_ack_0,sl_one,"type_cast_504_inst ",false,iNsTr_9_501,
    false,iNsTr_10_505);
    register_block_36 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_504_inst_req_0;
      type_cast_504_inst_ack_0 <= ack; 
      type_cast_504_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_9_501, dout => iNsTr_10_505, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_516_inst_req_0,type_cast_516_inst_ack_0,sl_one,"type_cast_516_inst ",false,iNsTr_12_513,
    false,iNsTr_13_517);
    register_block_37 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_516_inst_req_0;
      type_cast_516_inst_ack_0 <= ack; 
      type_cast_516_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_12_513, dout => iNsTr_13_517, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_526_inst_req_0,type_cast_526_inst_ack_0,sl_one,"type_cast_526_inst ",false,iNsTr_14_523,
    false,iNsTr_15_527);
    register_block_38 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_526_inst_req_0;
      type_cast_526_inst_ack_0 <= ack; 
      type_cast_526_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_14_523, dout => iNsTr_15_527, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_538_inst_req_0,type_cast_538_inst_ack_0,sl_one,"type_cast_538_inst ",false,iNsTr_17_535,
    false,iNsTr_18_539);
    register_block_39 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_538_inst_req_0;
      type_cast_538_inst_ack_0 <= ack; 
      type_cast_538_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_17_535, dout => iNsTr_18_539, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_548_inst_req_0,type_cast_548_inst_ack_0,sl_one,"type_cast_548_inst ",false,iNsTr_19_545,
    false,iNsTr_20_549);
    register_block_40 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_548_inst_req_0;
      type_cast_548_inst_ack_0 <= ack; 
      type_cast_548_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_19_545, dout => iNsTr_20_549, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_560_inst_req_0,type_cast_560_inst_ack_0,sl_one,"type_cast_560_inst ",false,iNsTr_22_557,
    false,iNsTr_23_561);
    register_block_41 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_560_inst_req_0;
      type_cast_560_inst_ack_0 <= ack; 
      type_cast_560_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_22_557, dout => iNsTr_23_561, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_570_inst_req_0,type_cast_570_inst_ack_0,sl_one,"type_cast_570_inst ",false,iNsTr_24_567,
    false,iNsTr_25_571);
    register_block_42 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_570_inst_req_0;
      type_cast_570_inst_ack_0 <= ack; 
      type_cast_570_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_24_567, dout => iNsTr_25_571, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_582_inst_req_0,type_cast_582_inst_ack_0,sl_one,"type_cast_582_inst ",false,iNsTr_27_579,
    false,iNsTr_28_583);
    register_block_43 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_582_inst_req_0;
      type_cast_582_inst_ack_0 <= ack; 
      type_cast_582_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_27_579, dout => iNsTr_28_583, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_592_inst_req_0,type_cast_592_inst_ack_0,sl_one,"type_cast_592_inst ",false,iNsTr_29_589,
    false,iNsTr_30_593);
    register_block_44 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_592_inst_req_0;
      type_cast_592_inst_ack_0 <= ack; 
      type_cast_592_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_29_589, dout => iNsTr_30_593, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_604_inst_req_0,type_cast_604_inst_ack_0,sl_one,"type_cast_604_inst ",false,iNsTr_32_601,
    false,iNsTr_33_605);
    register_block_45 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_604_inst_req_0;
      type_cast_604_inst_ack_0 <= ack; 
      type_cast_604_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_32_601, dout => iNsTr_33_605, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_614_inst_req_0,type_cast_614_inst_ack_0,sl_one,"type_cast_614_inst ",false,iNsTr_34_611,
    false,iNsTr_35_615);
    register_block_46 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_614_inst_req_0;
      type_cast_614_inst_ack_0 <= ack; 
      type_cast_614_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_34_611, dout => iNsTr_35_615, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_626_inst_req_0,type_cast_626_inst_ack_0,sl_one,"type_cast_626_inst ",false,iNsTr_37_623,
    false,iNsTr_38_627);
    register_block_47 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_626_inst_req_0;
      type_cast_626_inst_ack_0 <= ack; 
      type_cast_626_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_37_623, dout => iNsTr_38_627, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_636_inst_req_0,type_cast_636_inst_ack_0,sl_one,"type_cast_636_inst ",false,iNsTr_39_633,
    false,iNsTr_40_637);
    register_block_48 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_636_inst_req_0;
      type_cast_636_inst_ack_0 <= ack; 
      type_cast_636_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 8) 
        port map( din => iNsTr_39_633, dout => iNsTr_40_637, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_648_inst_req_0,type_cast_648_inst_ack_0,sl_one,"type_cast_648_inst ",false,iNsTr_42_645,
    false,iNsTr_43_649);
    register_block_49 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_648_inst_req_0;
      type_cast_648_inst_ack_0 <= ack; 
      type_cast_648_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_42_645, dout => iNsTr_43_649, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_665_inst_req_0,type_cast_665_inst_ack_0,sl_one,"type_cast_665_inst ",false,iNsTr_46_662,
    false,iNsTr_47_666);
    register_block_50 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_665_inst_req_0;
      type_cast_665_inst_ack_0 <= ack; 
      type_cast_665_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_46_662, dout => iNsTr_47_666, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_691_inst_req_0,type_cast_691_inst_ack_0,sl_one,"type_cast_691_inst ",false,iNsTr_52_688,
    false,iNsTr_53_692);
    register_block_51 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_691_inst_req_0;
      type_cast_691_inst_ack_0 <= ack; 
      type_cast_691_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_52_688, dout => iNsTr_53_692, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_708_inst_req_0,type_cast_708_inst_ack_0,sl_one,"type_cast_708_inst ",false,iNsTr_56_705,
    false,iNsTr_57_709);
    register_block_52 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_708_inst_req_0;
      type_cast_708_inst_ack_0 <= ack; 
      type_cast_708_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_56_705, dout => iNsTr_57_709, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_734_inst_req_0,type_cast_734_inst_ack_0,sl_one,"type_cast_734_inst ",false,iNsTr_62_731,
    false,iNsTr_63_735);
    register_block_53 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_734_inst_req_0;
      type_cast_734_inst_ack_0 <= ack; 
      type_cast_734_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_62_731, dout => iNsTr_63_735, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_751_inst_req_0,type_cast_751_inst_ack_0,sl_one,"type_cast_751_inst ",false,iNsTr_66_748,
    false,iNsTr_67_752);
    register_block_54 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_751_inst_req_0;
      type_cast_751_inst_ack_0 <= ack; 
      type_cast_751_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_66_748, dout => iNsTr_67_752, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_777_inst_req_0,type_cast_777_inst_ack_0,sl_one,"type_cast_777_inst ",false,iNsTr_72_774,
    false,iNsTr_73_778);
    register_block_55 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_777_inst_req_0;
      type_cast_777_inst_ack_0 <= ack; 
      type_cast_777_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_72_774, dout => iNsTr_73_778, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_794_inst_req_0,type_cast_794_inst_ack_0,sl_one,"type_cast_794_inst ",false,iNsTr_76_791,
    false,iNsTr_77_795);
    register_block_56 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_794_inst_req_0;
      type_cast_794_inst_ack_0 <= ack; 
      type_cast_794_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_76_791, dout => iNsTr_77_795, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_820_inst_req_0,type_cast_820_inst_ack_0,sl_one,"type_cast_820_inst ",false,iNsTr_82_817,
    false,iNsTr_83_821);
    register_block_57 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_820_inst_req_0;
      type_cast_820_inst_ack_0 <= ack; 
      type_cast_820_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_82_817, dout => iNsTr_83_821, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_837_inst_req_0,type_cast_837_inst_ack_0,sl_one,"type_cast_837_inst ",false,iNsTr_86_834,
    false,iNsTr_87_838);
    register_block_58 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_837_inst_req_0;
      type_cast_837_inst_ack_0 <= ack; 
      type_cast_837_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_86_834, dout => iNsTr_87_838, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_863_inst_req_0,type_cast_863_inst_ack_0,sl_one,"type_cast_863_inst ",false,iNsTr_92_860,
    false,iNsTr_93_864);
    register_block_59 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_863_inst_req_0;
      type_cast_863_inst_ack_0 <= ack; 
      type_cast_863_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_92_860, dout => iNsTr_93_864, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_880_inst_req_0,type_cast_880_inst_ack_0,sl_one,"type_cast_880_inst ",false,iNsTr_96_877,
    false,iNsTr_97_881);
    register_block_60 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_880_inst_req_0;
      type_cast_880_inst_ack_0 <= ack; 
      type_cast_880_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_96_877, dout => iNsTr_97_881, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_906_inst_req_0,type_cast_906_inst_ack_0,sl_one,"type_cast_906_inst ",false,iNsTr_102_903,
    false,iNsTr_103_907);
    register_block_61 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_906_inst_req_0;
      type_cast_906_inst_ack_0 <= ack; 
      type_cast_906_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_102_903, dout => iNsTr_103_907, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_923_inst_req_0,type_cast_923_inst_ack_0,sl_one,"type_cast_923_inst ",false,iNsTr_106_920,
    false,iNsTr_107_924);
    register_block_62 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_923_inst_req_0;
      type_cast_923_inst_ack_0 <= ack; 
      type_cast_923_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_106_920, dout => iNsTr_107_924, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_949_inst_req_0,type_cast_949_inst_ack_0,sl_one,"type_cast_949_inst ",false,iNsTr_112_946,
    false,iNsTr_113_950);
    register_block_63 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_949_inst_req_0;
      type_cast_949_inst_ack_0 <= ack; 
      type_cast_949_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_112_946, dout => iNsTr_113_950, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_966_inst_req_0,type_cast_966_inst_ack_0,sl_one,"type_cast_966_inst ",false,iNsTr_116_963,
    false,iNsTr_117_967);
    register_block_64 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_966_inst_req_0;
      type_cast_966_inst_ack_0 <= ack; 
      type_cast_966_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_116_963, dout => iNsTr_117_967, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_996_inst_req_0,type_cast_996_inst_ack_0,sl_one,"type_cast_996_inst ",false,iNsTr_123_993,
    false,iNsTr_124_997);
    register_block_65 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_996_inst_req_0;
      type_cast_996_inst_ack_0 <= ack; 
      type_cast_996_inst: RegisterBase --
        generic map(in_data_width => 8,out_data_width => 32) 
        port map( din => iNsTr_123_993, dout => iNsTr_124_997, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1000_index_0_rename_req_0,array_obj_ref_1000_index_0_rename_ack_0,sl_one,"array_obj_ref_1000_index_0_rename ",false,simple_obj_ref_999_resized,
    false,simple_obj_ref_999_scaled);
    array_obj_ref_1000_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1000_index_0_rename_ack_0 <= array_obj_ref_1000_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_999_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_999_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1000_index_0_resize_req_0,array_obj_ref_1000_index_0_resize_ack_0,sl_one,"array_obj_ref_1000_index_0_resize ",false,iNsTr_124_997,
    false,simple_obj_ref_999_resized);
    array_obj_ref_1000_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1000_index_0_resize_ack_0 <= array_obj_ref_1000_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_124_997;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_999_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1000_offset_inst_req_0,array_obj_ref_1000_offset_inst_ack_0,sl_one,"array_obj_ref_1000_offset_inst ",false,simple_obj_ref_999_scaled,
    false,array_obj_ref_1000_final_offset);
    array_obj_ref_1000_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1000_offset_inst_ack_0 <= array_obj_ref_1000_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_999_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1000_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1000_root_address_inst_req_0,array_obj_ref_1000_root_address_inst_ack_0,sl_one,"array_obj_ref_1000_root_address_inst ",false,array_obj_ref_1000_final_offset,
    false,array_obj_ref_1000_root_address);
    array_obj_ref_1000_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1000_root_address_inst_ack_0 <= array_obj_ref_1000_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1000_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1000_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1021_index_0_rename_req_0,array_obj_ref_1021_index_0_rename_ack_0,sl_one,"array_obj_ref_1021_index_0_rename ",false,simple_obj_ref_1020_resized,
    false,simple_obj_ref_1020_scaled);
    array_obj_ref_1021_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1021_index_0_rename_ack_0 <= array_obj_ref_1021_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1020_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1020_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1021_index_0_resize_req_0,array_obj_ref_1021_index_0_resize_ack_0,sl_one,"array_obj_ref_1021_index_0_resize ",false,iNsTr_129_1018,
    false,simple_obj_ref_1020_resized);
    array_obj_ref_1021_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1021_index_0_resize_ack_0 <= array_obj_ref_1021_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_129_1018;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1020_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1021_offset_inst_req_0,array_obj_ref_1021_offset_inst_ack_0,sl_one,"array_obj_ref_1021_offset_inst ",false,simple_obj_ref_1020_scaled,
    false,array_obj_ref_1021_final_offset);
    array_obj_ref_1021_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1021_offset_inst_ack_0 <= array_obj_ref_1021_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1020_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1021_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1021_root_address_inst_req_0,array_obj_ref_1021_root_address_inst_ack_0,sl_one,"array_obj_ref_1021_root_address_inst ",false,array_obj_ref_1021_final_offset,
    false,array_obj_ref_1021_root_address);
    array_obj_ref_1021_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1021_root_address_inst_ack_0 <= array_obj_ref_1021_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1021_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1021_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1042_index_0_rename_req_0,array_obj_ref_1042_index_0_rename_ack_0,sl_one,"array_obj_ref_1042_index_0_rename ",false,simple_obj_ref_1041_resized,
    false,simple_obj_ref_1041_scaled);
    array_obj_ref_1042_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1042_index_0_rename_ack_0 <= array_obj_ref_1042_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1041_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1041_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1042_index_0_resize_req_0,array_obj_ref_1042_index_0_resize_ack_0,sl_one,"array_obj_ref_1042_index_0_resize ",false,iNsTr_134_1039,
    false,simple_obj_ref_1041_resized);
    array_obj_ref_1042_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1042_index_0_resize_ack_0 <= array_obj_ref_1042_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_134_1039;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1041_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1042_offset_inst_req_0,array_obj_ref_1042_offset_inst_ack_0,sl_one,"array_obj_ref_1042_offset_inst ",false,simple_obj_ref_1041_scaled,
    false,array_obj_ref_1042_final_offset);
    array_obj_ref_1042_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1042_offset_inst_ack_0 <= array_obj_ref_1042_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1041_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1042_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1042_root_address_inst_req_0,array_obj_ref_1042_root_address_inst_ack_0,sl_one,"array_obj_ref_1042_root_address_inst ",false,array_obj_ref_1042_final_offset,
    false,array_obj_ref_1042_root_address);
    array_obj_ref_1042_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1042_root_address_inst_ack_0 <= array_obj_ref_1042_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1042_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1042_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1063_index_0_rename_req_0,array_obj_ref_1063_index_0_rename_ack_0,sl_one,"array_obj_ref_1063_index_0_rename ",false,simple_obj_ref_1062_resized,
    false,simple_obj_ref_1062_scaled);
    array_obj_ref_1063_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1063_index_0_rename_ack_0 <= array_obj_ref_1063_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1062_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1062_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1063_index_0_resize_req_0,array_obj_ref_1063_index_0_resize_ack_0,sl_one,"array_obj_ref_1063_index_0_resize ",false,iNsTr_139_1060,
    false,simple_obj_ref_1062_resized);
    array_obj_ref_1063_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1063_index_0_resize_ack_0 <= array_obj_ref_1063_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_139_1060;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1062_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1063_offset_inst_req_0,array_obj_ref_1063_offset_inst_ack_0,sl_one,"array_obj_ref_1063_offset_inst ",false,simple_obj_ref_1062_scaled,
    false,array_obj_ref_1063_final_offset);
    array_obj_ref_1063_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1063_offset_inst_ack_0 <= array_obj_ref_1063_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1062_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1063_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1063_root_address_inst_req_0,array_obj_ref_1063_root_address_inst_ack_0,sl_one,"array_obj_ref_1063_root_address_inst ",false,array_obj_ref_1063_final_offset,
    false,array_obj_ref_1063_root_address);
    array_obj_ref_1063_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1063_root_address_inst_ack_0 <= array_obj_ref_1063_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1063_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1063_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1084_index_0_rename_req_0,array_obj_ref_1084_index_0_rename_ack_0,sl_one,"array_obj_ref_1084_index_0_rename ",false,simple_obj_ref_1083_resized,
    false,simple_obj_ref_1083_scaled);
    array_obj_ref_1084_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1084_index_0_rename_ack_0 <= array_obj_ref_1084_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1083_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1083_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1084_index_0_resize_req_0,array_obj_ref_1084_index_0_resize_ack_0,sl_one,"array_obj_ref_1084_index_0_resize ",false,iNsTr_144_1081,
    false,simple_obj_ref_1083_resized);
    array_obj_ref_1084_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1084_index_0_resize_ack_0 <= array_obj_ref_1084_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_144_1081;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1083_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1084_offset_inst_req_0,array_obj_ref_1084_offset_inst_ack_0,sl_one,"array_obj_ref_1084_offset_inst ",false,simple_obj_ref_1083_scaled,
    false,array_obj_ref_1084_final_offset);
    array_obj_ref_1084_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1084_offset_inst_ack_0 <= array_obj_ref_1084_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1083_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1084_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1084_root_address_inst_req_0,array_obj_ref_1084_root_address_inst_ack_0,sl_one,"array_obj_ref_1084_root_address_inst ",false,array_obj_ref_1084_final_offset,
    false,array_obj_ref_1084_root_address);
    array_obj_ref_1084_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1084_root_address_inst_ack_0 <= array_obj_ref_1084_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1084_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1084_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1105_index_0_rename_req_0,array_obj_ref_1105_index_0_rename_ack_0,sl_one,"array_obj_ref_1105_index_0_rename ",false,simple_obj_ref_1104_resized,
    false,simple_obj_ref_1104_scaled);
    array_obj_ref_1105_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1105_index_0_rename_ack_0 <= array_obj_ref_1105_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1104_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1104_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1105_index_0_resize_req_0,array_obj_ref_1105_index_0_resize_ack_0,sl_one,"array_obj_ref_1105_index_0_resize ",false,iNsTr_149_1102,
    false,simple_obj_ref_1104_resized);
    array_obj_ref_1105_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1105_index_0_resize_ack_0 <= array_obj_ref_1105_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_149_1102;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1104_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1105_offset_inst_req_0,array_obj_ref_1105_offset_inst_ack_0,sl_one,"array_obj_ref_1105_offset_inst ",false,simple_obj_ref_1104_scaled,
    false,array_obj_ref_1105_final_offset);
    array_obj_ref_1105_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1105_offset_inst_ack_0 <= array_obj_ref_1105_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1104_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1105_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1105_root_address_inst_req_0,array_obj_ref_1105_root_address_inst_ack_0,sl_one,"array_obj_ref_1105_root_address_inst ",false,array_obj_ref_1105_final_offset,
    false,array_obj_ref_1105_root_address);
    array_obj_ref_1105_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1105_root_address_inst_ack_0 <= array_obj_ref_1105_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1105_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1105_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1126_index_0_rename_req_0,array_obj_ref_1126_index_0_rename_ack_0,sl_one,"array_obj_ref_1126_index_0_rename ",false,simple_obj_ref_1125_resized,
    false,simple_obj_ref_1125_scaled);
    array_obj_ref_1126_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1126_index_0_rename_ack_0 <= array_obj_ref_1126_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1125_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1125_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1126_index_0_resize_req_0,array_obj_ref_1126_index_0_resize_ack_0,sl_one,"array_obj_ref_1126_index_0_resize ",false,iNsTr_154_1123,
    false,simple_obj_ref_1125_resized);
    array_obj_ref_1126_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1126_index_0_resize_ack_0 <= array_obj_ref_1126_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_154_1123;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1125_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1126_offset_inst_req_0,array_obj_ref_1126_offset_inst_ack_0,sl_one,"array_obj_ref_1126_offset_inst ",false,simple_obj_ref_1125_scaled,
    false,array_obj_ref_1126_final_offset);
    array_obj_ref_1126_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1126_offset_inst_ack_0 <= array_obj_ref_1126_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1125_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1126_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1126_root_address_inst_req_0,array_obj_ref_1126_root_address_inst_ack_0,sl_one,"array_obj_ref_1126_root_address_inst ",false,array_obj_ref_1126_final_offset,
    false,array_obj_ref_1126_root_address);
    array_obj_ref_1126_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1126_root_address_inst_ack_0 <= array_obj_ref_1126_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1126_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1126_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1147_index_0_rename_req_0,array_obj_ref_1147_index_0_rename_ack_0,sl_one,"array_obj_ref_1147_index_0_rename ",false,simple_obj_ref_1146_resized,
    false,simple_obj_ref_1146_scaled);
    array_obj_ref_1147_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1147_index_0_rename_ack_0 <= array_obj_ref_1147_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_1146_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_1146_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1147_index_0_resize_req_0,array_obj_ref_1147_index_0_resize_ack_0,sl_one,"array_obj_ref_1147_index_0_resize ",false,iNsTr_159_1144,
    false,simple_obj_ref_1146_resized);
    array_obj_ref_1147_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1147_index_0_resize_ack_0 <= array_obj_ref_1147_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_159_1144;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_1146_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1147_offset_inst_req_0,array_obj_ref_1147_offset_inst_ack_0,sl_one,"array_obj_ref_1147_offset_inst ",false,simple_obj_ref_1146_scaled,
    false,array_obj_ref_1147_final_offset);
    array_obj_ref_1147_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1147_offset_inst_ack_0 <= array_obj_ref_1147_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_1146_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1147_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_1147_root_address_inst_req_0,array_obj_ref_1147_root_address_inst_ack_0,sl_one,"array_obj_ref_1147_root_address_inst ",false,array_obj_ref_1147_final_offset,
    false,array_obj_ref_1147_root_address);
    array_obj_ref_1147_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_1147_root_address_inst_ack_0 <= array_obj_ref_1147_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_1147_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_1147_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_652_index_0_rename_req_0,array_obj_ref_652_index_0_rename_ack_0,sl_one,"array_obj_ref_652_index_0_rename ",false,simple_obj_ref_651_resized,
    false,simple_obj_ref_651_scaled);
    array_obj_ref_652_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_652_index_0_rename_ack_0 <= array_obj_ref_652_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_651_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_651_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_652_index_0_resize_req_0,array_obj_ref_652_index_0_resize_ack_0,sl_one,"array_obj_ref_652_index_0_resize ",false,iNsTr_43_649,
    false,simple_obj_ref_651_resized);
    array_obj_ref_652_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_652_index_0_resize_ack_0 <= array_obj_ref_652_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_43_649;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_651_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_652_offset_inst_req_0,array_obj_ref_652_offset_inst_ack_0,sl_one,"array_obj_ref_652_offset_inst ",false,simple_obj_ref_651_scaled,
    false,array_obj_ref_652_final_offset);
    array_obj_ref_652_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_652_offset_inst_ack_0 <= array_obj_ref_652_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_651_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_652_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_652_root_address_inst_req_0,array_obj_ref_652_root_address_inst_ack_0,sl_one,"array_obj_ref_652_root_address_inst ",false,array_obj_ref_652_final_offset,
    false,array_obj_ref_652_root_address);
    array_obj_ref_652_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_652_root_address_inst_ack_0 <= array_obj_ref_652_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_652_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_652_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_669_index_0_rename_req_0,array_obj_ref_669_index_0_rename_ack_0,sl_one,"array_obj_ref_669_index_0_rename ",false,simple_obj_ref_668_resized,
    false,simple_obj_ref_668_scaled);
    array_obj_ref_669_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_669_index_0_rename_ack_0 <= array_obj_ref_669_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_668_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_668_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_669_index_0_resize_req_0,array_obj_ref_669_index_0_resize_ack_0,sl_one,"array_obj_ref_669_index_0_resize ",false,iNsTr_47_666,
    false,simple_obj_ref_668_resized);
    array_obj_ref_669_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_669_index_0_resize_ack_0 <= array_obj_ref_669_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_47_666;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_668_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_669_offset_inst_req_0,array_obj_ref_669_offset_inst_ack_0,sl_one,"array_obj_ref_669_offset_inst ",false,simple_obj_ref_668_scaled,
    false,array_obj_ref_669_final_offset);
    array_obj_ref_669_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_669_offset_inst_ack_0 <= array_obj_ref_669_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_668_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_669_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_669_root_address_inst_req_0,array_obj_ref_669_root_address_inst_ack_0,sl_one,"array_obj_ref_669_root_address_inst ",false,array_obj_ref_669_final_offset,
    false,array_obj_ref_669_root_address);
    array_obj_ref_669_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_669_root_address_inst_ack_0 <= array_obj_ref_669_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_669_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_669_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_695_index_0_rename_req_0,array_obj_ref_695_index_0_rename_ack_0,sl_one,"array_obj_ref_695_index_0_rename ",false,simple_obj_ref_694_resized,
    false,simple_obj_ref_694_scaled);
    array_obj_ref_695_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_695_index_0_rename_ack_0 <= array_obj_ref_695_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_694_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_694_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_695_index_0_resize_req_0,array_obj_ref_695_index_0_resize_ack_0,sl_one,"array_obj_ref_695_index_0_resize ",false,iNsTr_53_692,
    false,simple_obj_ref_694_resized);
    array_obj_ref_695_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_695_index_0_resize_ack_0 <= array_obj_ref_695_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_53_692;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_694_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_695_offset_inst_req_0,array_obj_ref_695_offset_inst_ack_0,sl_one,"array_obj_ref_695_offset_inst ",false,simple_obj_ref_694_scaled,
    false,array_obj_ref_695_final_offset);
    array_obj_ref_695_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_695_offset_inst_ack_0 <= array_obj_ref_695_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_694_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_695_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_695_root_address_inst_req_0,array_obj_ref_695_root_address_inst_ack_0,sl_one,"array_obj_ref_695_root_address_inst ",false,array_obj_ref_695_final_offset,
    false,array_obj_ref_695_root_address);
    array_obj_ref_695_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_695_root_address_inst_ack_0 <= array_obj_ref_695_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_695_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_695_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_712_index_0_rename_req_0,array_obj_ref_712_index_0_rename_ack_0,sl_one,"array_obj_ref_712_index_0_rename ",false,simple_obj_ref_711_resized,
    false,simple_obj_ref_711_scaled);
    array_obj_ref_712_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_712_index_0_rename_ack_0 <= array_obj_ref_712_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_711_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_711_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_712_index_0_resize_req_0,array_obj_ref_712_index_0_resize_ack_0,sl_one,"array_obj_ref_712_index_0_resize ",false,iNsTr_57_709,
    false,simple_obj_ref_711_resized);
    array_obj_ref_712_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_712_index_0_resize_ack_0 <= array_obj_ref_712_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_57_709;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_711_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_712_offset_inst_req_0,array_obj_ref_712_offset_inst_ack_0,sl_one,"array_obj_ref_712_offset_inst ",false,simple_obj_ref_711_scaled,
    false,array_obj_ref_712_final_offset);
    array_obj_ref_712_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_712_offset_inst_ack_0 <= array_obj_ref_712_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_711_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_712_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_712_root_address_inst_req_0,array_obj_ref_712_root_address_inst_ack_0,sl_one,"array_obj_ref_712_root_address_inst ",false,array_obj_ref_712_final_offset,
    false,array_obj_ref_712_root_address);
    array_obj_ref_712_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_712_root_address_inst_ack_0 <= array_obj_ref_712_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_712_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_712_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_738_index_0_rename_req_0,array_obj_ref_738_index_0_rename_ack_0,sl_one,"array_obj_ref_738_index_0_rename ",false,simple_obj_ref_737_resized,
    false,simple_obj_ref_737_scaled);
    array_obj_ref_738_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_738_index_0_rename_ack_0 <= array_obj_ref_738_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_737_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_737_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_738_index_0_resize_req_0,array_obj_ref_738_index_0_resize_ack_0,sl_one,"array_obj_ref_738_index_0_resize ",false,iNsTr_63_735,
    false,simple_obj_ref_737_resized);
    array_obj_ref_738_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_738_index_0_resize_ack_0 <= array_obj_ref_738_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_63_735;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_737_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_738_offset_inst_req_0,array_obj_ref_738_offset_inst_ack_0,sl_one,"array_obj_ref_738_offset_inst ",false,simple_obj_ref_737_scaled,
    false,array_obj_ref_738_final_offset);
    array_obj_ref_738_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_738_offset_inst_ack_0 <= array_obj_ref_738_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_737_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_738_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_738_root_address_inst_req_0,array_obj_ref_738_root_address_inst_ack_0,sl_one,"array_obj_ref_738_root_address_inst ",false,array_obj_ref_738_final_offset,
    false,array_obj_ref_738_root_address);
    array_obj_ref_738_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_738_root_address_inst_ack_0 <= array_obj_ref_738_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_738_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_738_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_755_index_0_rename_req_0,array_obj_ref_755_index_0_rename_ack_0,sl_one,"array_obj_ref_755_index_0_rename ",false,simple_obj_ref_754_resized,
    false,simple_obj_ref_754_scaled);
    array_obj_ref_755_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_755_index_0_rename_ack_0 <= array_obj_ref_755_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_754_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_754_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_755_index_0_resize_req_0,array_obj_ref_755_index_0_resize_ack_0,sl_one,"array_obj_ref_755_index_0_resize ",false,iNsTr_67_752,
    false,simple_obj_ref_754_resized);
    array_obj_ref_755_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_755_index_0_resize_ack_0 <= array_obj_ref_755_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_67_752;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_754_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_755_offset_inst_req_0,array_obj_ref_755_offset_inst_ack_0,sl_one,"array_obj_ref_755_offset_inst ",false,simple_obj_ref_754_scaled,
    false,array_obj_ref_755_final_offset);
    array_obj_ref_755_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_755_offset_inst_ack_0 <= array_obj_ref_755_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_754_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_755_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_755_root_address_inst_req_0,array_obj_ref_755_root_address_inst_ack_0,sl_one,"array_obj_ref_755_root_address_inst ",false,array_obj_ref_755_final_offset,
    false,array_obj_ref_755_root_address);
    array_obj_ref_755_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_755_root_address_inst_ack_0 <= array_obj_ref_755_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_755_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_755_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_781_index_0_rename_req_0,array_obj_ref_781_index_0_rename_ack_0,sl_one,"array_obj_ref_781_index_0_rename ",false,simple_obj_ref_780_resized,
    false,simple_obj_ref_780_scaled);
    array_obj_ref_781_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_781_index_0_rename_ack_0 <= array_obj_ref_781_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_780_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_780_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_781_index_0_resize_req_0,array_obj_ref_781_index_0_resize_ack_0,sl_one,"array_obj_ref_781_index_0_resize ",false,iNsTr_73_778,
    false,simple_obj_ref_780_resized);
    array_obj_ref_781_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_781_index_0_resize_ack_0 <= array_obj_ref_781_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_73_778;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_780_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_781_offset_inst_req_0,array_obj_ref_781_offset_inst_ack_0,sl_one,"array_obj_ref_781_offset_inst ",false,simple_obj_ref_780_scaled,
    false,array_obj_ref_781_final_offset);
    array_obj_ref_781_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_781_offset_inst_ack_0 <= array_obj_ref_781_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_780_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_781_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_781_root_address_inst_req_0,array_obj_ref_781_root_address_inst_ack_0,sl_one,"array_obj_ref_781_root_address_inst ",false,array_obj_ref_781_final_offset,
    false,array_obj_ref_781_root_address);
    array_obj_ref_781_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_781_root_address_inst_ack_0 <= array_obj_ref_781_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_781_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_781_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_798_index_0_rename_req_0,array_obj_ref_798_index_0_rename_ack_0,sl_one,"array_obj_ref_798_index_0_rename ",false,simple_obj_ref_797_resized,
    false,simple_obj_ref_797_scaled);
    array_obj_ref_798_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_798_index_0_rename_ack_0 <= array_obj_ref_798_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_797_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_797_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_798_index_0_resize_req_0,array_obj_ref_798_index_0_resize_ack_0,sl_one,"array_obj_ref_798_index_0_resize ",false,iNsTr_77_795,
    false,simple_obj_ref_797_resized);
    array_obj_ref_798_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_798_index_0_resize_ack_0 <= array_obj_ref_798_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_77_795;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_797_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_798_offset_inst_req_0,array_obj_ref_798_offset_inst_ack_0,sl_one,"array_obj_ref_798_offset_inst ",false,simple_obj_ref_797_scaled,
    false,array_obj_ref_798_final_offset);
    array_obj_ref_798_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_798_offset_inst_ack_0 <= array_obj_ref_798_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_797_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_798_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_798_root_address_inst_req_0,array_obj_ref_798_root_address_inst_ack_0,sl_one,"array_obj_ref_798_root_address_inst ",false,array_obj_ref_798_final_offset,
    false,array_obj_ref_798_root_address);
    array_obj_ref_798_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_798_root_address_inst_ack_0 <= array_obj_ref_798_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_798_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_798_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_824_index_0_rename_req_0,array_obj_ref_824_index_0_rename_ack_0,sl_one,"array_obj_ref_824_index_0_rename ",false,simple_obj_ref_823_resized,
    false,simple_obj_ref_823_scaled);
    array_obj_ref_824_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_824_index_0_rename_ack_0 <= array_obj_ref_824_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_823_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_823_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_824_index_0_resize_req_0,array_obj_ref_824_index_0_resize_ack_0,sl_one,"array_obj_ref_824_index_0_resize ",false,iNsTr_83_821,
    false,simple_obj_ref_823_resized);
    array_obj_ref_824_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_824_index_0_resize_ack_0 <= array_obj_ref_824_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_83_821;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_823_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_824_offset_inst_req_0,array_obj_ref_824_offset_inst_ack_0,sl_one,"array_obj_ref_824_offset_inst ",false,simple_obj_ref_823_scaled,
    false,array_obj_ref_824_final_offset);
    array_obj_ref_824_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_824_offset_inst_ack_0 <= array_obj_ref_824_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_823_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_824_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_824_root_address_inst_req_0,array_obj_ref_824_root_address_inst_ack_0,sl_one,"array_obj_ref_824_root_address_inst ",false,array_obj_ref_824_final_offset,
    false,array_obj_ref_824_root_address);
    array_obj_ref_824_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_824_root_address_inst_ack_0 <= array_obj_ref_824_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_824_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_824_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_841_index_0_rename_req_0,array_obj_ref_841_index_0_rename_ack_0,sl_one,"array_obj_ref_841_index_0_rename ",false,simple_obj_ref_840_resized,
    false,simple_obj_ref_840_scaled);
    array_obj_ref_841_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_841_index_0_rename_ack_0 <= array_obj_ref_841_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_840_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_840_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_841_index_0_resize_req_0,array_obj_ref_841_index_0_resize_ack_0,sl_one,"array_obj_ref_841_index_0_resize ",false,iNsTr_87_838,
    false,simple_obj_ref_840_resized);
    array_obj_ref_841_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_841_index_0_resize_ack_0 <= array_obj_ref_841_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_87_838;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_840_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_841_offset_inst_req_0,array_obj_ref_841_offset_inst_ack_0,sl_one,"array_obj_ref_841_offset_inst ",false,simple_obj_ref_840_scaled,
    false,array_obj_ref_841_final_offset);
    array_obj_ref_841_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_841_offset_inst_ack_0 <= array_obj_ref_841_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_840_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_841_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_841_root_address_inst_req_0,array_obj_ref_841_root_address_inst_ack_0,sl_one,"array_obj_ref_841_root_address_inst ",false,array_obj_ref_841_final_offset,
    false,array_obj_ref_841_root_address);
    array_obj_ref_841_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_841_root_address_inst_ack_0 <= array_obj_ref_841_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_841_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_841_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_867_index_0_rename_req_0,array_obj_ref_867_index_0_rename_ack_0,sl_one,"array_obj_ref_867_index_0_rename ",false,simple_obj_ref_866_resized,
    false,simple_obj_ref_866_scaled);
    array_obj_ref_867_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_867_index_0_rename_ack_0 <= array_obj_ref_867_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_866_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_866_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_867_index_0_resize_req_0,array_obj_ref_867_index_0_resize_ack_0,sl_one,"array_obj_ref_867_index_0_resize ",false,iNsTr_93_864,
    false,simple_obj_ref_866_resized);
    array_obj_ref_867_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_867_index_0_resize_ack_0 <= array_obj_ref_867_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_93_864;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_866_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_867_offset_inst_req_0,array_obj_ref_867_offset_inst_ack_0,sl_one,"array_obj_ref_867_offset_inst ",false,simple_obj_ref_866_scaled,
    false,array_obj_ref_867_final_offset);
    array_obj_ref_867_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_867_offset_inst_ack_0 <= array_obj_ref_867_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_866_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_867_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_867_root_address_inst_req_0,array_obj_ref_867_root_address_inst_ack_0,sl_one,"array_obj_ref_867_root_address_inst ",false,array_obj_ref_867_final_offset,
    false,array_obj_ref_867_root_address);
    array_obj_ref_867_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_867_root_address_inst_ack_0 <= array_obj_ref_867_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_867_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_867_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_884_index_0_rename_req_0,array_obj_ref_884_index_0_rename_ack_0,sl_one,"array_obj_ref_884_index_0_rename ",false,simple_obj_ref_883_resized,
    false,simple_obj_ref_883_scaled);
    array_obj_ref_884_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_884_index_0_rename_ack_0 <= array_obj_ref_884_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_883_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_883_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_884_index_0_resize_req_0,array_obj_ref_884_index_0_resize_ack_0,sl_one,"array_obj_ref_884_index_0_resize ",false,iNsTr_97_881,
    false,simple_obj_ref_883_resized);
    array_obj_ref_884_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_884_index_0_resize_ack_0 <= array_obj_ref_884_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_97_881;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_883_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_884_offset_inst_req_0,array_obj_ref_884_offset_inst_ack_0,sl_one,"array_obj_ref_884_offset_inst ",false,simple_obj_ref_883_scaled,
    false,array_obj_ref_884_final_offset);
    array_obj_ref_884_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_884_offset_inst_ack_0 <= array_obj_ref_884_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_883_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_884_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_884_root_address_inst_req_0,array_obj_ref_884_root_address_inst_ack_0,sl_one,"array_obj_ref_884_root_address_inst ",false,array_obj_ref_884_final_offset,
    false,array_obj_ref_884_root_address);
    array_obj_ref_884_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_884_root_address_inst_ack_0 <= array_obj_ref_884_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_884_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_884_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_910_index_0_rename_req_0,array_obj_ref_910_index_0_rename_ack_0,sl_one,"array_obj_ref_910_index_0_rename ",false,simple_obj_ref_909_resized,
    false,simple_obj_ref_909_scaled);
    array_obj_ref_910_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_910_index_0_rename_ack_0 <= array_obj_ref_910_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_909_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_909_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_910_index_0_resize_req_0,array_obj_ref_910_index_0_resize_ack_0,sl_one,"array_obj_ref_910_index_0_resize ",false,iNsTr_103_907,
    false,simple_obj_ref_909_resized);
    array_obj_ref_910_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_910_index_0_resize_ack_0 <= array_obj_ref_910_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_103_907;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_909_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_910_offset_inst_req_0,array_obj_ref_910_offset_inst_ack_0,sl_one,"array_obj_ref_910_offset_inst ",false,simple_obj_ref_909_scaled,
    false,array_obj_ref_910_final_offset);
    array_obj_ref_910_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_910_offset_inst_ack_0 <= array_obj_ref_910_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_909_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_910_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_910_root_address_inst_req_0,array_obj_ref_910_root_address_inst_ack_0,sl_one,"array_obj_ref_910_root_address_inst ",false,array_obj_ref_910_final_offset,
    false,array_obj_ref_910_root_address);
    array_obj_ref_910_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_910_root_address_inst_ack_0 <= array_obj_ref_910_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_910_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_910_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_927_index_0_rename_req_0,array_obj_ref_927_index_0_rename_ack_0,sl_one,"array_obj_ref_927_index_0_rename ",false,simple_obj_ref_926_resized,
    false,simple_obj_ref_926_scaled);
    array_obj_ref_927_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_927_index_0_rename_ack_0 <= array_obj_ref_927_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_926_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_926_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_927_index_0_resize_req_0,array_obj_ref_927_index_0_resize_ack_0,sl_one,"array_obj_ref_927_index_0_resize ",false,iNsTr_107_924,
    false,simple_obj_ref_926_resized);
    array_obj_ref_927_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_927_index_0_resize_ack_0 <= array_obj_ref_927_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_107_924;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_926_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_927_offset_inst_req_0,array_obj_ref_927_offset_inst_ack_0,sl_one,"array_obj_ref_927_offset_inst ",false,simple_obj_ref_926_scaled,
    false,array_obj_ref_927_final_offset);
    array_obj_ref_927_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_927_offset_inst_ack_0 <= array_obj_ref_927_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_926_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_927_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_927_root_address_inst_req_0,array_obj_ref_927_root_address_inst_ack_0,sl_one,"array_obj_ref_927_root_address_inst ",false,array_obj_ref_927_final_offset,
    false,array_obj_ref_927_root_address);
    array_obj_ref_927_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_927_root_address_inst_ack_0 <= array_obj_ref_927_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_927_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_927_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_953_index_0_rename_req_0,array_obj_ref_953_index_0_rename_ack_0,sl_one,"array_obj_ref_953_index_0_rename ",false,simple_obj_ref_952_resized,
    false,simple_obj_ref_952_scaled);
    array_obj_ref_953_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_953_index_0_rename_ack_0 <= array_obj_ref_953_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_952_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_952_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_953_index_0_resize_req_0,array_obj_ref_953_index_0_resize_ack_0,sl_one,"array_obj_ref_953_index_0_resize ",false,iNsTr_113_950,
    false,simple_obj_ref_952_resized);
    array_obj_ref_953_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_953_index_0_resize_ack_0 <= array_obj_ref_953_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_113_950;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_952_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_953_offset_inst_req_0,array_obj_ref_953_offset_inst_ack_0,sl_one,"array_obj_ref_953_offset_inst ",false,simple_obj_ref_952_scaled,
    false,array_obj_ref_953_final_offset);
    array_obj_ref_953_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_953_offset_inst_ack_0 <= array_obj_ref_953_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_952_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_953_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_953_root_address_inst_req_0,array_obj_ref_953_root_address_inst_ack_0,sl_one,"array_obj_ref_953_root_address_inst ",false,array_obj_ref_953_final_offset,
    false,array_obj_ref_953_root_address);
    array_obj_ref_953_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_953_root_address_inst_ack_0 <= array_obj_ref_953_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_953_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_953_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_970_index_0_rename_req_0,array_obj_ref_970_index_0_rename_ack_0,sl_one,"array_obj_ref_970_index_0_rename ",false,simple_obj_ref_969_resized,
    false,simple_obj_ref_969_scaled);
    array_obj_ref_970_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_970_index_0_rename_ack_0 <= array_obj_ref_970_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_969_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_969_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_970_index_0_resize_req_0,array_obj_ref_970_index_0_resize_ack_0,sl_one,"array_obj_ref_970_index_0_resize ",false,iNsTr_117_967,
    false,simple_obj_ref_969_resized);
    array_obj_ref_970_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_970_index_0_resize_ack_0 <= array_obj_ref_970_index_0_resize_req_0;
      in_aggregated_sig <= iNsTr_117_967;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_969_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_970_offset_inst_req_0,array_obj_ref_970_offset_inst_ack_0,sl_one,"array_obj_ref_970_offset_inst ",false,simple_obj_ref_969_scaled,
    false,array_obj_ref_970_final_offset);
    array_obj_ref_970_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_970_offset_inst_ack_0 <= array_obj_ref_970_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_969_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_970_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_970_root_address_inst_req_0,array_obj_ref_970_root_address_inst_ack_0,sl_one,"array_obj_ref_970_root_address_inst ",false,array_obj_ref_970_final_offset,
    false,array_obj_ref_970_root_address);
    array_obj_ref_970_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_970_root_address_inst_ack_0 <= array_obj_ref_970_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_970_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_970_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1004_addr_0_req_0,ptr_deref_1004_addr_0_ack_0,sl_one,"ptr_deref_1004_addr_0 ",false,ptr_deref_1004_root_address,
    false,ptr_deref_1004_word_address_0);
    ptr_deref_1004_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1004_addr_0_ack_0 <= ptr_deref_1004_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1004_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1004_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1004_base_resize_req_0,ptr_deref_1004_base_resize_ack_0,sl_one,"ptr_deref_1004_base_resize ",false,iNsTr_125_1002,
    false,ptr_deref_1004_resized_base_address);
    ptr_deref_1004_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1004_base_resize_ack_0 <= ptr_deref_1004_base_resize_req_0;
      in_aggregated_sig <= iNsTr_125_1002;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1004_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1004_gather_scatter_req_0,ptr_deref_1004_gather_scatter_ack_0,sl_one,"ptr_deref_1004_gather_scatter ",false,iNsTr_122_989,
    false,ptr_deref_1004_data_0);
    ptr_deref_1004_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1004_gather_scatter_ack_0 <= ptr_deref_1004_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_122_989;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1004_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1004_root_address_inst_req_0,ptr_deref_1004_root_address_inst_ack_0,sl_one,"ptr_deref_1004_root_address_inst ",false,ptr_deref_1004_resized_base_address,
    false,ptr_deref_1004_root_address);
    ptr_deref_1004_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1004_root_address_inst_ack_0 <= ptr_deref_1004_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1004_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1004_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1009_addr_0_req_0,ptr_deref_1009_addr_0_ack_0,sl_one,"ptr_deref_1009_addr_0 ",false,ptr_deref_1009_root_address,
    false,ptr_deref_1009_word_address_0);
    ptr_deref_1009_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1009_addr_0_ack_0 <= ptr_deref_1009_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1009_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1009_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1009_base_resize_req_0,ptr_deref_1009_base_resize_ack_0,sl_one,"ptr_deref_1009_base_resize ",false,c1_433,
    false,ptr_deref_1009_resized_base_address);
    ptr_deref_1009_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1009_base_resize_ack_0 <= ptr_deref_1009_base_resize_req_0;
      in_aggregated_sig <= c1_433;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1009_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1009_gather_scatter_req_0,ptr_deref_1009_gather_scatter_ack_0,sl_one,"ptr_deref_1009_gather_scatter ",false,ptr_deref_1009_data_0,
    false,iNsTr_127_1010);
    ptr_deref_1009_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1009_gather_scatter_ack_0 <= ptr_deref_1009_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1009_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_127_1010 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1009_root_address_inst_req_0,ptr_deref_1009_root_address_inst_ack_0,sl_one,"ptr_deref_1009_root_address_inst ",false,ptr_deref_1009_resized_base_address,
    false,ptr_deref_1009_root_address);
    ptr_deref_1009_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1009_root_address_inst_ack_0 <= ptr_deref_1009_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1009_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1009_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1013_addr_0_req_0,ptr_deref_1013_addr_0_ack_0,sl_one,"ptr_deref_1013_addr_0 ",false,ptr_deref_1013_root_address,
    false,ptr_deref_1013_word_address_0);
    ptr_deref_1013_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1013_addr_0_ack_0 <= ptr_deref_1013_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1013_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1013_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1013_base_resize_req_0,ptr_deref_1013_base_resize_ack_0,sl_one,"ptr_deref_1013_base_resize ",false,I1_401,
    false,ptr_deref_1013_resized_base_address);
    ptr_deref_1013_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1013_base_resize_ack_0 <= ptr_deref_1013_base_resize_req_0;
      in_aggregated_sig <= I1_401;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1013_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1013_gather_scatter_req_0,ptr_deref_1013_gather_scatter_ack_0,sl_one,"ptr_deref_1013_gather_scatter ",false,ptr_deref_1013_data_0,
    false,iNsTr_128_1014);
    ptr_deref_1013_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1013_gather_scatter_ack_0 <= ptr_deref_1013_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1013_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_128_1014 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1013_root_address_inst_req_0,ptr_deref_1013_root_address_inst_ack_0,sl_one,"ptr_deref_1013_root_address_inst ",false,ptr_deref_1013_resized_base_address,
    false,ptr_deref_1013_root_address);
    ptr_deref_1013_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1013_root_address_inst_ack_0 <= ptr_deref_1013_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1013_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1013_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1025_addr_0_req_0,ptr_deref_1025_addr_0_ack_0,sl_one,"ptr_deref_1025_addr_0 ",false,ptr_deref_1025_root_address,
    false,ptr_deref_1025_word_address_0);
    ptr_deref_1025_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1025_addr_0_ack_0 <= ptr_deref_1025_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1025_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1025_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1025_base_resize_req_0,ptr_deref_1025_base_resize_ack_0,sl_one,"ptr_deref_1025_base_resize ",false,iNsTr_130_1023,
    false,ptr_deref_1025_resized_base_address);
    ptr_deref_1025_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1025_base_resize_ack_0 <= ptr_deref_1025_base_resize_req_0;
      in_aggregated_sig <= iNsTr_130_1023;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1025_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1025_gather_scatter_req_0,ptr_deref_1025_gather_scatter_ack_0,sl_one,"ptr_deref_1025_gather_scatter ",false,iNsTr_127_1010,
    false,ptr_deref_1025_data_0);
    ptr_deref_1025_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1025_gather_scatter_ack_0 <= ptr_deref_1025_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_127_1010;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1025_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1025_root_address_inst_req_0,ptr_deref_1025_root_address_inst_ack_0,sl_one,"ptr_deref_1025_root_address_inst ",false,ptr_deref_1025_resized_base_address,
    false,ptr_deref_1025_root_address);
    ptr_deref_1025_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1025_root_address_inst_ack_0 <= ptr_deref_1025_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1025_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1025_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1030_addr_0_req_0,ptr_deref_1030_addr_0_ack_0,sl_one,"ptr_deref_1030_addr_0 ",false,ptr_deref_1030_root_address,
    false,ptr_deref_1030_word_address_0);
    ptr_deref_1030_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1030_addr_0_ack_0 <= ptr_deref_1030_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1030_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1030_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1030_base_resize_req_0,ptr_deref_1030_base_resize_ack_0,sl_one,"ptr_deref_1030_base_resize ",false,c2_437,
    false,ptr_deref_1030_resized_base_address);
    ptr_deref_1030_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1030_base_resize_ack_0 <= ptr_deref_1030_base_resize_req_0;
      in_aggregated_sig <= c2_437;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1030_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1030_gather_scatter_req_0,ptr_deref_1030_gather_scatter_ack_0,sl_one,"ptr_deref_1030_gather_scatter ",false,ptr_deref_1030_data_0,
    false,iNsTr_132_1031);
    ptr_deref_1030_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1030_gather_scatter_ack_0 <= ptr_deref_1030_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1030_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_132_1031 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1030_root_address_inst_req_0,ptr_deref_1030_root_address_inst_ack_0,sl_one,"ptr_deref_1030_root_address_inst ",false,ptr_deref_1030_resized_base_address,
    false,ptr_deref_1030_root_address);
    ptr_deref_1030_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1030_root_address_inst_ack_0 <= ptr_deref_1030_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1030_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1030_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1034_addr_0_req_0,ptr_deref_1034_addr_0_ack_0,sl_one,"ptr_deref_1034_addr_0 ",false,ptr_deref_1034_root_address,
    false,ptr_deref_1034_word_address_0);
    ptr_deref_1034_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1034_addr_0_ack_0 <= ptr_deref_1034_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1034_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1034_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1034_base_resize_req_0,ptr_deref_1034_base_resize_ack_0,sl_one,"ptr_deref_1034_base_resize ",false,I2_405,
    false,ptr_deref_1034_resized_base_address);
    ptr_deref_1034_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1034_base_resize_ack_0 <= ptr_deref_1034_base_resize_req_0;
      in_aggregated_sig <= I2_405;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1034_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1034_gather_scatter_req_0,ptr_deref_1034_gather_scatter_ack_0,sl_one,"ptr_deref_1034_gather_scatter ",false,ptr_deref_1034_data_0,
    false,iNsTr_133_1035);
    ptr_deref_1034_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1034_gather_scatter_ack_0 <= ptr_deref_1034_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1034_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_133_1035 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1034_root_address_inst_req_0,ptr_deref_1034_root_address_inst_ack_0,sl_one,"ptr_deref_1034_root_address_inst ",false,ptr_deref_1034_resized_base_address,
    false,ptr_deref_1034_root_address);
    ptr_deref_1034_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1034_root_address_inst_ack_0 <= ptr_deref_1034_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1034_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1034_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1046_addr_0_req_0,ptr_deref_1046_addr_0_ack_0,sl_one,"ptr_deref_1046_addr_0 ",false,ptr_deref_1046_root_address,
    false,ptr_deref_1046_word_address_0);
    ptr_deref_1046_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1046_addr_0_ack_0 <= ptr_deref_1046_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1046_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1046_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1046_base_resize_req_0,ptr_deref_1046_base_resize_ack_0,sl_one,"ptr_deref_1046_base_resize ",false,iNsTr_135_1044,
    false,ptr_deref_1046_resized_base_address);
    ptr_deref_1046_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1046_base_resize_ack_0 <= ptr_deref_1046_base_resize_req_0;
      in_aggregated_sig <= iNsTr_135_1044;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1046_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1046_gather_scatter_req_0,ptr_deref_1046_gather_scatter_ack_0,sl_one,"ptr_deref_1046_gather_scatter ",false,iNsTr_132_1031,
    false,ptr_deref_1046_data_0);
    ptr_deref_1046_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1046_gather_scatter_ack_0 <= ptr_deref_1046_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_132_1031;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1046_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1046_root_address_inst_req_0,ptr_deref_1046_root_address_inst_ack_0,sl_one,"ptr_deref_1046_root_address_inst ",false,ptr_deref_1046_resized_base_address,
    false,ptr_deref_1046_root_address);
    ptr_deref_1046_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1046_root_address_inst_ack_0 <= ptr_deref_1046_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1046_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1046_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1051_addr_0_req_0,ptr_deref_1051_addr_0_ack_0,sl_one,"ptr_deref_1051_addr_0 ",false,ptr_deref_1051_root_address,
    false,ptr_deref_1051_word_address_0);
    ptr_deref_1051_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1051_addr_0_ack_0 <= ptr_deref_1051_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1051_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1051_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1051_base_resize_req_0,ptr_deref_1051_base_resize_ack_0,sl_one,"ptr_deref_1051_base_resize ",false,c3_441,
    false,ptr_deref_1051_resized_base_address);
    ptr_deref_1051_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1051_base_resize_ack_0 <= ptr_deref_1051_base_resize_req_0;
      in_aggregated_sig <= c3_441;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1051_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1051_gather_scatter_req_0,ptr_deref_1051_gather_scatter_ack_0,sl_one,"ptr_deref_1051_gather_scatter ",false,ptr_deref_1051_data_0,
    false,iNsTr_137_1052);
    ptr_deref_1051_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1051_gather_scatter_ack_0 <= ptr_deref_1051_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1051_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_137_1052 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1051_root_address_inst_req_0,ptr_deref_1051_root_address_inst_ack_0,sl_one,"ptr_deref_1051_root_address_inst ",false,ptr_deref_1051_resized_base_address,
    false,ptr_deref_1051_root_address);
    ptr_deref_1051_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1051_root_address_inst_ack_0 <= ptr_deref_1051_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1051_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1051_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1055_addr_0_req_0,ptr_deref_1055_addr_0_ack_0,sl_one,"ptr_deref_1055_addr_0 ",false,ptr_deref_1055_root_address,
    false,ptr_deref_1055_word_address_0);
    ptr_deref_1055_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1055_addr_0_ack_0 <= ptr_deref_1055_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1055_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1055_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1055_base_resize_req_0,ptr_deref_1055_base_resize_ack_0,sl_one,"ptr_deref_1055_base_resize ",false,I3_409,
    false,ptr_deref_1055_resized_base_address);
    ptr_deref_1055_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1055_base_resize_ack_0 <= ptr_deref_1055_base_resize_req_0;
      in_aggregated_sig <= I3_409;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1055_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1055_gather_scatter_req_0,ptr_deref_1055_gather_scatter_ack_0,sl_one,"ptr_deref_1055_gather_scatter ",false,ptr_deref_1055_data_0,
    false,iNsTr_138_1056);
    ptr_deref_1055_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1055_gather_scatter_ack_0 <= ptr_deref_1055_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1055_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_138_1056 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1055_root_address_inst_req_0,ptr_deref_1055_root_address_inst_ack_0,sl_one,"ptr_deref_1055_root_address_inst ",false,ptr_deref_1055_resized_base_address,
    false,ptr_deref_1055_root_address);
    ptr_deref_1055_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1055_root_address_inst_ack_0 <= ptr_deref_1055_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1055_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1055_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1067_addr_0_req_0,ptr_deref_1067_addr_0_ack_0,sl_one,"ptr_deref_1067_addr_0 ",false,ptr_deref_1067_root_address,
    false,ptr_deref_1067_word_address_0);
    ptr_deref_1067_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1067_addr_0_ack_0 <= ptr_deref_1067_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1067_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1067_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1067_base_resize_req_0,ptr_deref_1067_base_resize_ack_0,sl_one,"ptr_deref_1067_base_resize ",false,iNsTr_140_1065,
    false,ptr_deref_1067_resized_base_address);
    ptr_deref_1067_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1067_base_resize_ack_0 <= ptr_deref_1067_base_resize_req_0;
      in_aggregated_sig <= iNsTr_140_1065;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1067_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1067_gather_scatter_req_0,ptr_deref_1067_gather_scatter_ack_0,sl_one,"ptr_deref_1067_gather_scatter ",false,iNsTr_137_1052,
    false,ptr_deref_1067_data_0);
    ptr_deref_1067_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1067_gather_scatter_ack_0 <= ptr_deref_1067_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_137_1052;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1067_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1067_root_address_inst_req_0,ptr_deref_1067_root_address_inst_ack_0,sl_one,"ptr_deref_1067_root_address_inst ",false,ptr_deref_1067_resized_base_address,
    false,ptr_deref_1067_root_address);
    ptr_deref_1067_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1067_root_address_inst_ack_0 <= ptr_deref_1067_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1067_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1067_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1072_addr_0_req_0,ptr_deref_1072_addr_0_ack_0,sl_one,"ptr_deref_1072_addr_0 ",false,ptr_deref_1072_root_address,
    false,ptr_deref_1072_word_address_0);
    ptr_deref_1072_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1072_addr_0_ack_0 <= ptr_deref_1072_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1072_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1072_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1072_base_resize_req_0,ptr_deref_1072_base_resize_ack_0,sl_one,"ptr_deref_1072_base_resize ",false,c4_445,
    false,ptr_deref_1072_resized_base_address);
    ptr_deref_1072_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1072_base_resize_ack_0 <= ptr_deref_1072_base_resize_req_0;
      in_aggregated_sig <= c4_445;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1072_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1072_gather_scatter_req_0,ptr_deref_1072_gather_scatter_ack_0,sl_one,"ptr_deref_1072_gather_scatter ",false,ptr_deref_1072_data_0,
    false,iNsTr_142_1073);
    ptr_deref_1072_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1072_gather_scatter_ack_0 <= ptr_deref_1072_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1072_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_142_1073 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1072_root_address_inst_req_0,ptr_deref_1072_root_address_inst_ack_0,sl_one,"ptr_deref_1072_root_address_inst ",false,ptr_deref_1072_resized_base_address,
    false,ptr_deref_1072_root_address);
    ptr_deref_1072_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1072_root_address_inst_ack_0 <= ptr_deref_1072_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1072_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1072_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1076_addr_0_req_0,ptr_deref_1076_addr_0_ack_0,sl_one,"ptr_deref_1076_addr_0 ",false,ptr_deref_1076_root_address,
    false,ptr_deref_1076_word_address_0);
    ptr_deref_1076_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1076_addr_0_ack_0 <= ptr_deref_1076_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1076_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1076_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1076_base_resize_req_0,ptr_deref_1076_base_resize_ack_0,sl_one,"ptr_deref_1076_base_resize ",false,I4_413,
    false,ptr_deref_1076_resized_base_address);
    ptr_deref_1076_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1076_base_resize_ack_0 <= ptr_deref_1076_base_resize_req_0;
      in_aggregated_sig <= I4_413;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1076_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1076_gather_scatter_req_0,ptr_deref_1076_gather_scatter_ack_0,sl_one,"ptr_deref_1076_gather_scatter ",false,ptr_deref_1076_data_0,
    false,iNsTr_143_1077);
    ptr_deref_1076_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1076_gather_scatter_ack_0 <= ptr_deref_1076_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1076_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_143_1077 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1076_root_address_inst_req_0,ptr_deref_1076_root_address_inst_ack_0,sl_one,"ptr_deref_1076_root_address_inst ",false,ptr_deref_1076_resized_base_address,
    false,ptr_deref_1076_root_address);
    ptr_deref_1076_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1076_root_address_inst_ack_0 <= ptr_deref_1076_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1076_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1076_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1088_addr_0_req_0,ptr_deref_1088_addr_0_ack_0,sl_one,"ptr_deref_1088_addr_0 ",false,ptr_deref_1088_root_address,
    false,ptr_deref_1088_word_address_0);
    ptr_deref_1088_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1088_addr_0_ack_0 <= ptr_deref_1088_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1088_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1088_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1088_base_resize_req_0,ptr_deref_1088_base_resize_ack_0,sl_one,"ptr_deref_1088_base_resize ",false,iNsTr_145_1086,
    false,ptr_deref_1088_resized_base_address);
    ptr_deref_1088_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1088_base_resize_ack_0 <= ptr_deref_1088_base_resize_req_0;
      in_aggregated_sig <= iNsTr_145_1086;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1088_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1088_gather_scatter_req_0,ptr_deref_1088_gather_scatter_ack_0,sl_one,"ptr_deref_1088_gather_scatter ",false,iNsTr_142_1073,
    false,ptr_deref_1088_data_0);
    ptr_deref_1088_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1088_gather_scatter_ack_0 <= ptr_deref_1088_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_142_1073;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1088_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1088_root_address_inst_req_0,ptr_deref_1088_root_address_inst_ack_0,sl_one,"ptr_deref_1088_root_address_inst ",false,ptr_deref_1088_resized_base_address,
    false,ptr_deref_1088_root_address);
    ptr_deref_1088_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1088_root_address_inst_ack_0 <= ptr_deref_1088_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1088_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1088_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1093_addr_0_req_0,ptr_deref_1093_addr_0_ack_0,sl_one,"ptr_deref_1093_addr_0 ",false,ptr_deref_1093_root_address,
    false,ptr_deref_1093_word_address_0);
    ptr_deref_1093_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1093_addr_0_ack_0 <= ptr_deref_1093_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1093_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1093_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1093_base_resize_req_0,ptr_deref_1093_base_resize_ack_0,sl_one,"ptr_deref_1093_base_resize ",false,c5_449,
    false,ptr_deref_1093_resized_base_address);
    ptr_deref_1093_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1093_base_resize_ack_0 <= ptr_deref_1093_base_resize_req_0;
      in_aggregated_sig <= c5_449;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1093_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1093_gather_scatter_req_0,ptr_deref_1093_gather_scatter_ack_0,sl_one,"ptr_deref_1093_gather_scatter ",false,ptr_deref_1093_data_0,
    false,iNsTr_147_1094);
    ptr_deref_1093_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1093_gather_scatter_ack_0 <= ptr_deref_1093_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1093_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_147_1094 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1093_root_address_inst_req_0,ptr_deref_1093_root_address_inst_ack_0,sl_one,"ptr_deref_1093_root_address_inst ",false,ptr_deref_1093_resized_base_address,
    false,ptr_deref_1093_root_address);
    ptr_deref_1093_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1093_root_address_inst_ack_0 <= ptr_deref_1093_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1093_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1093_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1097_addr_0_req_0,ptr_deref_1097_addr_0_ack_0,sl_one,"ptr_deref_1097_addr_0 ",false,ptr_deref_1097_root_address,
    false,ptr_deref_1097_word_address_0);
    ptr_deref_1097_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1097_addr_0_ack_0 <= ptr_deref_1097_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1097_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1097_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1097_base_resize_req_0,ptr_deref_1097_base_resize_ack_0,sl_one,"ptr_deref_1097_base_resize ",false,I5_417,
    false,ptr_deref_1097_resized_base_address);
    ptr_deref_1097_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1097_base_resize_ack_0 <= ptr_deref_1097_base_resize_req_0;
      in_aggregated_sig <= I5_417;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1097_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1097_gather_scatter_req_0,ptr_deref_1097_gather_scatter_ack_0,sl_one,"ptr_deref_1097_gather_scatter ",false,ptr_deref_1097_data_0,
    false,iNsTr_148_1098);
    ptr_deref_1097_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1097_gather_scatter_ack_0 <= ptr_deref_1097_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1097_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_148_1098 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1097_root_address_inst_req_0,ptr_deref_1097_root_address_inst_ack_0,sl_one,"ptr_deref_1097_root_address_inst ",false,ptr_deref_1097_resized_base_address,
    false,ptr_deref_1097_root_address);
    ptr_deref_1097_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1097_root_address_inst_ack_0 <= ptr_deref_1097_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1097_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1097_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1109_addr_0_req_0,ptr_deref_1109_addr_0_ack_0,sl_one,"ptr_deref_1109_addr_0 ",false,ptr_deref_1109_root_address,
    false,ptr_deref_1109_word_address_0);
    ptr_deref_1109_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1109_addr_0_ack_0 <= ptr_deref_1109_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1109_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1109_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1109_base_resize_req_0,ptr_deref_1109_base_resize_ack_0,sl_one,"ptr_deref_1109_base_resize ",false,iNsTr_150_1107,
    false,ptr_deref_1109_resized_base_address);
    ptr_deref_1109_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1109_base_resize_ack_0 <= ptr_deref_1109_base_resize_req_0;
      in_aggregated_sig <= iNsTr_150_1107;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1109_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1109_gather_scatter_req_0,ptr_deref_1109_gather_scatter_ack_0,sl_one,"ptr_deref_1109_gather_scatter ",false,iNsTr_147_1094,
    false,ptr_deref_1109_data_0);
    ptr_deref_1109_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1109_gather_scatter_ack_0 <= ptr_deref_1109_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_147_1094;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1109_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1109_root_address_inst_req_0,ptr_deref_1109_root_address_inst_ack_0,sl_one,"ptr_deref_1109_root_address_inst ",false,ptr_deref_1109_resized_base_address,
    false,ptr_deref_1109_root_address);
    ptr_deref_1109_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1109_root_address_inst_ack_0 <= ptr_deref_1109_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1109_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1109_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1114_addr_0_req_0,ptr_deref_1114_addr_0_ack_0,sl_one,"ptr_deref_1114_addr_0 ",false,ptr_deref_1114_root_address,
    false,ptr_deref_1114_word_address_0);
    ptr_deref_1114_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1114_addr_0_ack_0 <= ptr_deref_1114_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1114_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1114_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1114_base_resize_req_0,ptr_deref_1114_base_resize_ack_0,sl_one,"ptr_deref_1114_base_resize ",false,c6_453,
    false,ptr_deref_1114_resized_base_address);
    ptr_deref_1114_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1114_base_resize_ack_0 <= ptr_deref_1114_base_resize_req_0;
      in_aggregated_sig <= c6_453;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1114_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1114_gather_scatter_req_0,ptr_deref_1114_gather_scatter_ack_0,sl_one,"ptr_deref_1114_gather_scatter ",false,ptr_deref_1114_data_0,
    false,iNsTr_152_1115);
    ptr_deref_1114_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1114_gather_scatter_ack_0 <= ptr_deref_1114_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1114_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_152_1115 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1114_root_address_inst_req_0,ptr_deref_1114_root_address_inst_ack_0,sl_one,"ptr_deref_1114_root_address_inst ",false,ptr_deref_1114_resized_base_address,
    false,ptr_deref_1114_root_address);
    ptr_deref_1114_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1114_root_address_inst_ack_0 <= ptr_deref_1114_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1114_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1114_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1118_addr_0_req_0,ptr_deref_1118_addr_0_ack_0,sl_one,"ptr_deref_1118_addr_0 ",false,ptr_deref_1118_root_address,
    false,ptr_deref_1118_word_address_0);
    ptr_deref_1118_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1118_addr_0_ack_0 <= ptr_deref_1118_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1118_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1118_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1118_base_resize_req_0,ptr_deref_1118_base_resize_ack_0,sl_one,"ptr_deref_1118_base_resize ",false,I6_421,
    false,ptr_deref_1118_resized_base_address);
    ptr_deref_1118_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1118_base_resize_ack_0 <= ptr_deref_1118_base_resize_req_0;
      in_aggregated_sig <= I6_421;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1118_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1118_gather_scatter_req_0,ptr_deref_1118_gather_scatter_ack_0,sl_one,"ptr_deref_1118_gather_scatter ",false,ptr_deref_1118_data_0,
    false,iNsTr_153_1119);
    ptr_deref_1118_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1118_gather_scatter_ack_0 <= ptr_deref_1118_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1118_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_153_1119 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1118_root_address_inst_req_0,ptr_deref_1118_root_address_inst_ack_0,sl_one,"ptr_deref_1118_root_address_inst ",false,ptr_deref_1118_resized_base_address,
    false,ptr_deref_1118_root_address);
    ptr_deref_1118_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1118_root_address_inst_ack_0 <= ptr_deref_1118_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1118_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1118_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1130_addr_0_req_0,ptr_deref_1130_addr_0_ack_0,sl_one,"ptr_deref_1130_addr_0 ",false,ptr_deref_1130_root_address,
    false,ptr_deref_1130_word_address_0);
    ptr_deref_1130_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1130_addr_0_ack_0 <= ptr_deref_1130_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1130_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1130_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1130_base_resize_req_0,ptr_deref_1130_base_resize_ack_0,sl_one,"ptr_deref_1130_base_resize ",false,iNsTr_155_1128,
    false,ptr_deref_1130_resized_base_address);
    ptr_deref_1130_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1130_base_resize_ack_0 <= ptr_deref_1130_base_resize_req_0;
      in_aggregated_sig <= iNsTr_155_1128;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1130_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1130_gather_scatter_req_0,ptr_deref_1130_gather_scatter_ack_0,sl_one,"ptr_deref_1130_gather_scatter ",false,iNsTr_152_1115,
    false,ptr_deref_1130_data_0);
    ptr_deref_1130_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1130_gather_scatter_ack_0 <= ptr_deref_1130_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_152_1115;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1130_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1130_root_address_inst_req_0,ptr_deref_1130_root_address_inst_ack_0,sl_one,"ptr_deref_1130_root_address_inst ",false,ptr_deref_1130_resized_base_address,
    false,ptr_deref_1130_root_address);
    ptr_deref_1130_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1130_root_address_inst_ack_0 <= ptr_deref_1130_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1130_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1130_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1135_addr_0_req_0,ptr_deref_1135_addr_0_ack_0,sl_one,"ptr_deref_1135_addr_0 ",false,ptr_deref_1135_root_address,
    false,ptr_deref_1135_word_address_0);
    ptr_deref_1135_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1135_addr_0_ack_0 <= ptr_deref_1135_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1135_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1135_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1135_base_resize_req_0,ptr_deref_1135_base_resize_ack_0,sl_one,"ptr_deref_1135_base_resize ",false,c7_457,
    false,ptr_deref_1135_resized_base_address);
    ptr_deref_1135_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1135_base_resize_ack_0 <= ptr_deref_1135_base_resize_req_0;
      in_aggregated_sig <= c7_457;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1135_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1135_gather_scatter_req_0,ptr_deref_1135_gather_scatter_ack_0,sl_one,"ptr_deref_1135_gather_scatter ",false,ptr_deref_1135_data_0,
    false,iNsTr_157_1136);
    ptr_deref_1135_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1135_gather_scatter_ack_0 <= ptr_deref_1135_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1135_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_157_1136 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1135_root_address_inst_req_0,ptr_deref_1135_root_address_inst_ack_0,sl_one,"ptr_deref_1135_root_address_inst ",false,ptr_deref_1135_resized_base_address,
    false,ptr_deref_1135_root_address);
    ptr_deref_1135_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1135_root_address_inst_ack_0 <= ptr_deref_1135_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1135_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1135_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1139_addr_0_req_0,ptr_deref_1139_addr_0_ack_0,sl_one,"ptr_deref_1139_addr_0 ",false,ptr_deref_1139_root_address,
    false,ptr_deref_1139_word_address_0);
    ptr_deref_1139_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1139_addr_0_ack_0 <= ptr_deref_1139_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1139_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1139_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1139_base_resize_req_0,ptr_deref_1139_base_resize_ack_0,sl_one,"ptr_deref_1139_base_resize ",false,I7_425,
    false,ptr_deref_1139_resized_base_address);
    ptr_deref_1139_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1139_base_resize_ack_0 <= ptr_deref_1139_base_resize_req_0;
      in_aggregated_sig <= I7_425;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1139_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1139_gather_scatter_req_0,ptr_deref_1139_gather_scatter_ack_0,sl_one,"ptr_deref_1139_gather_scatter ",false,ptr_deref_1139_data_0,
    false,iNsTr_158_1140);
    ptr_deref_1139_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1139_gather_scatter_ack_0 <= ptr_deref_1139_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1139_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_158_1140 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1139_root_address_inst_req_0,ptr_deref_1139_root_address_inst_ack_0,sl_one,"ptr_deref_1139_root_address_inst ",false,ptr_deref_1139_resized_base_address,
    false,ptr_deref_1139_root_address);
    ptr_deref_1139_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1139_root_address_inst_ack_0 <= ptr_deref_1139_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1139_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1139_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1151_addr_0_req_0,ptr_deref_1151_addr_0_ack_0,sl_one,"ptr_deref_1151_addr_0 ",false,ptr_deref_1151_root_address,
    false,ptr_deref_1151_word_address_0);
    ptr_deref_1151_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1151_addr_0_ack_0 <= ptr_deref_1151_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1151_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1151_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1151_base_resize_req_0,ptr_deref_1151_base_resize_ack_0,sl_one,"ptr_deref_1151_base_resize ",false,iNsTr_160_1149,
    false,ptr_deref_1151_resized_base_address);
    ptr_deref_1151_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1151_base_resize_ack_0 <= ptr_deref_1151_base_resize_req_0;
      in_aggregated_sig <= iNsTr_160_1149;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_1151_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1151_gather_scatter_req_0,ptr_deref_1151_gather_scatter_ack_0,sl_one,"ptr_deref_1151_gather_scatter ",false,iNsTr_157_1136,
    false,ptr_deref_1151_data_0);
    ptr_deref_1151_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_1151_gather_scatter_ack_0 <= ptr_deref_1151_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_157_1136;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1151_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1151_root_address_inst_req_0,ptr_deref_1151_root_address_inst_ack_0,sl_one,"ptr_deref_1151_root_address_inst ",false,ptr_deref_1151_resized_base_address,
    false,ptr_deref_1151_root_address);
    ptr_deref_1151_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_1151_root_address_inst_ack_0 <= ptr_deref_1151_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1151_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1151_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1158_addr_0_req_0,ptr_deref_1158_addr_0_ack_0,sl_one,"ptr_deref_1158_addr_0 ",false,ptr_deref_1158_root_address,
    false,ptr_deref_1158_word_address_0);
    ptr_deref_1158_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1158_addr_0_ack_0 <= ptr_deref_1158_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1158_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1158_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1158_base_resize_req_0,ptr_deref_1158_base_resize_ack_0,sl_one,"ptr_deref_1158_base_resize ",false,I_397,
    false,ptr_deref_1158_resized_base_address);
    ptr_deref_1158_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1158_base_resize_ack_0 <= ptr_deref_1158_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1158_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1158_gather_scatter_req_0,ptr_deref_1158_gather_scatter_ack_0,sl_one,"ptr_deref_1158_gather_scatter ",false,ptr_deref_1158_data_0,
    false,iNsTr_164_1159);
    ptr_deref_1158_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1158_gather_scatter_ack_0 <= ptr_deref_1158_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_1158_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_164_1159 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1158_root_address_inst_req_0,ptr_deref_1158_root_address_inst_ack_0,sl_one,"ptr_deref_1158_root_address_inst ",false,ptr_deref_1158_resized_base_address,
    false,ptr_deref_1158_root_address);
    ptr_deref_1158_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1158_root_address_inst_ack_0 <= ptr_deref_1158_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1158_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1158_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1175_addr_0_req_0,ptr_deref_1175_addr_0_ack_0,sl_one,"ptr_deref_1175_addr_0 ",false,ptr_deref_1175_root_address,
    false,ptr_deref_1175_word_address_0);
    ptr_deref_1175_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1175_addr_0_ack_0 <= ptr_deref_1175_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_1175_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1175_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1175_base_resize_req_0,ptr_deref_1175_base_resize_ack_0,sl_one,"ptr_deref_1175_base_resize ",false,I_397,
    false,ptr_deref_1175_resized_base_address);
    ptr_deref_1175_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1175_base_resize_ack_0 <= ptr_deref_1175_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_1175_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1175_gather_scatter_req_0,ptr_deref_1175_gather_scatter_ack_0,sl_one,"ptr_deref_1175_gather_scatter ",false,iNsTr_167_1173,
    false,ptr_deref_1175_data_0);
    ptr_deref_1175_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_1175_gather_scatter_ack_0 <= ptr_deref_1175_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_167_1173;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1175_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_1175_root_address_inst_req_0,ptr_deref_1175_root_address_inst_ack_0,sl_one,"ptr_deref_1175_root_address_inst ",false,ptr_deref_1175_resized_base_address,
    false,ptr_deref_1175_root_address);
    ptr_deref_1175_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_1175_root_address_inst_ack_0 <= ptr_deref_1175_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_1175_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_1175_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_459_addr_0_req_0,ptr_deref_459_addr_0_ack_0,sl_one,"ptr_deref_459_addr_0 ",false,ptr_deref_459_root_address,
    false,ptr_deref_459_word_address_0);
    ptr_deref_459_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_459_addr_0_ack_0 <= ptr_deref_459_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_459_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_459_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_459_base_resize_req_0,ptr_deref_459_base_resize_ack_0,sl_one,"ptr_deref_459_base_resize ",false,I_397,
    false,ptr_deref_459_resized_base_address);
    ptr_deref_459_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_459_base_resize_ack_0 <= ptr_deref_459_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_459_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_459_gather_scatter_req_0,ptr_deref_459_gather_scatter_ack_0,sl_one,"ptr_deref_459_gather_scatter ",false,type_cast_461_wire_constant,
    false,ptr_deref_459_data_0);
    ptr_deref_459_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_459_gather_scatter_ack_0 <= ptr_deref_459_gather_scatter_req_0;
      in_aggregated_sig <= type_cast_461_wire_constant;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_459_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_459_root_address_inst_req_0,ptr_deref_459_root_address_inst_ack_0,sl_one,"ptr_deref_459_root_address_inst ",false,ptr_deref_459_resized_base_address,
    false,ptr_deref_459_root_address);
    ptr_deref_459_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_459_root_address_inst_ack_0 <= ptr_deref_459_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_459_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_459_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_467_addr_0_req_0,ptr_deref_467_addr_0_ack_0,sl_one,"ptr_deref_467_addr_0 ",false,ptr_deref_467_root_address,
    false,ptr_deref_467_word_address_0);
    ptr_deref_467_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_467_addr_0_ack_0 <= ptr_deref_467_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_467_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_467_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_467_base_resize_req_0,ptr_deref_467_base_resize_ack_0,sl_one,"ptr_deref_467_base_resize ",false,I_397,
    false,ptr_deref_467_resized_base_address);
    ptr_deref_467_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_467_base_resize_ack_0 <= ptr_deref_467_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_467_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_467_gather_scatter_req_0,ptr_deref_467_gather_scatter_ack_0,sl_one,"ptr_deref_467_gather_scatter ",false,ptr_deref_467_data_0,
    false,iNsTr_2_468);
    ptr_deref_467_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_467_gather_scatter_ack_0 <= ptr_deref_467_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_467_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_2_468 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_467_root_address_inst_req_0,ptr_deref_467_root_address_inst_ack_0,sl_one,"ptr_deref_467_root_address_inst ",false,ptr_deref_467_resized_base_address,
    false,ptr_deref_467_root_address);
    ptr_deref_467_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_467_root_address_inst_ack_0 <= ptr_deref_467_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_467_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_467_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_490_addr_0_req_0,ptr_deref_490_addr_0_ack_0,sl_one,"ptr_deref_490_addr_0 ",false,ptr_deref_490_root_address,
    false,ptr_deref_490_word_address_0);
    ptr_deref_490_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_490_addr_0_ack_0 <= ptr_deref_490_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_490_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_490_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_490_base_resize_req_0,ptr_deref_490_base_resize_ack_0,sl_one,"ptr_deref_490_base_resize ",false,I_397,
    false,ptr_deref_490_resized_base_address);
    ptr_deref_490_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_490_base_resize_ack_0 <= ptr_deref_490_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_490_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_490_gather_scatter_req_0,ptr_deref_490_gather_scatter_ack_0,sl_one,"ptr_deref_490_gather_scatter ",false,ptr_deref_490_data_0,
    false,iNsTr_7_491);
    ptr_deref_490_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_490_gather_scatter_ack_0 <= ptr_deref_490_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_490_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_7_491 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_490_root_address_inst_req_0,ptr_deref_490_root_address_inst_ack_0,sl_one,"ptr_deref_490_root_address_inst ",false,ptr_deref_490_resized_base_address,
    false,ptr_deref_490_root_address);
    ptr_deref_490_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_490_root_address_inst_ack_0 <= ptr_deref_490_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_490_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_490_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_507_addr_0_req_0,ptr_deref_507_addr_0_ack_0,sl_one,"ptr_deref_507_addr_0 ",false,ptr_deref_507_root_address,
    false,ptr_deref_507_word_address_0);
    ptr_deref_507_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_507_addr_0_ack_0 <= ptr_deref_507_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_507_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_507_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_507_base_resize_req_0,ptr_deref_507_base_resize_ack_0,sl_one,"ptr_deref_507_base_resize ",false,I1_401,
    false,ptr_deref_507_resized_base_address);
    ptr_deref_507_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_507_base_resize_ack_0 <= ptr_deref_507_base_resize_req_0;
      in_aggregated_sig <= I1_401;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_507_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_507_gather_scatter_req_0,ptr_deref_507_gather_scatter_ack_0,sl_one,"ptr_deref_507_gather_scatter ",false,iNsTr_10_505,
    false,ptr_deref_507_data_0);
    ptr_deref_507_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_507_gather_scatter_ack_0 <= ptr_deref_507_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_10_505;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_507_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_507_root_address_inst_req_0,ptr_deref_507_root_address_inst_ack_0,sl_one,"ptr_deref_507_root_address_inst ",false,ptr_deref_507_resized_base_address,
    false,ptr_deref_507_root_address);
    ptr_deref_507_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_507_root_address_inst_ack_0 <= ptr_deref_507_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_507_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_507_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_512_addr_0_req_0,ptr_deref_512_addr_0_ack_0,sl_one,"ptr_deref_512_addr_0 ",false,ptr_deref_512_root_address,
    false,ptr_deref_512_word_address_0);
    ptr_deref_512_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_512_addr_0_ack_0 <= ptr_deref_512_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_512_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_512_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_512_base_resize_req_0,ptr_deref_512_base_resize_ack_0,sl_one,"ptr_deref_512_base_resize ",false,I_397,
    false,ptr_deref_512_resized_base_address);
    ptr_deref_512_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_512_base_resize_ack_0 <= ptr_deref_512_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_512_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_512_gather_scatter_req_0,ptr_deref_512_gather_scatter_ack_0,sl_one,"ptr_deref_512_gather_scatter ",false,ptr_deref_512_data_0,
    false,iNsTr_12_513);
    ptr_deref_512_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_512_gather_scatter_ack_0 <= ptr_deref_512_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_512_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_12_513 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_512_root_address_inst_req_0,ptr_deref_512_root_address_inst_ack_0,sl_one,"ptr_deref_512_root_address_inst ",false,ptr_deref_512_resized_base_address,
    false,ptr_deref_512_root_address);
    ptr_deref_512_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_512_root_address_inst_ack_0 <= ptr_deref_512_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_512_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_512_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_529_addr_0_req_0,ptr_deref_529_addr_0_ack_0,sl_one,"ptr_deref_529_addr_0 ",false,ptr_deref_529_root_address,
    false,ptr_deref_529_word_address_0);
    ptr_deref_529_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_529_addr_0_ack_0 <= ptr_deref_529_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_529_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_529_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_529_base_resize_req_0,ptr_deref_529_base_resize_ack_0,sl_one,"ptr_deref_529_base_resize ",false,I2_405,
    false,ptr_deref_529_resized_base_address);
    ptr_deref_529_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_529_base_resize_ack_0 <= ptr_deref_529_base_resize_req_0;
      in_aggregated_sig <= I2_405;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_529_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_529_gather_scatter_req_0,ptr_deref_529_gather_scatter_ack_0,sl_one,"ptr_deref_529_gather_scatter ",false,iNsTr_15_527,
    false,ptr_deref_529_data_0);
    ptr_deref_529_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_529_gather_scatter_ack_0 <= ptr_deref_529_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_15_527;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_529_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_529_root_address_inst_req_0,ptr_deref_529_root_address_inst_ack_0,sl_one,"ptr_deref_529_root_address_inst ",false,ptr_deref_529_resized_base_address,
    false,ptr_deref_529_root_address);
    ptr_deref_529_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_529_root_address_inst_ack_0 <= ptr_deref_529_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_529_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_529_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_534_addr_0_req_0,ptr_deref_534_addr_0_ack_0,sl_one,"ptr_deref_534_addr_0 ",false,ptr_deref_534_root_address,
    false,ptr_deref_534_word_address_0);
    ptr_deref_534_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_534_addr_0_ack_0 <= ptr_deref_534_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_534_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_534_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_534_base_resize_req_0,ptr_deref_534_base_resize_ack_0,sl_one,"ptr_deref_534_base_resize ",false,I_397,
    false,ptr_deref_534_resized_base_address);
    ptr_deref_534_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_534_base_resize_ack_0 <= ptr_deref_534_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_534_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_534_gather_scatter_req_0,ptr_deref_534_gather_scatter_ack_0,sl_one,"ptr_deref_534_gather_scatter ",false,ptr_deref_534_data_0,
    false,iNsTr_17_535);
    ptr_deref_534_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_534_gather_scatter_ack_0 <= ptr_deref_534_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_534_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_17_535 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_534_root_address_inst_req_0,ptr_deref_534_root_address_inst_ack_0,sl_one,"ptr_deref_534_root_address_inst ",false,ptr_deref_534_resized_base_address,
    false,ptr_deref_534_root_address);
    ptr_deref_534_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_534_root_address_inst_ack_0 <= ptr_deref_534_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_534_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_534_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_551_addr_0_req_0,ptr_deref_551_addr_0_ack_0,sl_one,"ptr_deref_551_addr_0 ",false,ptr_deref_551_root_address,
    false,ptr_deref_551_word_address_0);
    ptr_deref_551_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_551_addr_0_ack_0 <= ptr_deref_551_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_551_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_551_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_551_base_resize_req_0,ptr_deref_551_base_resize_ack_0,sl_one,"ptr_deref_551_base_resize ",false,I3_409,
    false,ptr_deref_551_resized_base_address);
    ptr_deref_551_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_551_base_resize_ack_0 <= ptr_deref_551_base_resize_req_0;
      in_aggregated_sig <= I3_409;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_551_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_551_gather_scatter_req_0,ptr_deref_551_gather_scatter_ack_0,sl_one,"ptr_deref_551_gather_scatter ",false,iNsTr_20_549,
    false,ptr_deref_551_data_0);
    ptr_deref_551_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_551_gather_scatter_ack_0 <= ptr_deref_551_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_20_549;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_551_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_551_root_address_inst_req_0,ptr_deref_551_root_address_inst_ack_0,sl_one,"ptr_deref_551_root_address_inst ",false,ptr_deref_551_resized_base_address,
    false,ptr_deref_551_root_address);
    ptr_deref_551_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_551_root_address_inst_ack_0 <= ptr_deref_551_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_551_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_551_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_556_addr_0_req_0,ptr_deref_556_addr_0_ack_0,sl_one,"ptr_deref_556_addr_0 ",false,ptr_deref_556_root_address,
    false,ptr_deref_556_word_address_0);
    ptr_deref_556_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_556_addr_0_ack_0 <= ptr_deref_556_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_556_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_556_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_556_base_resize_req_0,ptr_deref_556_base_resize_ack_0,sl_one,"ptr_deref_556_base_resize ",false,I_397,
    false,ptr_deref_556_resized_base_address);
    ptr_deref_556_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_556_base_resize_ack_0 <= ptr_deref_556_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_556_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_556_gather_scatter_req_0,ptr_deref_556_gather_scatter_ack_0,sl_one,"ptr_deref_556_gather_scatter ",false,ptr_deref_556_data_0,
    false,iNsTr_22_557);
    ptr_deref_556_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_556_gather_scatter_ack_0 <= ptr_deref_556_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_556_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_22_557 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_556_root_address_inst_req_0,ptr_deref_556_root_address_inst_ack_0,sl_one,"ptr_deref_556_root_address_inst ",false,ptr_deref_556_resized_base_address,
    false,ptr_deref_556_root_address);
    ptr_deref_556_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_556_root_address_inst_ack_0 <= ptr_deref_556_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_556_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_556_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_573_addr_0_req_0,ptr_deref_573_addr_0_ack_0,sl_one,"ptr_deref_573_addr_0 ",false,ptr_deref_573_root_address,
    false,ptr_deref_573_word_address_0);
    ptr_deref_573_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_573_addr_0_ack_0 <= ptr_deref_573_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_573_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_573_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_573_base_resize_req_0,ptr_deref_573_base_resize_ack_0,sl_one,"ptr_deref_573_base_resize ",false,I4_413,
    false,ptr_deref_573_resized_base_address);
    ptr_deref_573_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_573_base_resize_ack_0 <= ptr_deref_573_base_resize_req_0;
      in_aggregated_sig <= I4_413;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_573_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_573_gather_scatter_req_0,ptr_deref_573_gather_scatter_ack_0,sl_one,"ptr_deref_573_gather_scatter ",false,iNsTr_25_571,
    false,ptr_deref_573_data_0);
    ptr_deref_573_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_573_gather_scatter_ack_0 <= ptr_deref_573_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_25_571;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_573_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_573_root_address_inst_req_0,ptr_deref_573_root_address_inst_ack_0,sl_one,"ptr_deref_573_root_address_inst ",false,ptr_deref_573_resized_base_address,
    false,ptr_deref_573_root_address);
    ptr_deref_573_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_573_root_address_inst_ack_0 <= ptr_deref_573_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_573_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_573_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_578_addr_0_req_0,ptr_deref_578_addr_0_ack_0,sl_one,"ptr_deref_578_addr_0 ",false,ptr_deref_578_root_address,
    false,ptr_deref_578_word_address_0);
    ptr_deref_578_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_578_addr_0_ack_0 <= ptr_deref_578_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_578_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_578_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_578_base_resize_req_0,ptr_deref_578_base_resize_ack_0,sl_one,"ptr_deref_578_base_resize ",false,I_397,
    false,ptr_deref_578_resized_base_address);
    ptr_deref_578_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_578_base_resize_ack_0 <= ptr_deref_578_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_578_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_578_gather_scatter_req_0,ptr_deref_578_gather_scatter_ack_0,sl_one,"ptr_deref_578_gather_scatter ",false,ptr_deref_578_data_0,
    false,iNsTr_27_579);
    ptr_deref_578_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_578_gather_scatter_ack_0 <= ptr_deref_578_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_578_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_27_579 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_578_root_address_inst_req_0,ptr_deref_578_root_address_inst_ack_0,sl_one,"ptr_deref_578_root_address_inst ",false,ptr_deref_578_resized_base_address,
    false,ptr_deref_578_root_address);
    ptr_deref_578_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_578_root_address_inst_ack_0 <= ptr_deref_578_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_578_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_578_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_595_addr_0_req_0,ptr_deref_595_addr_0_ack_0,sl_one,"ptr_deref_595_addr_0 ",false,ptr_deref_595_root_address,
    false,ptr_deref_595_word_address_0);
    ptr_deref_595_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_595_addr_0_ack_0 <= ptr_deref_595_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_595_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_595_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_595_base_resize_req_0,ptr_deref_595_base_resize_ack_0,sl_one,"ptr_deref_595_base_resize ",false,I5_417,
    false,ptr_deref_595_resized_base_address);
    ptr_deref_595_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_595_base_resize_ack_0 <= ptr_deref_595_base_resize_req_0;
      in_aggregated_sig <= I5_417;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_595_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_595_gather_scatter_req_0,ptr_deref_595_gather_scatter_ack_0,sl_one,"ptr_deref_595_gather_scatter ",false,iNsTr_30_593,
    false,ptr_deref_595_data_0);
    ptr_deref_595_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_595_gather_scatter_ack_0 <= ptr_deref_595_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_30_593;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_595_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_595_root_address_inst_req_0,ptr_deref_595_root_address_inst_ack_0,sl_one,"ptr_deref_595_root_address_inst ",false,ptr_deref_595_resized_base_address,
    false,ptr_deref_595_root_address);
    ptr_deref_595_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_595_root_address_inst_ack_0 <= ptr_deref_595_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_595_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_595_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_600_addr_0_req_0,ptr_deref_600_addr_0_ack_0,sl_one,"ptr_deref_600_addr_0 ",false,ptr_deref_600_root_address,
    false,ptr_deref_600_word_address_0);
    ptr_deref_600_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_600_addr_0_ack_0 <= ptr_deref_600_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_600_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_600_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_600_base_resize_req_0,ptr_deref_600_base_resize_ack_0,sl_one,"ptr_deref_600_base_resize ",false,I_397,
    false,ptr_deref_600_resized_base_address);
    ptr_deref_600_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_600_base_resize_ack_0 <= ptr_deref_600_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_600_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_600_gather_scatter_req_0,ptr_deref_600_gather_scatter_ack_0,sl_one,"ptr_deref_600_gather_scatter ",false,ptr_deref_600_data_0,
    false,iNsTr_32_601);
    ptr_deref_600_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_600_gather_scatter_ack_0 <= ptr_deref_600_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_600_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_32_601 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_600_root_address_inst_req_0,ptr_deref_600_root_address_inst_ack_0,sl_one,"ptr_deref_600_root_address_inst ",false,ptr_deref_600_resized_base_address,
    false,ptr_deref_600_root_address);
    ptr_deref_600_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_600_root_address_inst_ack_0 <= ptr_deref_600_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_600_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_600_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_617_addr_0_req_0,ptr_deref_617_addr_0_ack_0,sl_one,"ptr_deref_617_addr_0 ",false,ptr_deref_617_root_address,
    false,ptr_deref_617_word_address_0);
    ptr_deref_617_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_617_addr_0_ack_0 <= ptr_deref_617_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_617_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_617_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_617_base_resize_req_0,ptr_deref_617_base_resize_ack_0,sl_one,"ptr_deref_617_base_resize ",false,I6_421,
    false,ptr_deref_617_resized_base_address);
    ptr_deref_617_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_617_base_resize_ack_0 <= ptr_deref_617_base_resize_req_0;
      in_aggregated_sig <= I6_421;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_617_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_617_gather_scatter_req_0,ptr_deref_617_gather_scatter_ack_0,sl_one,"ptr_deref_617_gather_scatter ",false,iNsTr_35_615,
    false,ptr_deref_617_data_0);
    ptr_deref_617_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_617_gather_scatter_ack_0 <= ptr_deref_617_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_35_615;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_617_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_617_root_address_inst_req_0,ptr_deref_617_root_address_inst_ack_0,sl_one,"ptr_deref_617_root_address_inst ",false,ptr_deref_617_resized_base_address,
    false,ptr_deref_617_root_address);
    ptr_deref_617_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_617_root_address_inst_ack_0 <= ptr_deref_617_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_617_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_617_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_622_addr_0_req_0,ptr_deref_622_addr_0_ack_0,sl_one,"ptr_deref_622_addr_0 ",false,ptr_deref_622_root_address,
    false,ptr_deref_622_word_address_0);
    ptr_deref_622_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_622_addr_0_ack_0 <= ptr_deref_622_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_622_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_622_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_622_base_resize_req_0,ptr_deref_622_base_resize_ack_0,sl_one,"ptr_deref_622_base_resize ",false,I_397,
    false,ptr_deref_622_resized_base_address);
    ptr_deref_622_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_622_base_resize_ack_0 <= ptr_deref_622_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_622_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_622_gather_scatter_req_0,ptr_deref_622_gather_scatter_ack_0,sl_one,"ptr_deref_622_gather_scatter ",false,ptr_deref_622_data_0,
    false,iNsTr_37_623);
    ptr_deref_622_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_622_gather_scatter_ack_0 <= ptr_deref_622_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_622_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_37_623 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_622_root_address_inst_req_0,ptr_deref_622_root_address_inst_ack_0,sl_one,"ptr_deref_622_root_address_inst ",false,ptr_deref_622_resized_base_address,
    false,ptr_deref_622_root_address);
    ptr_deref_622_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_622_root_address_inst_ack_0 <= ptr_deref_622_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_622_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_622_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_639_addr_0_req_0,ptr_deref_639_addr_0_ack_0,sl_one,"ptr_deref_639_addr_0 ",false,ptr_deref_639_root_address,
    false,ptr_deref_639_word_address_0);
    ptr_deref_639_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_639_addr_0_ack_0 <= ptr_deref_639_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_639_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_639_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_639_base_resize_req_0,ptr_deref_639_base_resize_ack_0,sl_one,"ptr_deref_639_base_resize ",false,I7_425,
    false,ptr_deref_639_resized_base_address);
    ptr_deref_639_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_639_base_resize_ack_0 <= ptr_deref_639_base_resize_req_0;
      in_aggregated_sig <= I7_425;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_639_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_639_gather_scatter_req_0,ptr_deref_639_gather_scatter_ack_0,sl_one,"ptr_deref_639_gather_scatter ",false,iNsTr_40_637,
    false,ptr_deref_639_data_0);
    ptr_deref_639_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_639_gather_scatter_ack_0 <= ptr_deref_639_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_40_637;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_639_data_0 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_639_root_address_inst_req_0,ptr_deref_639_root_address_inst_ack_0,sl_one,"ptr_deref_639_root_address_inst ",false,ptr_deref_639_resized_base_address,
    false,ptr_deref_639_root_address);
    ptr_deref_639_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_639_root_address_inst_ack_0 <= ptr_deref_639_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_639_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_639_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_644_addr_0_req_0,ptr_deref_644_addr_0_ack_0,sl_one,"ptr_deref_644_addr_0 ",false,ptr_deref_644_root_address,
    false,ptr_deref_644_word_address_0);
    ptr_deref_644_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_644_addr_0_ack_0 <= ptr_deref_644_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_644_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_644_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_644_base_resize_req_0,ptr_deref_644_base_resize_ack_0,sl_one,"ptr_deref_644_base_resize ",false,I_397,
    false,ptr_deref_644_resized_base_address);
    ptr_deref_644_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_644_base_resize_ack_0 <= ptr_deref_644_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_644_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_644_gather_scatter_req_0,ptr_deref_644_gather_scatter_ack_0,sl_one,"ptr_deref_644_gather_scatter ",false,ptr_deref_644_data_0,
    false,iNsTr_42_645);
    ptr_deref_644_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_644_gather_scatter_ack_0 <= ptr_deref_644_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_644_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_42_645 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_644_root_address_inst_req_0,ptr_deref_644_root_address_inst_ack_0,sl_one,"ptr_deref_644_root_address_inst ",false,ptr_deref_644_resized_base_address,
    false,ptr_deref_644_root_address);
    ptr_deref_644_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_644_root_address_inst_ack_0 <= ptr_deref_644_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_644_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_644_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_657_addr_0_req_0,ptr_deref_657_addr_0_ack_0,sl_one,"ptr_deref_657_addr_0 ",false,ptr_deref_657_root_address,
    false,ptr_deref_657_word_address_0);
    ptr_deref_657_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_657_addr_0_ack_0 <= ptr_deref_657_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_657_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_657_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_657_base_resize_req_0,ptr_deref_657_base_resize_ack_0,sl_one,"ptr_deref_657_base_resize ",false,iNsTr_44_654,
    false,ptr_deref_657_resized_base_address);
    ptr_deref_657_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_657_base_resize_ack_0 <= ptr_deref_657_base_resize_req_0;
      in_aggregated_sig <= iNsTr_44_654;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_657_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_657_gather_scatter_req_0,ptr_deref_657_gather_scatter_ack_0,sl_one,"ptr_deref_657_gather_scatter ",false,ptr_deref_657_data_0,
    false,iNsTr_45_658);
    ptr_deref_657_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_657_gather_scatter_ack_0 <= ptr_deref_657_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_657_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_45_658 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_657_root_address_inst_req_0,ptr_deref_657_root_address_inst_ack_0,sl_one,"ptr_deref_657_root_address_inst ",false,ptr_deref_657_resized_base_address,
    false,ptr_deref_657_root_address);
    ptr_deref_657_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_657_root_address_inst_ack_0 <= ptr_deref_657_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_657_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_657_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_661_addr_0_req_0,ptr_deref_661_addr_0_ack_0,sl_one,"ptr_deref_661_addr_0 ",false,ptr_deref_661_root_address,
    false,ptr_deref_661_word_address_0);
    ptr_deref_661_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_661_addr_0_ack_0 <= ptr_deref_661_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_661_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_661_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_661_base_resize_req_0,ptr_deref_661_base_resize_ack_0,sl_one,"ptr_deref_661_base_resize ",false,I_397,
    false,ptr_deref_661_resized_base_address);
    ptr_deref_661_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_661_base_resize_ack_0 <= ptr_deref_661_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_661_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_661_gather_scatter_req_0,ptr_deref_661_gather_scatter_ack_0,sl_one,"ptr_deref_661_gather_scatter ",false,ptr_deref_661_data_0,
    false,iNsTr_46_662);
    ptr_deref_661_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_661_gather_scatter_ack_0 <= ptr_deref_661_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_661_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_46_662 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_661_root_address_inst_req_0,ptr_deref_661_root_address_inst_ack_0,sl_one,"ptr_deref_661_root_address_inst ",false,ptr_deref_661_resized_base_address,
    false,ptr_deref_661_root_address);
    ptr_deref_661_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_661_root_address_inst_ack_0 <= ptr_deref_661_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_661_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_661_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_674_addr_0_req_0,ptr_deref_674_addr_0_ack_0,sl_one,"ptr_deref_674_addr_0 ",false,ptr_deref_674_root_address,
    false,ptr_deref_674_word_address_0);
    ptr_deref_674_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_674_addr_0_ack_0 <= ptr_deref_674_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_674_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_674_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_674_base_resize_req_0,ptr_deref_674_base_resize_ack_0,sl_one,"ptr_deref_674_base_resize ",false,iNsTr_48_671,
    false,ptr_deref_674_resized_base_address);
    ptr_deref_674_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_674_base_resize_ack_0 <= ptr_deref_674_base_resize_req_0;
      in_aggregated_sig <= iNsTr_48_671;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_674_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_674_gather_scatter_req_0,ptr_deref_674_gather_scatter_ack_0,sl_one,"ptr_deref_674_gather_scatter ",false,ptr_deref_674_data_0,
    false,iNsTr_49_675);
    ptr_deref_674_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_674_gather_scatter_ack_0 <= ptr_deref_674_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_674_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_49_675 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_674_root_address_inst_req_0,ptr_deref_674_root_address_inst_ack_0,sl_one,"ptr_deref_674_root_address_inst ",false,ptr_deref_674_resized_base_address,
    false,ptr_deref_674_root_address);
    ptr_deref_674_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_674_root_address_inst_ack_0 <= ptr_deref_674_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_674_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_674_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_682_addr_0_req_0,ptr_deref_682_addr_0_ack_0,sl_one,"ptr_deref_682_addr_0 ",false,ptr_deref_682_root_address,
    false,ptr_deref_682_word_address_0);
    ptr_deref_682_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_682_addr_0_ack_0 <= ptr_deref_682_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_682_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_682_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_682_base_resize_req_0,ptr_deref_682_base_resize_ack_0,sl_one,"ptr_deref_682_base_resize ",false,c0_429,
    false,ptr_deref_682_resized_base_address);
    ptr_deref_682_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_682_base_resize_ack_0 <= ptr_deref_682_base_resize_req_0;
      in_aggregated_sig <= c0_429;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_682_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_682_gather_scatter_req_0,ptr_deref_682_gather_scatter_ack_0,sl_one,"ptr_deref_682_gather_scatter ",false,iNsTr_50_680,
    false,ptr_deref_682_data_0);
    ptr_deref_682_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_682_gather_scatter_ack_0 <= ptr_deref_682_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_50_680;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_682_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_682_root_address_inst_req_0,ptr_deref_682_root_address_inst_ack_0,sl_one,"ptr_deref_682_root_address_inst ",false,ptr_deref_682_resized_base_address,
    false,ptr_deref_682_root_address);
    ptr_deref_682_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_682_root_address_inst_ack_0 <= ptr_deref_682_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_682_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_682_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_687_addr_0_req_0,ptr_deref_687_addr_0_ack_0,sl_one,"ptr_deref_687_addr_0 ",false,ptr_deref_687_root_address,
    false,ptr_deref_687_word_address_0);
    ptr_deref_687_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_687_addr_0_ack_0 <= ptr_deref_687_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_687_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_687_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_687_base_resize_req_0,ptr_deref_687_base_resize_ack_0,sl_one,"ptr_deref_687_base_resize ",false,I1_401,
    false,ptr_deref_687_resized_base_address);
    ptr_deref_687_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_687_base_resize_ack_0 <= ptr_deref_687_base_resize_req_0;
      in_aggregated_sig <= I1_401;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_687_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_687_gather_scatter_req_0,ptr_deref_687_gather_scatter_ack_0,sl_one,"ptr_deref_687_gather_scatter ",false,ptr_deref_687_data_0,
    false,iNsTr_52_688);
    ptr_deref_687_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_687_gather_scatter_ack_0 <= ptr_deref_687_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_687_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_52_688 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_687_root_address_inst_req_0,ptr_deref_687_root_address_inst_ack_0,sl_one,"ptr_deref_687_root_address_inst ",false,ptr_deref_687_resized_base_address,
    false,ptr_deref_687_root_address);
    ptr_deref_687_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_687_root_address_inst_ack_0 <= ptr_deref_687_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_687_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_687_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_700_addr_0_req_0,ptr_deref_700_addr_0_ack_0,sl_one,"ptr_deref_700_addr_0 ",false,ptr_deref_700_root_address,
    false,ptr_deref_700_word_address_0);
    ptr_deref_700_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_700_addr_0_ack_0 <= ptr_deref_700_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_700_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_700_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_700_base_resize_req_0,ptr_deref_700_base_resize_ack_0,sl_one,"ptr_deref_700_base_resize ",false,iNsTr_54_697,
    false,ptr_deref_700_resized_base_address);
    ptr_deref_700_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_700_base_resize_ack_0 <= ptr_deref_700_base_resize_req_0;
      in_aggregated_sig <= iNsTr_54_697;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_700_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_700_gather_scatter_req_0,ptr_deref_700_gather_scatter_ack_0,sl_one,"ptr_deref_700_gather_scatter ",false,ptr_deref_700_data_0,
    false,iNsTr_55_701);
    ptr_deref_700_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_700_gather_scatter_ack_0 <= ptr_deref_700_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_700_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_55_701 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_700_root_address_inst_req_0,ptr_deref_700_root_address_inst_ack_0,sl_one,"ptr_deref_700_root_address_inst ",false,ptr_deref_700_resized_base_address,
    false,ptr_deref_700_root_address);
    ptr_deref_700_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_700_root_address_inst_ack_0 <= ptr_deref_700_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_700_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_700_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_704_addr_0_req_0,ptr_deref_704_addr_0_ack_0,sl_one,"ptr_deref_704_addr_0 ",false,ptr_deref_704_root_address,
    false,ptr_deref_704_word_address_0);
    ptr_deref_704_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_704_addr_0_ack_0 <= ptr_deref_704_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_704_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_704_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_704_base_resize_req_0,ptr_deref_704_base_resize_ack_0,sl_one,"ptr_deref_704_base_resize ",false,I1_401,
    false,ptr_deref_704_resized_base_address);
    ptr_deref_704_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_704_base_resize_ack_0 <= ptr_deref_704_base_resize_req_0;
      in_aggregated_sig <= I1_401;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_704_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_704_gather_scatter_req_0,ptr_deref_704_gather_scatter_ack_0,sl_one,"ptr_deref_704_gather_scatter ",false,ptr_deref_704_data_0,
    false,iNsTr_56_705);
    ptr_deref_704_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_704_gather_scatter_ack_0 <= ptr_deref_704_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_704_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_56_705 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_704_root_address_inst_req_0,ptr_deref_704_root_address_inst_ack_0,sl_one,"ptr_deref_704_root_address_inst ",false,ptr_deref_704_resized_base_address,
    false,ptr_deref_704_root_address);
    ptr_deref_704_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_704_root_address_inst_ack_0 <= ptr_deref_704_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_704_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_704_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_717_addr_0_req_0,ptr_deref_717_addr_0_ack_0,sl_one,"ptr_deref_717_addr_0 ",false,ptr_deref_717_root_address,
    false,ptr_deref_717_word_address_0);
    ptr_deref_717_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_717_addr_0_ack_0 <= ptr_deref_717_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_717_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_717_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_717_base_resize_req_0,ptr_deref_717_base_resize_ack_0,sl_one,"ptr_deref_717_base_resize ",false,iNsTr_58_714,
    false,ptr_deref_717_resized_base_address);
    ptr_deref_717_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_717_base_resize_ack_0 <= ptr_deref_717_base_resize_req_0;
      in_aggregated_sig <= iNsTr_58_714;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_717_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_717_gather_scatter_req_0,ptr_deref_717_gather_scatter_ack_0,sl_one,"ptr_deref_717_gather_scatter ",false,ptr_deref_717_data_0,
    false,iNsTr_59_718);
    ptr_deref_717_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_717_gather_scatter_ack_0 <= ptr_deref_717_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_717_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_59_718 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_717_root_address_inst_req_0,ptr_deref_717_root_address_inst_ack_0,sl_one,"ptr_deref_717_root_address_inst ",false,ptr_deref_717_resized_base_address,
    false,ptr_deref_717_root_address);
    ptr_deref_717_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_717_root_address_inst_ack_0 <= ptr_deref_717_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_717_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_717_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_725_addr_0_req_0,ptr_deref_725_addr_0_ack_0,sl_one,"ptr_deref_725_addr_0 ",false,ptr_deref_725_root_address,
    false,ptr_deref_725_word_address_0);
    ptr_deref_725_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_725_addr_0_ack_0 <= ptr_deref_725_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_725_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_725_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_725_base_resize_req_0,ptr_deref_725_base_resize_ack_0,sl_one,"ptr_deref_725_base_resize ",false,c1_433,
    false,ptr_deref_725_resized_base_address);
    ptr_deref_725_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_725_base_resize_ack_0 <= ptr_deref_725_base_resize_req_0;
      in_aggregated_sig <= c1_433;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_725_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_725_gather_scatter_req_0,ptr_deref_725_gather_scatter_ack_0,sl_one,"ptr_deref_725_gather_scatter ",false,iNsTr_60_723,
    false,ptr_deref_725_data_0);
    ptr_deref_725_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_725_gather_scatter_ack_0 <= ptr_deref_725_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_60_723;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_725_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_725_root_address_inst_req_0,ptr_deref_725_root_address_inst_ack_0,sl_one,"ptr_deref_725_root_address_inst ",false,ptr_deref_725_resized_base_address,
    false,ptr_deref_725_root_address);
    ptr_deref_725_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_725_root_address_inst_ack_0 <= ptr_deref_725_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_725_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_725_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_730_addr_0_req_0,ptr_deref_730_addr_0_ack_0,sl_one,"ptr_deref_730_addr_0 ",false,ptr_deref_730_root_address,
    false,ptr_deref_730_word_address_0);
    ptr_deref_730_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_730_addr_0_ack_0 <= ptr_deref_730_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_730_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_730_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_730_base_resize_req_0,ptr_deref_730_base_resize_ack_0,sl_one,"ptr_deref_730_base_resize ",false,I2_405,
    false,ptr_deref_730_resized_base_address);
    ptr_deref_730_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_730_base_resize_ack_0 <= ptr_deref_730_base_resize_req_0;
      in_aggregated_sig <= I2_405;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_730_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_730_gather_scatter_req_0,ptr_deref_730_gather_scatter_ack_0,sl_one,"ptr_deref_730_gather_scatter ",false,ptr_deref_730_data_0,
    false,iNsTr_62_731);
    ptr_deref_730_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_730_gather_scatter_ack_0 <= ptr_deref_730_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_730_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_62_731 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_730_root_address_inst_req_0,ptr_deref_730_root_address_inst_ack_0,sl_one,"ptr_deref_730_root_address_inst ",false,ptr_deref_730_resized_base_address,
    false,ptr_deref_730_root_address);
    ptr_deref_730_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_730_root_address_inst_ack_0 <= ptr_deref_730_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_730_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_730_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_743_addr_0_req_0,ptr_deref_743_addr_0_ack_0,sl_one,"ptr_deref_743_addr_0 ",false,ptr_deref_743_root_address,
    false,ptr_deref_743_word_address_0);
    ptr_deref_743_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_743_addr_0_ack_0 <= ptr_deref_743_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_743_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_743_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_743_base_resize_req_0,ptr_deref_743_base_resize_ack_0,sl_one,"ptr_deref_743_base_resize ",false,iNsTr_64_740,
    false,ptr_deref_743_resized_base_address);
    ptr_deref_743_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_743_base_resize_ack_0 <= ptr_deref_743_base_resize_req_0;
      in_aggregated_sig <= iNsTr_64_740;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_743_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_743_gather_scatter_req_0,ptr_deref_743_gather_scatter_ack_0,sl_one,"ptr_deref_743_gather_scatter ",false,ptr_deref_743_data_0,
    false,iNsTr_65_744);
    ptr_deref_743_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_743_gather_scatter_ack_0 <= ptr_deref_743_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_743_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_65_744 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_743_root_address_inst_req_0,ptr_deref_743_root_address_inst_ack_0,sl_one,"ptr_deref_743_root_address_inst ",false,ptr_deref_743_resized_base_address,
    false,ptr_deref_743_root_address);
    ptr_deref_743_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_743_root_address_inst_ack_0 <= ptr_deref_743_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_743_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_743_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_747_addr_0_req_0,ptr_deref_747_addr_0_ack_0,sl_one,"ptr_deref_747_addr_0 ",false,ptr_deref_747_root_address,
    false,ptr_deref_747_word_address_0);
    ptr_deref_747_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_747_addr_0_ack_0 <= ptr_deref_747_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_747_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_747_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_747_base_resize_req_0,ptr_deref_747_base_resize_ack_0,sl_one,"ptr_deref_747_base_resize ",false,I2_405,
    false,ptr_deref_747_resized_base_address);
    ptr_deref_747_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_747_base_resize_ack_0 <= ptr_deref_747_base_resize_req_0;
      in_aggregated_sig <= I2_405;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_747_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_747_gather_scatter_req_0,ptr_deref_747_gather_scatter_ack_0,sl_one,"ptr_deref_747_gather_scatter ",false,ptr_deref_747_data_0,
    false,iNsTr_66_748);
    ptr_deref_747_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_747_gather_scatter_ack_0 <= ptr_deref_747_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_747_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_66_748 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_747_root_address_inst_req_0,ptr_deref_747_root_address_inst_ack_0,sl_one,"ptr_deref_747_root_address_inst ",false,ptr_deref_747_resized_base_address,
    false,ptr_deref_747_root_address);
    ptr_deref_747_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_747_root_address_inst_ack_0 <= ptr_deref_747_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_747_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_747_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_760_addr_0_req_0,ptr_deref_760_addr_0_ack_0,sl_one,"ptr_deref_760_addr_0 ",false,ptr_deref_760_root_address,
    false,ptr_deref_760_word_address_0);
    ptr_deref_760_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_760_addr_0_ack_0 <= ptr_deref_760_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_760_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_760_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_760_base_resize_req_0,ptr_deref_760_base_resize_ack_0,sl_one,"ptr_deref_760_base_resize ",false,iNsTr_68_757,
    false,ptr_deref_760_resized_base_address);
    ptr_deref_760_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_760_base_resize_ack_0 <= ptr_deref_760_base_resize_req_0;
      in_aggregated_sig <= iNsTr_68_757;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_760_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_760_gather_scatter_req_0,ptr_deref_760_gather_scatter_ack_0,sl_one,"ptr_deref_760_gather_scatter ",false,ptr_deref_760_data_0,
    false,iNsTr_69_761);
    ptr_deref_760_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_760_gather_scatter_ack_0 <= ptr_deref_760_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_760_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_69_761 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_760_root_address_inst_req_0,ptr_deref_760_root_address_inst_ack_0,sl_one,"ptr_deref_760_root_address_inst ",false,ptr_deref_760_resized_base_address,
    false,ptr_deref_760_root_address);
    ptr_deref_760_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_760_root_address_inst_ack_0 <= ptr_deref_760_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_760_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_760_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_768_addr_0_req_0,ptr_deref_768_addr_0_ack_0,sl_one,"ptr_deref_768_addr_0 ",false,ptr_deref_768_root_address,
    false,ptr_deref_768_word_address_0);
    ptr_deref_768_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_768_addr_0_ack_0 <= ptr_deref_768_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_768_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_768_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_768_base_resize_req_0,ptr_deref_768_base_resize_ack_0,sl_one,"ptr_deref_768_base_resize ",false,c2_437,
    false,ptr_deref_768_resized_base_address);
    ptr_deref_768_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_768_base_resize_ack_0 <= ptr_deref_768_base_resize_req_0;
      in_aggregated_sig <= c2_437;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_768_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_768_gather_scatter_req_0,ptr_deref_768_gather_scatter_ack_0,sl_one,"ptr_deref_768_gather_scatter ",false,iNsTr_70_766,
    false,ptr_deref_768_data_0);
    ptr_deref_768_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_768_gather_scatter_ack_0 <= ptr_deref_768_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_70_766;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_768_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_768_root_address_inst_req_0,ptr_deref_768_root_address_inst_ack_0,sl_one,"ptr_deref_768_root_address_inst ",false,ptr_deref_768_resized_base_address,
    false,ptr_deref_768_root_address);
    ptr_deref_768_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_768_root_address_inst_ack_0 <= ptr_deref_768_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_768_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_768_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_773_addr_0_req_0,ptr_deref_773_addr_0_ack_0,sl_one,"ptr_deref_773_addr_0 ",false,ptr_deref_773_root_address,
    false,ptr_deref_773_word_address_0);
    ptr_deref_773_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_773_addr_0_ack_0 <= ptr_deref_773_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_773_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_773_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_773_base_resize_req_0,ptr_deref_773_base_resize_ack_0,sl_one,"ptr_deref_773_base_resize ",false,I3_409,
    false,ptr_deref_773_resized_base_address);
    ptr_deref_773_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_773_base_resize_ack_0 <= ptr_deref_773_base_resize_req_0;
      in_aggregated_sig <= I3_409;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_773_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_773_gather_scatter_req_0,ptr_deref_773_gather_scatter_ack_0,sl_one,"ptr_deref_773_gather_scatter ",false,ptr_deref_773_data_0,
    false,iNsTr_72_774);
    ptr_deref_773_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_773_gather_scatter_ack_0 <= ptr_deref_773_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_773_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_72_774 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_773_root_address_inst_req_0,ptr_deref_773_root_address_inst_ack_0,sl_one,"ptr_deref_773_root_address_inst ",false,ptr_deref_773_resized_base_address,
    false,ptr_deref_773_root_address);
    ptr_deref_773_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_773_root_address_inst_ack_0 <= ptr_deref_773_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_773_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_773_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_786_addr_0_req_0,ptr_deref_786_addr_0_ack_0,sl_one,"ptr_deref_786_addr_0 ",false,ptr_deref_786_root_address,
    false,ptr_deref_786_word_address_0);
    ptr_deref_786_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_786_addr_0_ack_0 <= ptr_deref_786_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_786_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_786_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_786_base_resize_req_0,ptr_deref_786_base_resize_ack_0,sl_one,"ptr_deref_786_base_resize ",false,iNsTr_74_783,
    false,ptr_deref_786_resized_base_address);
    ptr_deref_786_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_786_base_resize_ack_0 <= ptr_deref_786_base_resize_req_0;
      in_aggregated_sig <= iNsTr_74_783;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_786_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_786_gather_scatter_req_0,ptr_deref_786_gather_scatter_ack_0,sl_one,"ptr_deref_786_gather_scatter ",false,ptr_deref_786_data_0,
    false,iNsTr_75_787);
    ptr_deref_786_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_786_gather_scatter_ack_0 <= ptr_deref_786_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_786_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_75_787 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_786_root_address_inst_req_0,ptr_deref_786_root_address_inst_ack_0,sl_one,"ptr_deref_786_root_address_inst ",false,ptr_deref_786_resized_base_address,
    false,ptr_deref_786_root_address);
    ptr_deref_786_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_786_root_address_inst_ack_0 <= ptr_deref_786_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_786_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_786_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_790_addr_0_req_0,ptr_deref_790_addr_0_ack_0,sl_one,"ptr_deref_790_addr_0 ",false,ptr_deref_790_root_address,
    false,ptr_deref_790_word_address_0);
    ptr_deref_790_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_790_addr_0_ack_0 <= ptr_deref_790_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_790_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_790_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_790_base_resize_req_0,ptr_deref_790_base_resize_ack_0,sl_one,"ptr_deref_790_base_resize ",false,I3_409,
    false,ptr_deref_790_resized_base_address);
    ptr_deref_790_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_790_base_resize_ack_0 <= ptr_deref_790_base_resize_req_0;
      in_aggregated_sig <= I3_409;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_790_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_790_gather_scatter_req_0,ptr_deref_790_gather_scatter_ack_0,sl_one,"ptr_deref_790_gather_scatter ",false,ptr_deref_790_data_0,
    false,iNsTr_76_791);
    ptr_deref_790_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_790_gather_scatter_ack_0 <= ptr_deref_790_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_790_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_76_791 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_790_root_address_inst_req_0,ptr_deref_790_root_address_inst_ack_0,sl_one,"ptr_deref_790_root_address_inst ",false,ptr_deref_790_resized_base_address,
    false,ptr_deref_790_root_address);
    ptr_deref_790_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_790_root_address_inst_ack_0 <= ptr_deref_790_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_790_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_790_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_803_addr_0_req_0,ptr_deref_803_addr_0_ack_0,sl_one,"ptr_deref_803_addr_0 ",false,ptr_deref_803_root_address,
    false,ptr_deref_803_word_address_0);
    ptr_deref_803_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_803_addr_0_ack_0 <= ptr_deref_803_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_803_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_803_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_803_base_resize_req_0,ptr_deref_803_base_resize_ack_0,sl_one,"ptr_deref_803_base_resize ",false,iNsTr_78_800,
    false,ptr_deref_803_resized_base_address);
    ptr_deref_803_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_803_base_resize_ack_0 <= ptr_deref_803_base_resize_req_0;
      in_aggregated_sig <= iNsTr_78_800;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_803_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_803_gather_scatter_req_0,ptr_deref_803_gather_scatter_ack_0,sl_one,"ptr_deref_803_gather_scatter ",false,ptr_deref_803_data_0,
    false,iNsTr_79_804);
    ptr_deref_803_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_803_gather_scatter_ack_0 <= ptr_deref_803_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_803_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_79_804 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_803_root_address_inst_req_0,ptr_deref_803_root_address_inst_ack_0,sl_one,"ptr_deref_803_root_address_inst ",false,ptr_deref_803_resized_base_address,
    false,ptr_deref_803_root_address);
    ptr_deref_803_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_803_root_address_inst_ack_0 <= ptr_deref_803_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_803_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_803_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_811_addr_0_req_0,ptr_deref_811_addr_0_ack_0,sl_one,"ptr_deref_811_addr_0 ",false,ptr_deref_811_root_address,
    false,ptr_deref_811_word_address_0);
    ptr_deref_811_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_811_addr_0_ack_0 <= ptr_deref_811_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_811_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_811_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_811_base_resize_req_0,ptr_deref_811_base_resize_ack_0,sl_one,"ptr_deref_811_base_resize ",false,c3_441,
    false,ptr_deref_811_resized_base_address);
    ptr_deref_811_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_811_base_resize_ack_0 <= ptr_deref_811_base_resize_req_0;
      in_aggregated_sig <= c3_441;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_811_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_811_gather_scatter_req_0,ptr_deref_811_gather_scatter_ack_0,sl_one,"ptr_deref_811_gather_scatter ",false,iNsTr_80_809,
    false,ptr_deref_811_data_0);
    ptr_deref_811_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_811_gather_scatter_ack_0 <= ptr_deref_811_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_80_809;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_811_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_811_root_address_inst_req_0,ptr_deref_811_root_address_inst_ack_0,sl_one,"ptr_deref_811_root_address_inst ",false,ptr_deref_811_resized_base_address,
    false,ptr_deref_811_root_address);
    ptr_deref_811_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_811_root_address_inst_ack_0 <= ptr_deref_811_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_811_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_811_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_816_addr_0_req_0,ptr_deref_816_addr_0_ack_0,sl_one,"ptr_deref_816_addr_0 ",false,ptr_deref_816_root_address,
    false,ptr_deref_816_word_address_0);
    ptr_deref_816_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_816_addr_0_ack_0 <= ptr_deref_816_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_816_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_816_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_816_base_resize_req_0,ptr_deref_816_base_resize_ack_0,sl_one,"ptr_deref_816_base_resize ",false,I4_413,
    false,ptr_deref_816_resized_base_address);
    ptr_deref_816_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_816_base_resize_ack_0 <= ptr_deref_816_base_resize_req_0;
      in_aggregated_sig <= I4_413;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_816_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_816_gather_scatter_req_0,ptr_deref_816_gather_scatter_ack_0,sl_one,"ptr_deref_816_gather_scatter ",false,ptr_deref_816_data_0,
    false,iNsTr_82_817);
    ptr_deref_816_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_816_gather_scatter_ack_0 <= ptr_deref_816_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_816_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_82_817 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_816_root_address_inst_req_0,ptr_deref_816_root_address_inst_ack_0,sl_one,"ptr_deref_816_root_address_inst ",false,ptr_deref_816_resized_base_address,
    false,ptr_deref_816_root_address);
    ptr_deref_816_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_816_root_address_inst_ack_0 <= ptr_deref_816_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_816_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_816_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_829_addr_0_req_0,ptr_deref_829_addr_0_ack_0,sl_one,"ptr_deref_829_addr_0 ",false,ptr_deref_829_root_address,
    false,ptr_deref_829_word_address_0);
    ptr_deref_829_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_829_addr_0_ack_0 <= ptr_deref_829_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_829_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_829_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_829_base_resize_req_0,ptr_deref_829_base_resize_ack_0,sl_one,"ptr_deref_829_base_resize ",false,iNsTr_84_826,
    false,ptr_deref_829_resized_base_address);
    ptr_deref_829_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_829_base_resize_ack_0 <= ptr_deref_829_base_resize_req_0;
      in_aggregated_sig <= iNsTr_84_826;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_829_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_829_gather_scatter_req_0,ptr_deref_829_gather_scatter_ack_0,sl_one,"ptr_deref_829_gather_scatter ",false,ptr_deref_829_data_0,
    false,iNsTr_85_830);
    ptr_deref_829_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_829_gather_scatter_ack_0 <= ptr_deref_829_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_829_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_85_830 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_829_root_address_inst_req_0,ptr_deref_829_root_address_inst_ack_0,sl_one,"ptr_deref_829_root_address_inst ",false,ptr_deref_829_resized_base_address,
    false,ptr_deref_829_root_address);
    ptr_deref_829_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_829_root_address_inst_ack_0 <= ptr_deref_829_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_829_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_829_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_833_addr_0_req_0,ptr_deref_833_addr_0_ack_0,sl_one,"ptr_deref_833_addr_0 ",false,ptr_deref_833_root_address,
    false,ptr_deref_833_word_address_0);
    ptr_deref_833_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_833_addr_0_ack_0 <= ptr_deref_833_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_833_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_833_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_833_base_resize_req_0,ptr_deref_833_base_resize_ack_0,sl_one,"ptr_deref_833_base_resize ",false,I4_413,
    false,ptr_deref_833_resized_base_address);
    ptr_deref_833_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_833_base_resize_ack_0 <= ptr_deref_833_base_resize_req_0;
      in_aggregated_sig <= I4_413;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_833_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_833_gather_scatter_req_0,ptr_deref_833_gather_scatter_ack_0,sl_one,"ptr_deref_833_gather_scatter ",false,ptr_deref_833_data_0,
    false,iNsTr_86_834);
    ptr_deref_833_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_833_gather_scatter_ack_0 <= ptr_deref_833_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_833_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_86_834 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_833_root_address_inst_req_0,ptr_deref_833_root_address_inst_ack_0,sl_one,"ptr_deref_833_root_address_inst ",false,ptr_deref_833_resized_base_address,
    false,ptr_deref_833_root_address);
    ptr_deref_833_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_833_root_address_inst_ack_0 <= ptr_deref_833_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_833_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_833_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_846_addr_0_req_0,ptr_deref_846_addr_0_ack_0,sl_one,"ptr_deref_846_addr_0 ",false,ptr_deref_846_root_address,
    false,ptr_deref_846_word_address_0);
    ptr_deref_846_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_846_addr_0_ack_0 <= ptr_deref_846_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_846_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_846_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_846_base_resize_req_0,ptr_deref_846_base_resize_ack_0,sl_one,"ptr_deref_846_base_resize ",false,iNsTr_88_843,
    false,ptr_deref_846_resized_base_address);
    ptr_deref_846_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_846_base_resize_ack_0 <= ptr_deref_846_base_resize_req_0;
      in_aggregated_sig <= iNsTr_88_843;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_846_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_846_gather_scatter_req_0,ptr_deref_846_gather_scatter_ack_0,sl_one,"ptr_deref_846_gather_scatter ",false,ptr_deref_846_data_0,
    false,iNsTr_89_847);
    ptr_deref_846_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_846_gather_scatter_ack_0 <= ptr_deref_846_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_846_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_89_847 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_846_root_address_inst_req_0,ptr_deref_846_root_address_inst_ack_0,sl_one,"ptr_deref_846_root_address_inst ",false,ptr_deref_846_resized_base_address,
    false,ptr_deref_846_root_address);
    ptr_deref_846_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_846_root_address_inst_ack_0 <= ptr_deref_846_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_846_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_846_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_854_addr_0_req_0,ptr_deref_854_addr_0_ack_0,sl_one,"ptr_deref_854_addr_0 ",false,ptr_deref_854_root_address,
    false,ptr_deref_854_word_address_0);
    ptr_deref_854_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_854_addr_0_ack_0 <= ptr_deref_854_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_854_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_854_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_854_base_resize_req_0,ptr_deref_854_base_resize_ack_0,sl_one,"ptr_deref_854_base_resize ",false,c4_445,
    false,ptr_deref_854_resized_base_address);
    ptr_deref_854_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_854_base_resize_ack_0 <= ptr_deref_854_base_resize_req_0;
      in_aggregated_sig <= c4_445;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_854_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_854_gather_scatter_req_0,ptr_deref_854_gather_scatter_ack_0,sl_one,"ptr_deref_854_gather_scatter ",false,iNsTr_90_852,
    false,ptr_deref_854_data_0);
    ptr_deref_854_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_854_gather_scatter_ack_0 <= ptr_deref_854_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_90_852;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_854_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_854_root_address_inst_req_0,ptr_deref_854_root_address_inst_ack_0,sl_one,"ptr_deref_854_root_address_inst ",false,ptr_deref_854_resized_base_address,
    false,ptr_deref_854_root_address);
    ptr_deref_854_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_854_root_address_inst_ack_0 <= ptr_deref_854_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_854_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_854_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_859_addr_0_req_0,ptr_deref_859_addr_0_ack_0,sl_one,"ptr_deref_859_addr_0 ",false,ptr_deref_859_root_address,
    false,ptr_deref_859_word_address_0);
    ptr_deref_859_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_859_addr_0_ack_0 <= ptr_deref_859_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_859_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_859_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_859_base_resize_req_0,ptr_deref_859_base_resize_ack_0,sl_one,"ptr_deref_859_base_resize ",false,I5_417,
    false,ptr_deref_859_resized_base_address);
    ptr_deref_859_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_859_base_resize_ack_0 <= ptr_deref_859_base_resize_req_0;
      in_aggregated_sig <= I5_417;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_859_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_859_gather_scatter_req_0,ptr_deref_859_gather_scatter_ack_0,sl_one,"ptr_deref_859_gather_scatter ",false,ptr_deref_859_data_0,
    false,iNsTr_92_860);
    ptr_deref_859_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_859_gather_scatter_ack_0 <= ptr_deref_859_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_859_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_92_860 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_859_root_address_inst_req_0,ptr_deref_859_root_address_inst_ack_0,sl_one,"ptr_deref_859_root_address_inst ",false,ptr_deref_859_resized_base_address,
    false,ptr_deref_859_root_address);
    ptr_deref_859_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_859_root_address_inst_ack_0 <= ptr_deref_859_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_859_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_859_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_872_addr_0_req_0,ptr_deref_872_addr_0_ack_0,sl_one,"ptr_deref_872_addr_0 ",false,ptr_deref_872_root_address,
    false,ptr_deref_872_word_address_0);
    ptr_deref_872_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_872_addr_0_ack_0 <= ptr_deref_872_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_872_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_872_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_872_base_resize_req_0,ptr_deref_872_base_resize_ack_0,sl_one,"ptr_deref_872_base_resize ",false,iNsTr_94_869,
    false,ptr_deref_872_resized_base_address);
    ptr_deref_872_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_872_base_resize_ack_0 <= ptr_deref_872_base_resize_req_0;
      in_aggregated_sig <= iNsTr_94_869;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_872_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_872_gather_scatter_req_0,ptr_deref_872_gather_scatter_ack_0,sl_one,"ptr_deref_872_gather_scatter ",false,ptr_deref_872_data_0,
    false,iNsTr_95_873);
    ptr_deref_872_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_872_gather_scatter_ack_0 <= ptr_deref_872_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_872_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_95_873 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_872_root_address_inst_req_0,ptr_deref_872_root_address_inst_ack_0,sl_one,"ptr_deref_872_root_address_inst ",false,ptr_deref_872_resized_base_address,
    false,ptr_deref_872_root_address);
    ptr_deref_872_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_872_root_address_inst_ack_0 <= ptr_deref_872_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_872_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_872_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_876_addr_0_req_0,ptr_deref_876_addr_0_ack_0,sl_one,"ptr_deref_876_addr_0 ",false,ptr_deref_876_root_address,
    false,ptr_deref_876_word_address_0);
    ptr_deref_876_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_876_addr_0_ack_0 <= ptr_deref_876_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_876_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_876_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_876_base_resize_req_0,ptr_deref_876_base_resize_ack_0,sl_one,"ptr_deref_876_base_resize ",false,I5_417,
    false,ptr_deref_876_resized_base_address);
    ptr_deref_876_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_876_base_resize_ack_0 <= ptr_deref_876_base_resize_req_0;
      in_aggregated_sig <= I5_417;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_876_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_876_gather_scatter_req_0,ptr_deref_876_gather_scatter_ack_0,sl_one,"ptr_deref_876_gather_scatter ",false,ptr_deref_876_data_0,
    false,iNsTr_96_877);
    ptr_deref_876_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_876_gather_scatter_ack_0 <= ptr_deref_876_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_876_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_96_877 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_876_root_address_inst_req_0,ptr_deref_876_root_address_inst_ack_0,sl_one,"ptr_deref_876_root_address_inst ",false,ptr_deref_876_resized_base_address,
    false,ptr_deref_876_root_address);
    ptr_deref_876_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_876_root_address_inst_ack_0 <= ptr_deref_876_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_876_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_876_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_889_addr_0_req_0,ptr_deref_889_addr_0_ack_0,sl_one,"ptr_deref_889_addr_0 ",false,ptr_deref_889_root_address,
    false,ptr_deref_889_word_address_0);
    ptr_deref_889_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_889_addr_0_ack_0 <= ptr_deref_889_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_889_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_889_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_889_base_resize_req_0,ptr_deref_889_base_resize_ack_0,sl_one,"ptr_deref_889_base_resize ",false,iNsTr_98_886,
    false,ptr_deref_889_resized_base_address);
    ptr_deref_889_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_889_base_resize_ack_0 <= ptr_deref_889_base_resize_req_0;
      in_aggregated_sig <= iNsTr_98_886;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_889_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_889_gather_scatter_req_0,ptr_deref_889_gather_scatter_ack_0,sl_one,"ptr_deref_889_gather_scatter ",false,ptr_deref_889_data_0,
    false,iNsTr_99_890);
    ptr_deref_889_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_889_gather_scatter_ack_0 <= ptr_deref_889_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_889_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_99_890 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_889_root_address_inst_req_0,ptr_deref_889_root_address_inst_ack_0,sl_one,"ptr_deref_889_root_address_inst ",false,ptr_deref_889_resized_base_address,
    false,ptr_deref_889_root_address);
    ptr_deref_889_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_889_root_address_inst_ack_0 <= ptr_deref_889_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_889_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_889_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_897_addr_0_req_0,ptr_deref_897_addr_0_ack_0,sl_one,"ptr_deref_897_addr_0 ",false,ptr_deref_897_root_address,
    false,ptr_deref_897_word_address_0);
    ptr_deref_897_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_897_addr_0_ack_0 <= ptr_deref_897_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_897_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_897_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_897_base_resize_req_0,ptr_deref_897_base_resize_ack_0,sl_one,"ptr_deref_897_base_resize ",false,c5_449,
    false,ptr_deref_897_resized_base_address);
    ptr_deref_897_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_897_base_resize_ack_0 <= ptr_deref_897_base_resize_req_0;
      in_aggregated_sig <= c5_449;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_897_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_897_gather_scatter_req_0,ptr_deref_897_gather_scatter_ack_0,sl_one,"ptr_deref_897_gather_scatter ",false,iNsTr_100_895,
    false,ptr_deref_897_data_0);
    ptr_deref_897_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_897_gather_scatter_ack_0 <= ptr_deref_897_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_100_895;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_897_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_897_root_address_inst_req_0,ptr_deref_897_root_address_inst_ack_0,sl_one,"ptr_deref_897_root_address_inst ",false,ptr_deref_897_resized_base_address,
    false,ptr_deref_897_root_address);
    ptr_deref_897_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_897_root_address_inst_ack_0 <= ptr_deref_897_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_897_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_897_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_902_addr_0_req_0,ptr_deref_902_addr_0_ack_0,sl_one,"ptr_deref_902_addr_0 ",false,ptr_deref_902_root_address,
    false,ptr_deref_902_word_address_0);
    ptr_deref_902_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_902_addr_0_ack_0 <= ptr_deref_902_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_902_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_902_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_902_base_resize_req_0,ptr_deref_902_base_resize_ack_0,sl_one,"ptr_deref_902_base_resize ",false,I6_421,
    false,ptr_deref_902_resized_base_address);
    ptr_deref_902_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_902_base_resize_ack_0 <= ptr_deref_902_base_resize_req_0;
      in_aggregated_sig <= I6_421;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_902_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_902_gather_scatter_req_0,ptr_deref_902_gather_scatter_ack_0,sl_one,"ptr_deref_902_gather_scatter ",false,ptr_deref_902_data_0,
    false,iNsTr_102_903);
    ptr_deref_902_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_902_gather_scatter_ack_0 <= ptr_deref_902_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_902_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_102_903 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_902_root_address_inst_req_0,ptr_deref_902_root_address_inst_ack_0,sl_one,"ptr_deref_902_root_address_inst ",false,ptr_deref_902_resized_base_address,
    false,ptr_deref_902_root_address);
    ptr_deref_902_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_902_root_address_inst_ack_0 <= ptr_deref_902_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_902_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_902_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_915_addr_0_req_0,ptr_deref_915_addr_0_ack_0,sl_one,"ptr_deref_915_addr_0 ",false,ptr_deref_915_root_address,
    false,ptr_deref_915_word_address_0);
    ptr_deref_915_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_915_addr_0_ack_0 <= ptr_deref_915_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_915_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_915_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_915_base_resize_req_0,ptr_deref_915_base_resize_ack_0,sl_one,"ptr_deref_915_base_resize ",false,iNsTr_104_912,
    false,ptr_deref_915_resized_base_address);
    ptr_deref_915_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_915_base_resize_ack_0 <= ptr_deref_915_base_resize_req_0;
      in_aggregated_sig <= iNsTr_104_912;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_915_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_915_gather_scatter_req_0,ptr_deref_915_gather_scatter_ack_0,sl_one,"ptr_deref_915_gather_scatter ",false,ptr_deref_915_data_0,
    false,iNsTr_105_916);
    ptr_deref_915_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_915_gather_scatter_ack_0 <= ptr_deref_915_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_915_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_105_916 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_915_root_address_inst_req_0,ptr_deref_915_root_address_inst_ack_0,sl_one,"ptr_deref_915_root_address_inst ",false,ptr_deref_915_resized_base_address,
    false,ptr_deref_915_root_address);
    ptr_deref_915_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_915_root_address_inst_ack_0 <= ptr_deref_915_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_915_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_915_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_919_addr_0_req_0,ptr_deref_919_addr_0_ack_0,sl_one,"ptr_deref_919_addr_0 ",false,ptr_deref_919_root_address,
    false,ptr_deref_919_word_address_0);
    ptr_deref_919_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_919_addr_0_ack_0 <= ptr_deref_919_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_919_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_919_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_919_base_resize_req_0,ptr_deref_919_base_resize_ack_0,sl_one,"ptr_deref_919_base_resize ",false,I6_421,
    false,ptr_deref_919_resized_base_address);
    ptr_deref_919_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_919_base_resize_ack_0 <= ptr_deref_919_base_resize_req_0;
      in_aggregated_sig <= I6_421;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_919_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_919_gather_scatter_req_0,ptr_deref_919_gather_scatter_ack_0,sl_one,"ptr_deref_919_gather_scatter ",false,ptr_deref_919_data_0,
    false,iNsTr_106_920);
    ptr_deref_919_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_919_gather_scatter_ack_0 <= ptr_deref_919_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_919_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_106_920 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_919_root_address_inst_req_0,ptr_deref_919_root_address_inst_ack_0,sl_one,"ptr_deref_919_root_address_inst ",false,ptr_deref_919_resized_base_address,
    false,ptr_deref_919_root_address);
    ptr_deref_919_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_919_root_address_inst_ack_0 <= ptr_deref_919_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_919_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_919_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_932_addr_0_req_0,ptr_deref_932_addr_0_ack_0,sl_one,"ptr_deref_932_addr_0 ",false,ptr_deref_932_root_address,
    false,ptr_deref_932_word_address_0);
    ptr_deref_932_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_932_addr_0_ack_0 <= ptr_deref_932_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_932_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_932_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_932_base_resize_req_0,ptr_deref_932_base_resize_ack_0,sl_one,"ptr_deref_932_base_resize ",false,iNsTr_108_929,
    false,ptr_deref_932_resized_base_address);
    ptr_deref_932_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_932_base_resize_ack_0 <= ptr_deref_932_base_resize_req_0;
      in_aggregated_sig <= iNsTr_108_929;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_932_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_932_gather_scatter_req_0,ptr_deref_932_gather_scatter_ack_0,sl_one,"ptr_deref_932_gather_scatter ",false,ptr_deref_932_data_0,
    false,iNsTr_109_933);
    ptr_deref_932_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_932_gather_scatter_ack_0 <= ptr_deref_932_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_932_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_109_933 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_932_root_address_inst_req_0,ptr_deref_932_root_address_inst_ack_0,sl_one,"ptr_deref_932_root_address_inst ",false,ptr_deref_932_resized_base_address,
    false,ptr_deref_932_root_address);
    ptr_deref_932_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_932_root_address_inst_ack_0 <= ptr_deref_932_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_932_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_932_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_940_addr_0_req_0,ptr_deref_940_addr_0_ack_0,sl_one,"ptr_deref_940_addr_0 ",false,ptr_deref_940_root_address,
    false,ptr_deref_940_word_address_0);
    ptr_deref_940_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_940_addr_0_ack_0 <= ptr_deref_940_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_940_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_940_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_940_base_resize_req_0,ptr_deref_940_base_resize_ack_0,sl_one,"ptr_deref_940_base_resize ",false,c6_453,
    false,ptr_deref_940_resized_base_address);
    ptr_deref_940_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_940_base_resize_ack_0 <= ptr_deref_940_base_resize_req_0;
      in_aggregated_sig <= c6_453;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_940_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_940_gather_scatter_req_0,ptr_deref_940_gather_scatter_ack_0,sl_one,"ptr_deref_940_gather_scatter ",false,iNsTr_110_938,
    false,ptr_deref_940_data_0);
    ptr_deref_940_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_940_gather_scatter_ack_0 <= ptr_deref_940_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_110_938;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_940_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_940_root_address_inst_req_0,ptr_deref_940_root_address_inst_ack_0,sl_one,"ptr_deref_940_root_address_inst ",false,ptr_deref_940_resized_base_address,
    false,ptr_deref_940_root_address);
    ptr_deref_940_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_940_root_address_inst_ack_0 <= ptr_deref_940_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_940_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_940_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_945_addr_0_req_0,ptr_deref_945_addr_0_ack_0,sl_one,"ptr_deref_945_addr_0 ",false,ptr_deref_945_root_address,
    false,ptr_deref_945_word_address_0);
    ptr_deref_945_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_945_addr_0_ack_0 <= ptr_deref_945_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_945_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_945_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_945_base_resize_req_0,ptr_deref_945_base_resize_ack_0,sl_one,"ptr_deref_945_base_resize ",false,I7_425,
    false,ptr_deref_945_resized_base_address);
    ptr_deref_945_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_945_base_resize_ack_0 <= ptr_deref_945_base_resize_req_0;
      in_aggregated_sig <= I7_425;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_945_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_945_gather_scatter_req_0,ptr_deref_945_gather_scatter_ack_0,sl_one,"ptr_deref_945_gather_scatter ",false,ptr_deref_945_data_0,
    false,iNsTr_112_946);
    ptr_deref_945_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_945_gather_scatter_ack_0 <= ptr_deref_945_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_945_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_112_946 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_945_root_address_inst_req_0,ptr_deref_945_root_address_inst_ack_0,sl_one,"ptr_deref_945_root_address_inst ",false,ptr_deref_945_resized_base_address,
    false,ptr_deref_945_root_address);
    ptr_deref_945_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_945_root_address_inst_ack_0 <= ptr_deref_945_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_945_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_945_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_958_addr_0_req_0,ptr_deref_958_addr_0_ack_0,sl_one,"ptr_deref_958_addr_0 ",false,ptr_deref_958_root_address,
    false,ptr_deref_958_word_address_0);
    ptr_deref_958_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_958_addr_0_ack_0 <= ptr_deref_958_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_958_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_958_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_958_base_resize_req_0,ptr_deref_958_base_resize_ack_0,sl_one,"ptr_deref_958_base_resize ",false,iNsTr_114_955,
    false,ptr_deref_958_resized_base_address);
    ptr_deref_958_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_958_base_resize_ack_0 <= ptr_deref_958_base_resize_req_0;
      in_aggregated_sig <= iNsTr_114_955;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_958_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_958_gather_scatter_req_0,ptr_deref_958_gather_scatter_ack_0,sl_one,"ptr_deref_958_gather_scatter ",false,ptr_deref_958_data_0,
    false,iNsTr_115_959);
    ptr_deref_958_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_958_gather_scatter_ack_0 <= ptr_deref_958_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_958_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_115_959 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_958_root_address_inst_req_0,ptr_deref_958_root_address_inst_ack_0,sl_one,"ptr_deref_958_root_address_inst ",false,ptr_deref_958_resized_base_address,
    false,ptr_deref_958_root_address);
    ptr_deref_958_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_958_root_address_inst_ack_0 <= ptr_deref_958_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_958_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_958_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_962_addr_0_req_0,ptr_deref_962_addr_0_ack_0,sl_one,"ptr_deref_962_addr_0 ",false,ptr_deref_962_root_address,
    false,ptr_deref_962_word_address_0);
    ptr_deref_962_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_962_addr_0_ack_0 <= ptr_deref_962_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_962_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_962_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_962_base_resize_req_0,ptr_deref_962_base_resize_ack_0,sl_one,"ptr_deref_962_base_resize ",false,I7_425,
    false,ptr_deref_962_resized_base_address);
    ptr_deref_962_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_962_base_resize_ack_0 <= ptr_deref_962_base_resize_req_0;
      in_aggregated_sig <= I7_425;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_962_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_962_gather_scatter_req_0,ptr_deref_962_gather_scatter_ack_0,sl_one,"ptr_deref_962_gather_scatter ",false,ptr_deref_962_data_0,
    false,iNsTr_116_963);
    ptr_deref_962_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_962_gather_scatter_ack_0 <= ptr_deref_962_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_962_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_116_963 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_962_root_address_inst_req_0,ptr_deref_962_root_address_inst_ack_0,sl_one,"ptr_deref_962_root_address_inst ",false,ptr_deref_962_resized_base_address,
    false,ptr_deref_962_root_address);
    ptr_deref_962_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_962_root_address_inst_ack_0 <= ptr_deref_962_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_962_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_962_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_975_addr_0_req_0,ptr_deref_975_addr_0_ack_0,sl_one,"ptr_deref_975_addr_0 ",false,ptr_deref_975_root_address,
    false,ptr_deref_975_word_address_0);
    ptr_deref_975_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_975_addr_0_ack_0 <= ptr_deref_975_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_975_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_975_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_975_base_resize_req_0,ptr_deref_975_base_resize_ack_0,sl_one,"ptr_deref_975_base_resize ",false,iNsTr_118_972,
    false,ptr_deref_975_resized_base_address);
    ptr_deref_975_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_975_base_resize_ack_0 <= ptr_deref_975_base_resize_req_0;
      in_aggregated_sig <= iNsTr_118_972;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_975_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_975_gather_scatter_req_0,ptr_deref_975_gather_scatter_ack_0,sl_one,"ptr_deref_975_gather_scatter ",false,ptr_deref_975_data_0,
    false,iNsTr_119_976);
    ptr_deref_975_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_975_gather_scatter_ack_0 <= ptr_deref_975_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_975_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_119_976 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_975_root_address_inst_req_0,ptr_deref_975_root_address_inst_ack_0,sl_one,"ptr_deref_975_root_address_inst ",false,ptr_deref_975_resized_base_address,
    false,ptr_deref_975_root_address);
    ptr_deref_975_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_975_root_address_inst_ack_0 <= ptr_deref_975_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_975_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_975_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_983_addr_0_req_0,ptr_deref_983_addr_0_ack_0,sl_one,"ptr_deref_983_addr_0 ",false,ptr_deref_983_root_address,
    false,ptr_deref_983_word_address_0);
    ptr_deref_983_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_983_addr_0_ack_0 <= ptr_deref_983_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_983_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_983_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_983_base_resize_req_0,ptr_deref_983_base_resize_ack_0,sl_one,"ptr_deref_983_base_resize ",false,c7_457,
    false,ptr_deref_983_resized_base_address);
    ptr_deref_983_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_983_base_resize_ack_0 <= ptr_deref_983_base_resize_req_0;
      in_aggregated_sig <= c7_457;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_983_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_983_gather_scatter_req_0,ptr_deref_983_gather_scatter_ack_0,sl_one,"ptr_deref_983_gather_scatter ",false,iNsTr_120_981,
    false,ptr_deref_983_data_0);
    ptr_deref_983_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_983_gather_scatter_ack_0 <= ptr_deref_983_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_120_981;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_983_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_983_root_address_inst_req_0,ptr_deref_983_root_address_inst_ack_0,sl_one,"ptr_deref_983_root_address_inst ",false,ptr_deref_983_resized_base_address,
    false,ptr_deref_983_root_address);
    ptr_deref_983_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_983_root_address_inst_ack_0 <= ptr_deref_983_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_983_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_983_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_988_addr_0_req_0,ptr_deref_988_addr_0_ack_0,sl_one,"ptr_deref_988_addr_0 ",false,ptr_deref_988_root_address,
    false,ptr_deref_988_word_address_0);
    ptr_deref_988_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_988_addr_0_ack_0 <= ptr_deref_988_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_988_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_988_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_988_base_resize_req_0,ptr_deref_988_base_resize_ack_0,sl_one,"ptr_deref_988_base_resize ",false,c0_429,
    false,ptr_deref_988_resized_base_address);
    ptr_deref_988_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_988_base_resize_ack_0 <= ptr_deref_988_base_resize_req_0;
      in_aggregated_sig <= c0_429;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_988_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_988_gather_scatter_req_0,ptr_deref_988_gather_scatter_ack_0,sl_one,"ptr_deref_988_gather_scatter ",false,ptr_deref_988_data_0,
    false,iNsTr_122_989);
    ptr_deref_988_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_988_gather_scatter_ack_0 <= ptr_deref_988_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_988_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_122_989 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_988_root_address_inst_req_0,ptr_deref_988_root_address_inst_ack_0,sl_one,"ptr_deref_988_root_address_inst ",false,ptr_deref_988_resized_base_address,
    false,ptr_deref_988_root_address);
    ptr_deref_988_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_988_root_address_inst_ack_0 <= ptr_deref_988_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_988_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_988_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_992_addr_0_req_0,ptr_deref_992_addr_0_ack_0,sl_one,"ptr_deref_992_addr_0 ",false,ptr_deref_992_root_address,
    false,ptr_deref_992_word_address_0);
    ptr_deref_992_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_992_addr_0_ack_0 <= ptr_deref_992_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_992_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_992_word_address_0 <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_992_base_resize_req_0,ptr_deref_992_base_resize_ack_0,sl_one,"ptr_deref_992_base_resize ",false,I_397,
    false,ptr_deref_992_resized_base_address);
    ptr_deref_992_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_992_base_resize_ack_0 <= ptr_deref_992_base_resize_req_0;
      in_aggregated_sig <= I_397;
      out_aggregated_sig <= in_aggregated_sig(0 downto 0);
      ptr_deref_992_resized_base_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_992_gather_scatter_req_0,ptr_deref_992_gather_scatter_ack_0,sl_one,"ptr_deref_992_gather_scatter ",false,ptr_deref_992_data_0,
    false,iNsTr_123_993);
    ptr_deref_992_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(7 downto 0);
      signal out_aggregated_sig: std_logic_vector(7 downto 0);
      --
    begin -- 
      ptr_deref_992_gather_scatter_ack_0 <= ptr_deref_992_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_992_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_123_993 <= out_aggregated_sig(7 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_992_root_address_inst_req_0,ptr_deref_992_root_address_inst_ack_0,sl_one,"ptr_deref_992_root_address_inst ",false,ptr_deref_992_resized_base_address,
    false,ptr_deref_992_root_address);
    ptr_deref_992_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(0 downto 0);
      signal out_aggregated_sig: std_logic_vector(0 downto 0);
      --
    begin -- 
      ptr_deref_992_root_address_inst_ack_0 <= ptr_deref_992_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_992_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_992_root_address <= out_aggregated_sig(0 downto 0);
      --
    end Block;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_481_branch_req_0," req0 if_stmt_481_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_481_branch_ack_0," ack0 if_stmt_481_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_481_branch_ack_1," ack1 if_stmt_481_branch");
    if_stmt_481_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_4_480;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_481_branch_req_0,
          ack0 => if_stmt_481_branch_ack_0,
          ack1 => if_stmt_481_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_1168_inst_req_0,binary_1168_inst_ack_0,binary_1168_inst_req_1,binary_1168_inst_ack_1,sl_one,"binary_1168_inst",false,iNsTr_165_1163 & type_cast_1167_wire_constant,
    false,iNsTr_166_1169);
    -- shared split operator group (0) : binary_1168_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_165_1163;
      iNsTr_166_1169 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_1168_inst_req_0;
      reqR(0) <= binary_1168_inst_req_1;
      binary_1168_inst_ack_0 <= ackL(0); 
      binary_1168_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_479_inst_req_0,binary_479_inst_ack_0,binary_479_inst_req_1,binary_479_inst_ack_1,sl_one,"binary_479_inst",false,type_cast_475_wire & type_cast_478_wire_constant,
    false,iNsTr_4_480);
    -- shared split operator group (1) : binary_479_inst 
    ApIntSlt_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_475_wire;
      iNsTr_4_480 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_479_inst_req_0;
      reqR(0) <= binary_479_inst_req_1;
      binary_479_inst_ack_0 <= ackL(0); 
      binary_479_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_500_inst_req_0,binary_500_inst_ack_0,binary_500_inst_req_1,binary_500_inst_ack_1,sl_one,"binary_500_inst",false,iNsTr_8_495 & type_cast_499_wire_constant,
    false,iNsTr_9_501);
    -- shared split operator group (2) : binary_500_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_8_495;
      iNsTr_9_501 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_500_inst_req_0;
      reqR(0) <= binary_500_inst_req_1;
      binary_500_inst_ack_0 <= ackL(0); 
      binary_500_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_522_inst_req_0,binary_522_inst_ack_0,binary_522_inst_req_1,binary_522_inst_ack_1,sl_one,"binary_522_inst",false,iNsTr_13_517 & type_cast_521_wire_constant,
    false,iNsTr_14_523);
    -- shared split operator group (3) : binary_522_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_13_517;
      iNsTr_14_523 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_522_inst_req_0;
      reqR(0) <= binary_522_inst_req_1;
      binary_522_inst_ack_0 <= ackL(0); 
      binary_522_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_544_inst_req_0,binary_544_inst_ack_0,binary_544_inst_req_1,binary_544_inst_ack_1,sl_one,"binary_544_inst",false,iNsTr_18_539 & type_cast_543_wire_constant,
    false,iNsTr_19_545);
    -- shared split operator group (4) : binary_544_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_18_539;
      iNsTr_19_545 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_544_inst_req_0;
      reqR(0) <= binary_544_inst_req_1;
      binary_544_inst_ack_0 <= ackL(0); 
      binary_544_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_566_inst_req_0,binary_566_inst_ack_0,binary_566_inst_req_1,binary_566_inst_ack_1,sl_one,"binary_566_inst",false,iNsTr_23_561 & type_cast_565_wire_constant,
    false,iNsTr_24_567);
    -- shared split operator group (5) : binary_566_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_23_561;
      iNsTr_24_567 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_566_inst_req_0;
      reqR(0) <= binary_566_inst_req_1;
      binary_566_inst_ack_0 <= ackL(0); 
      binary_566_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_588_inst_req_0,binary_588_inst_ack_0,binary_588_inst_req_1,binary_588_inst_ack_1,sl_one,"binary_588_inst",false,iNsTr_28_583 & type_cast_587_wire_constant,
    false,iNsTr_29_589);
    -- shared split operator group (6) : binary_588_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_28_583;
      iNsTr_29_589 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_588_inst_req_0;
      reqR(0) <= binary_588_inst_req_1;
      binary_588_inst_ack_0 <= ackL(0); 
      binary_588_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_610_inst_req_0,binary_610_inst_ack_0,binary_610_inst_req_1,binary_610_inst_ack_1,sl_one,"binary_610_inst",false,iNsTr_33_605 & type_cast_609_wire_constant,
    false,iNsTr_34_611);
    -- shared split operator group (7) : binary_610_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_33_605;
      iNsTr_34_611 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_610_inst_req_0;
      reqR(0) <= binary_610_inst_req_1;
      binary_610_inst_ack_0 <= ackL(0); 
      binary_610_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_632_inst_req_0,binary_632_inst_ack_0,binary_632_inst_req_1,binary_632_inst_ack_1,sl_one,"binary_632_inst",false,iNsTr_38_627 & type_cast_631_wire_constant,
    false,iNsTr_39_633);
    -- shared split operator group (8) : binary_632_inst 
    ApIntAdd_group_8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_38_627;
      iNsTr_39_633 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_632_inst_req_0;
      reqR(0) <= binary_632_inst_req_1;
      binary_632_inst_ack_0 <= ackL(0); 
      binary_632_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_679_inst_req_0,binary_679_inst_ack_0,binary_679_inst_req_1,binary_679_inst_ack_1,sl_one,"binary_679_inst",false,iNsTr_45_658 & iNsTr_49_675,
    false,iNsTr_50_680);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_722_inst_req_0,binary_722_inst_ack_0,binary_722_inst_req_1,binary_722_inst_ack_1,sl_one,"binary_722_inst",false,iNsTr_55_701 & iNsTr_59_718,
    false,iNsTr_60_723);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_765_inst_req_0,binary_765_inst_ack_0,binary_765_inst_req_1,binary_765_inst_ack_1,sl_one,"binary_765_inst",false,iNsTr_65_744 & iNsTr_69_761,
    false,iNsTr_70_766);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_980_inst_req_0,binary_980_inst_ack_0,binary_980_inst_req_1,binary_980_inst_ack_1,sl_one,"binary_980_inst",false,iNsTr_115_959 & iNsTr_119_976,
    false,iNsTr_120_981);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_808_inst_req_0,binary_808_inst_ack_0,binary_808_inst_req_1,binary_808_inst_ack_1,sl_one,"binary_808_inst",false,iNsTr_75_787 & iNsTr_79_804,
    false,iNsTr_80_809);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_851_inst_req_0,binary_851_inst_ack_0,binary_851_inst_req_1,binary_851_inst_ack_1,sl_one,"binary_851_inst",false,iNsTr_85_830 & iNsTr_89_847,
    false,iNsTr_90_852);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_894_inst_req_0,binary_894_inst_ack_0,binary_894_inst_req_1,binary_894_inst_ack_1,sl_one,"binary_894_inst",false,iNsTr_95_873 & iNsTr_99_890,
    false,iNsTr_100_895);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_937_inst_req_0,binary_937_inst_ack_0,binary_937_inst_req_1,binary_937_inst_ack_1,sl_one,"binary_937_inst",false,iNsTr_105_916 & iNsTr_109_933,
    false,iNsTr_110_938);
    -- shared split operator group (9) : binary_679_inst binary_722_inst binary_765_inst binary_980_inst binary_808_inst binary_851_inst binary_894_inst binary_937_inst 
    ApFloatAdd_group_9: Block -- 
      signal data_in: std_logic_vector(511 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_45_658 & iNsTr_49_675 & iNsTr_55_701 & iNsTr_59_718 & iNsTr_65_744 & iNsTr_69_761 & iNsTr_115_959 & iNsTr_119_976 & iNsTr_75_787 & iNsTr_79_804 & iNsTr_85_830 & iNsTr_89_847 & iNsTr_95_873 & iNsTr_99_890 & iNsTr_105_916 & iNsTr_109_933;
      iNsTr_50_680 <= data_out(255 downto 224);
      iNsTr_60_723 <= data_out(223 downto 192);
      iNsTr_70_766 <= data_out(191 downto 160);
      iNsTr_120_981 <= data_out(159 downto 128);
      iNsTr_80_809 <= data_out(127 downto 96);
      iNsTr_90_852 <= data_out(95 downto 64);
      iNsTr_100_895 <= data_out(63 downto 32);
      iNsTr_110_938 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      reqL_unguarded(7) <= binary_679_inst_req_0;
      reqL_unguarded(6) <= binary_722_inst_req_0;
      reqL_unguarded(5) <= binary_765_inst_req_0;
      reqL_unguarded(4) <= binary_980_inst_req_0;
      reqL_unguarded(3) <= binary_808_inst_req_0;
      reqL_unguarded(2) <= binary_851_inst_req_0;
      reqL_unguarded(1) <= binary_894_inst_req_0;
      reqL_unguarded(0) <= binary_937_inst_req_0;
      binary_679_inst_ack_0 <= ackL_unguarded(7);
      binary_722_inst_ack_0 <= ackL_unguarded(6);
      binary_765_inst_ack_0 <= ackL_unguarded(5);
      binary_980_inst_ack_0 <= ackL_unguarded(4);
      binary_808_inst_ack_0 <= ackL_unguarded(3);
      binary_851_inst_ack_0 <= ackL_unguarded(2);
      binary_894_inst_ack_0 <= ackL_unguarded(1);
      binary_937_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= binary_679_inst_req_1;
      reqR_unguarded(6) <= binary_722_inst_req_1;
      reqR_unguarded(5) <= binary_765_inst_req_1;
      reqR_unguarded(4) <= binary_980_inst_req_1;
      reqR_unguarded(3) <= binary_808_inst_req_1;
      reqR_unguarded(2) <= binary_851_inst_req_1;
      reqR_unguarded(1) <= binary_894_inst_req_1;
      reqR_unguarded(0) <= binary_937_inst_req_1;
      binary_679_inst_ack_1 <= ackR_unguarded(7);
      binary_722_inst_ack_1 <= ackR_unguarded(6);
      binary_765_inst_ack_1 <= ackR_unguarded(5);
      binary_980_inst_ack_1 <= ackR_unguarded(4);
      binary_808_inst_ack_1 <= ackR_unguarded(3);
      binary_851_inst_ack_1 <= ackR_unguarded(2);
      binary_894_inst_ack_1 <= ackR_unguarded(1);
      binary_937_inst_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 8 -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1009_load_0_req_0,ptr_deref_1009_load_0_ack_0,ptr_deref_1009_load_0_req_1,ptr_deref_1009_load_0_ack_1,sl_one,"ptr_deref_1009_load_0",false,ptr_deref_1009_word_address_0,
    false,ptr_deref_1009_data_0);
    -- shared load operator group (0) : ptr_deref_1009_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1009_load_0_req_0,
        ptr_deref_1009_load_0_ack_0,
        ptr_deref_1009_load_0_req_1,
        ptr_deref_1009_load_0_ack_1,
        "ptr_deref_1009_load_0",
        "memory_space_16" ,
        ptr_deref_1009_data_0,
        ptr_deref_1009_word_address_0,
        "ptr_deref_1009_data_0",
        "ptr_deref_1009_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1009_load_0_req_0;
      ptr_deref_1009_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1009_load_0_req_1;
      ptr_deref_1009_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1009_word_address_0;
      ptr_deref_1009_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_16_lr_req(0),
          mack => memory_space_16_lr_ack(0),
          maddr => memory_space_16_lr_addr(0 downto 0),
          mtag => memory_space_16_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_16_lc_req(0),
          mack => memory_space_16_lc_ack(0),
          mdata => memory_space_16_lc_data(31 downto 0),
          mtag => memory_space_16_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_687_load_0_req_0,ptr_deref_687_load_0_ack_0,ptr_deref_687_load_0_req_1,ptr_deref_687_load_0_ack_1,sl_one,"ptr_deref_687_load_0",false,ptr_deref_687_word_address_0,
    false,ptr_deref_687_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_704_load_0_req_0,ptr_deref_704_load_0_ack_0,ptr_deref_704_load_0_req_1,ptr_deref_704_load_0_ack_1,sl_one,"ptr_deref_704_load_0",false,ptr_deref_704_word_address_0,
    false,ptr_deref_704_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1013_load_0_req_0,ptr_deref_1013_load_0_ack_0,ptr_deref_1013_load_0_req_1,ptr_deref_1013_load_0_ack_1,sl_one,"ptr_deref_1013_load_0",false,ptr_deref_1013_word_address_0,
    false,ptr_deref_1013_data_0);
    -- shared load operator group (1) : ptr_deref_687_load_0 ptr_deref_704_load_0 ptr_deref_1013_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_687_load_0_req_0,
        ptr_deref_687_load_0_ack_0,
        ptr_deref_687_load_0_req_1,
        ptr_deref_687_load_0_ack_1,
        "ptr_deref_687_load_0",
        "memory_space_8" ,
        ptr_deref_687_data_0,
        ptr_deref_687_word_address_0,
        "ptr_deref_687_data_0",
        "ptr_deref_687_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_704_load_0_req_0,
        ptr_deref_704_load_0_ack_0,
        ptr_deref_704_load_0_req_1,
        ptr_deref_704_load_0_ack_1,
        "ptr_deref_704_load_0",
        "memory_space_8" ,
        ptr_deref_704_data_0,
        ptr_deref_704_word_address_0,
        "ptr_deref_704_data_0",
        "ptr_deref_704_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1013_load_0_req_0,
        ptr_deref_1013_load_0_ack_0,
        ptr_deref_1013_load_0_req_1,
        ptr_deref_1013_load_0_ack_1,
        "ptr_deref_1013_load_0",
        "memory_space_8" ,
        ptr_deref_1013_data_0,
        ptr_deref_1013_word_address_0,
        "ptr_deref_1013_data_0",
        "ptr_deref_1013_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_687_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_704_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1013_load_0_req_0;
      ptr_deref_687_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_704_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1013_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_687_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_704_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1013_load_0_req_1;
      ptr_deref_687_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_704_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1013_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_687_word_address_0 & ptr_deref_704_word_address_0 & ptr_deref_1013_word_address_0;
      ptr_deref_687_data_0 <= data_out(23 downto 16);
      ptr_deref_704_data_0 <= data_out(15 downto 8);
      ptr_deref_1013_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(7 downto 0),
          mtag => memory_space_8_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1030_load_0_req_0,ptr_deref_1030_load_0_ack_0,ptr_deref_1030_load_0_req_1,ptr_deref_1030_load_0_ack_1,sl_one,"ptr_deref_1030_load_0",false,ptr_deref_1030_word_address_0,
    false,ptr_deref_1030_data_0);
    -- shared load operator group (2) : ptr_deref_1030_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1030_load_0_req_0,
        ptr_deref_1030_load_0_ack_0,
        ptr_deref_1030_load_0_req_1,
        ptr_deref_1030_load_0_ack_1,
        "ptr_deref_1030_load_0",
        "memory_space_17" ,
        ptr_deref_1030_data_0,
        ptr_deref_1030_word_address_0,
        "ptr_deref_1030_data_0",
        "ptr_deref_1030_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1030_load_0_req_0;
      ptr_deref_1030_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1030_load_0_req_1;
      ptr_deref_1030_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1030_word_address_0;
      ptr_deref_1030_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_17_lr_req(0),
          mack => memory_space_17_lr_ack(0),
          maddr => memory_space_17_lr_addr(0 downto 0),
          mtag => memory_space_17_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_17_lc_req(0),
          mack => memory_space_17_lc_ack(0),
          mdata => memory_space_17_lc_data(31 downto 0),
          mtag => memory_space_17_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1034_load_0_req_0,ptr_deref_1034_load_0_ack_0,ptr_deref_1034_load_0_req_1,ptr_deref_1034_load_0_ack_1,sl_one,"ptr_deref_1034_load_0",false,ptr_deref_1034_word_address_0,
    false,ptr_deref_1034_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_747_load_0_req_0,ptr_deref_747_load_0_ack_0,ptr_deref_747_load_0_req_1,ptr_deref_747_load_0_ack_1,sl_one,"ptr_deref_747_load_0",false,ptr_deref_747_word_address_0,
    false,ptr_deref_747_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_730_load_0_req_0,ptr_deref_730_load_0_ack_0,ptr_deref_730_load_0_req_1,ptr_deref_730_load_0_ack_1,sl_one,"ptr_deref_730_load_0",false,ptr_deref_730_word_address_0,
    false,ptr_deref_730_data_0);
    -- shared load operator group (3) : ptr_deref_1034_load_0 ptr_deref_747_load_0 ptr_deref_730_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1034_load_0_req_0,
        ptr_deref_1034_load_0_ack_0,
        ptr_deref_1034_load_0_req_1,
        ptr_deref_1034_load_0_ack_1,
        "ptr_deref_1034_load_0",
        "memory_space_9" ,
        ptr_deref_1034_data_0,
        ptr_deref_1034_word_address_0,
        "ptr_deref_1034_data_0",
        "ptr_deref_1034_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_747_load_0_req_0,
        ptr_deref_747_load_0_ack_0,
        ptr_deref_747_load_0_req_1,
        ptr_deref_747_load_0_ack_1,
        "ptr_deref_747_load_0",
        "memory_space_9" ,
        ptr_deref_747_data_0,
        ptr_deref_747_word_address_0,
        "ptr_deref_747_data_0",
        "ptr_deref_747_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_730_load_0_req_0,
        ptr_deref_730_load_0_ack_0,
        ptr_deref_730_load_0_req_1,
        ptr_deref_730_load_0_ack_1,
        "ptr_deref_730_load_0",
        "memory_space_9" ,
        ptr_deref_730_data_0,
        ptr_deref_730_word_address_0,
        "ptr_deref_730_data_0",
        "ptr_deref_730_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1034_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_747_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_730_load_0_req_0;
      ptr_deref_1034_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_747_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_730_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1034_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_747_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_730_load_0_req_1;
      ptr_deref_1034_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_747_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_730_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1034_word_address_0 & ptr_deref_747_word_address_0 & ptr_deref_730_word_address_0;
      ptr_deref_1034_data_0 <= data_out(23 downto 16);
      ptr_deref_747_data_0 <= data_out(15 downto 8);
      ptr_deref_730_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(0 downto 0),
          mtag => memory_space_9_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(7 downto 0),
          mtag => memory_space_9_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1051_load_0_req_0,ptr_deref_1051_load_0_ack_0,ptr_deref_1051_load_0_req_1,ptr_deref_1051_load_0_ack_1,sl_one,"ptr_deref_1051_load_0",false,ptr_deref_1051_word_address_0,
    false,ptr_deref_1051_data_0);
    -- shared load operator group (4) : ptr_deref_1051_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1051_load_0_req_0,
        ptr_deref_1051_load_0_ack_0,
        ptr_deref_1051_load_0_req_1,
        ptr_deref_1051_load_0_ack_1,
        "ptr_deref_1051_load_0",
        "memory_space_18" ,
        ptr_deref_1051_data_0,
        ptr_deref_1051_word_address_0,
        "ptr_deref_1051_data_0",
        "ptr_deref_1051_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1051_load_0_req_0;
      ptr_deref_1051_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1051_load_0_req_1;
      ptr_deref_1051_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1051_word_address_0;
      ptr_deref_1051_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_18_lr_req(0),
          mack => memory_space_18_lr_ack(0),
          maddr => memory_space_18_lr_addr(0 downto 0),
          mtag => memory_space_18_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_18_lc_req(0),
          mack => memory_space_18_lc_ack(0),
          mdata => memory_space_18_lc_data(31 downto 0),
          mtag => memory_space_18_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1055_load_0_req_0,ptr_deref_1055_load_0_ack_0,ptr_deref_1055_load_0_req_1,ptr_deref_1055_load_0_ack_1,sl_one,"ptr_deref_1055_load_0",false,ptr_deref_1055_word_address_0,
    false,ptr_deref_1055_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_790_load_0_req_0,ptr_deref_790_load_0_ack_0,ptr_deref_790_load_0_req_1,ptr_deref_790_load_0_ack_1,sl_one,"ptr_deref_790_load_0",false,ptr_deref_790_word_address_0,
    false,ptr_deref_790_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_773_load_0_req_0,ptr_deref_773_load_0_ack_0,ptr_deref_773_load_0_req_1,ptr_deref_773_load_0_ack_1,sl_one,"ptr_deref_773_load_0",false,ptr_deref_773_word_address_0,
    false,ptr_deref_773_data_0);
    -- shared load operator group (5) : ptr_deref_1055_load_0 ptr_deref_790_load_0 ptr_deref_773_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1055_load_0_req_0,
        ptr_deref_1055_load_0_ack_0,
        ptr_deref_1055_load_0_req_1,
        ptr_deref_1055_load_0_ack_1,
        "ptr_deref_1055_load_0",
        "memory_space_10" ,
        ptr_deref_1055_data_0,
        ptr_deref_1055_word_address_0,
        "ptr_deref_1055_data_0",
        "ptr_deref_1055_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_790_load_0_req_0,
        ptr_deref_790_load_0_ack_0,
        ptr_deref_790_load_0_req_1,
        ptr_deref_790_load_0_ack_1,
        "ptr_deref_790_load_0",
        "memory_space_10" ,
        ptr_deref_790_data_0,
        ptr_deref_790_word_address_0,
        "ptr_deref_790_data_0",
        "ptr_deref_790_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_773_load_0_req_0,
        ptr_deref_773_load_0_ack_0,
        ptr_deref_773_load_0_req_1,
        ptr_deref_773_load_0_ack_1,
        "ptr_deref_773_load_0",
        "memory_space_10" ,
        ptr_deref_773_data_0,
        ptr_deref_773_word_address_0,
        "ptr_deref_773_data_0",
        "ptr_deref_773_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1055_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_790_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_773_load_0_req_0;
      ptr_deref_1055_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_790_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_773_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1055_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_790_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_773_load_0_req_1;
      ptr_deref_1055_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_790_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_773_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1055_word_address_0 & ptr_deref_790_word_address_0 & ptr_deref_773_word_address_0;
      ptr_deref_1055_data_0 <= data_out(23 downto 16);
      ptr_deref_790_data_0 <= data_out(15 downto 8);
      ptr_deref_773_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_10_lr_req(0),
          mack => memory_space_10_lr_ack(0),
          maddr => memory_space_10_lr_addr(0 downto 0),
          mtag => memory_space_10_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_10_lc_req(0),
          mack => memory_space_10_lc_ack(0),
          mdata => memory_space_10_lc_data(7 downto 0),
          mtag => memory_space_10_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1072_load_0_req_0,ptr_deref_1072_load_0_ack_0,ptr_deref_1072_load_0_req_1,ptr_deref_1072_load_0_ack_1,sl_one,"ptr_deref_1072_load_0",false,ptr_deref_1072_word_address_0,
    false,ptr_deref_1072_data_0);
    -- shared load operator group (6) : ptr_deref_1072_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1072_load_0_req_0,
        ptr_deref_1072_load_0_ack_0,
        ptr_deref_1072_load_0_req_1,
        ptr_deref_1072_load_0_ack_1,
        "ptr_deref_1072_load_0",
        "memory_space_19" ,
        ptr_deref_1072_data_0,
        ptr_deref_1072_word_address_0,
        "ptr_deref_1072_data_0",
        "ptr_deref_1072_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1072_load_0_req_0;
      ptr_deref_1072_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1072_load_0_req_1;
      ptr_deref_1072_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1072_word_address_0;
      ptr_deref_1072_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_19_lr_req(0),
          mack => memory_space_19_lr_ack(0),
          maddr => memory_space_19_lr_addr(0 downto 0),
          mtag => memory_space_19_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_19_lc_req(0),
          mack => memory_space_19_lc_ack(0),
          mdata => memory_space_19_lc_data(31 downto 0),
          mtag => memory_space_19_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1076_load_0_req_0,ptr_deref_1076_load_0_ack_0,ptr_deref_1076_load_0_req_1,ptr_deref_1076_load_0_ack_1,sl_one,"ptr_deref_1076_load_0",false,ptr_deref_1076_word_address_0,
    false,ptr_deref_1076_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_816_load_0_req_0,ptr_deref_816_load_0_ack_0,ptr_deref_816_load_0_req_1,ptr_deref_816_load_0_ack_1,sl_one,"ptr_deref_816_load_0",false,ptr_deref_816_word_address_0,
    false,ptr_deref_816_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_833_load_0_req_0,ptr_deref_833_load_0_ack_0,ptr_deref_833_load_0_req_1,ptr_deref_833_load_0_ack_1,sl_one,"ptr_deref_833_load_0",false,ptr_deref_833_word_address_0,
    false,ptr_deref_833_data_0);
    -- shared load operator group (7) : ptr_deref_1076_load_0 ptr_deref_816_load_0 ptr_deref_833_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1076_load_0_req_0,
        ptr_deref_1076_load_0_ack_0,
        ptr_deref_1076_load_0_req_1,
        ptr_deref_1076_load_0_ack_1,
        "ptr_deref_1076_load_0",
        "memory_space_11" ,
        ptr_deref_1076_data_0,
        ptr_deref_1076_word_address_0,
        "ptr_deref_1076_data_0",
        "ptr_deref_1076_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_816_load_0_req_0,
        ptr_deref_816_load_0_ack_0,
        ptr_deref_816_load_0_req_1,
        ptr_deref_816_load_0_ack_1,
        "ptr_deref_816_load_0",
        "memory_space_11" ,
        ptr_deref_816_data_0,
        ptr_deref_816_word_address_0,
        "ptr_deref_816_data_0",
        "ptr_deref_816_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_833_load_0_req_0,
        ptr_deref_833_load_0_ack_0,
        ptr_deref_833_load_0_req_1,
        ptr_deref_833_load_0_ack_1,
        "ptr_deref_833_load_0",
        "memory_space_11" ,
        ptr_deref_833_data_0,
        ptr_deref_833_word_address_0,
        "ptr_deref_833_data_0",
        "ptr_deref_833_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1076_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_816_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_833_load_0_req_0;
      ptr_deref_1076_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_816_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_833_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1076_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_816_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_833_load_0_req_1;
      ptr_deref_1076_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_816_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_833_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1076_word_address_0 & ptr_deref_816_word_address_0 & ptr_deref_833_word_address_0;
      ptr_deref_1076_data_0 <= data_out(23 downto 16);
      ptr_deref_816_data_0 <= data_out(15 downto 8);
      ptr_deref_833_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_11_lr_req(0),
          mack => memory_space_11_lr_ack(0),
          maddr => memory_space_11_lr_addr(0 downto 0),
          mtag => memory_space_11_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_11_lc_req(0),
          mack => memory_space_11_lc_ack(0),
          mdata => memory_space_11_lc_data(7 downto 0),
          mtag => memory_space_11_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1093_load_0_req_0,ptr_deref_1093_load_0_ack_0,ptr_deref_1093_load_0_req_1,ptr_deref_1093_load_0_ack_1,sl_one,"ptr_deref_1093_load_0",false,ptr_deref_1093_word_address_0,
    false,ptr_deref_1093_data_0);
    -- shared load operator group (8) : ptr_deref_1093_load_0 
    LoadGroup8: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1093_load_0_req_0,
        ptr_deref_1093_load_0_ack_0,
        ptr_deref_1093_load_0_req_1,
        ptr_deref_1093_load_0_ack_1,
        "ptr_deref_1093_load_0",
        "memory_space_20" ,
        ptr_deref_1093_data_0,
        ptr_deref_1093_word_address_0,
        "ptr_deref_1093_data_0",
        "ptr_deref_1093_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1093_load_0_req_0;
      ptr_deref_1093_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1093_load_0_req_1;
      ptr_deref_1093_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1093_word_address_0;
      ptr_deref_1093_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_20_lr_req(0),
          mack => memory_space_20_lr_ack(0),
          maddr => memory_space_20_lr_addr(0 downto 0),
          mtag => memory_space_20_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_20_lc_req(0),
          mack => memory_space_20_lc_ack(0),
          mdata => memory_space_20_lc_data(31 downto 0),
          mtag => memory_space_20_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 8
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1097_load_0_req_0,ptr_deref_1097_load_0_ack_0,ptr_deref_1097_load_0_req_1,ptr_deref_1097_load_0_ack_1,sl_one,"ptr_deref_1097_load_0",false,ptr_deref_1097_word_address_0,
    false,ptr_deref_1097_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_859_load_0_req_0,ptr_deref_859_load_0_ack_0,ptr_deref_859_load_0_req_1,ptr_deref_859_load_0_ack_1,sl_one,"ptr_deref_859_load_0",false,ptr_deref_859_word_address_0,
    false,ptr_deref_859_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_876_load_0_req_0,ptr_deref_876_load_0_ack_0,ptr_deref_876_load_0_req_1,ptr_deref_876_load_0_ack_1,sl_one,"ptr_deref_876_load_0",false,ptr_deref_876_word_address_0,
    false,ptr_deref_876_data_0);
    -- shared load operator group (9) : ptr_deref_1097_load_0 ptr_deref_859_load_0 ptr_deref_876_load_0 
    LoadGroup9: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1097_load_0_req_0,
        ptr_deref_1097_load_0_ack_0,
        ptr_deref_1097_load_0_req_1,
        ptr_deref_1097_load_0_ack_1,
        "ptr_deref_1097_load_0",
        "memory_space_12" ,
        ptr_deref_1097_data_0,
        ptr_deref_1097_word_address_0,
        "ptr_deref_1097_data_0",
        "ptr_deref_1097_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_859_load_0_req_0,
        ptr_deref_859_load_0_ack_0,
        ptr_deref_859_load_0_req_1,
        ptr_deref_859_load_0_ack_1,
        "ptr_deref_859_load_0",
        "memory_space_12" ,
        ptr_deref_859_data_0,
        ptr_deref_859_word_address_0,
        "ptr_deref_859_data_0",
        "ptr_deref_859_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_876_load_0_req_0,
        ptr_deref_876_load_0_ack_0,
        ptr_deref_876_load_0_req_1,
        ptr_deref_876_load_0_ack_1,
        "ptr_deref_876_load_0",
        "memory_space_12" ,
        ptr_deref_876_data_0,
        ptr_deref_876_word_address_0,
        "ptr_deref_876_data_0",
        "ptr_deref_876_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1097_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_859_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_876_load_0_req_0;
      ptr_deref_1097_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_859_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_876_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1097_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_859_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_876_load_0_req_1;
      ptr_deref_1097_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_859_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_876_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1097_word_address_0 & ptr_deref_859_word_address_0 & ptr_deref_876_word_address_0;
      ptr_deref_1097_data_0 <= data_out(23 downto 16);
      ptr_deref_859_data_0 <= data_out(15 downto 8);
      ptr_deref_876_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_12_lr_req(0),
          mack => memory_space_12_lr_ack(0),
          maddr => memory_space_12_lr_addr(0 downto 0),
          mtag => memory_space_12_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_12_lc_req(0),
          mack => memory_space_12_lc_ack(0),
          mdata => memory_space_12_lc_data(7 downto 0),
          mtag => memory_space_12_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 9
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1114_load_0_req_0,ptr_deref_1114_load_0_ack_0,ptr_deref_1114_load_0_req_1,ptr_deref_1114_load_0_ack_1,sl_one,"ptr_deref_1114_load_0",false,ptr_deref_1114_word_address_0,
    false,ptr_deref_1114_data_0);
    -- shared load operator group (10) : ptr_deref_1114_load_0 
    LoadGroup10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1114_load_0_req_0,
        ptr_deref_1114_load_0_ack_0,
        ptr_deref_1114_load_0_req_1,
        ptr_deref_1114_load_0_ack_1,
        "ptr_deref_1114_load_0",
        "memory_space_21" ,
        ptr_deref_1114_data_0,
        ptr_deref_1114_word_address_0,
        "ptr_deref_1114_data_0",
        "ptr_deref_1114_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1114_load_0_req_0;
      ptr_deref_1114_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1114_load_0_req_1;
      ptr_deref_1114_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1114_word_address_0;
      ptr_deref_1114_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_21_lr_req(0),
          mack => memory_space_21_lr_ack(0),
          maddr => memory_space_21_lr_addr(0 downto 0),
          mtag => memory_space_21_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_21_lc_req(0),
          mack => memory_space_21_lc_ack(0),
          mdata => memory_space_21_lc_data(31 downto 0),
          mtag => memory_space_21_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 10
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1118_load_0_req_0,ptr_deref_1118_load_0_ack_0,ptr_deref_1118_load_0_req_1,ptr_deref_1118_load_0_ack_1,sl_one,"ptr_deref_1118_load_0",false,ptr_deref_1118_word_address_0,
    false,ptr_deref_1118_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_902_load_0_req_0,ptr_deref_902_load_0_ack_0,ptr_deref_902_load_0_req_1,ptr_deref_902_load_0_ack_1,sl_one,"ptr_deref_902_load_0",false,ptr_deref_902_word_address_0,
    false,ptr_deref_902_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_919_load_0_req_0,ptr_deref_919_load_0_ack_0,ptr_deref_919_load_0_req_1,ptr_deref_919_load_0_ack_1,sl_one,"ptr_deref_919_load_0",false,ptr_deref_919_word_address_0,
    false,ptr_deref_919_data_0);
    -- shared load operator group (11) : ptr_deref_1118_load_0 ptr_deref_902_load_0 ptr_deref_919_load_0 
    LoadGroup11: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1118_load_0_req_0,
        ptr_deref_1118_load_0_ack_0,
        ptr_deref_1118_load_0_req_1,
        ptr_deref_1118_load_0_ack_1,
        "ptr_deref_1118_load_0",
        "memory_space_13" ,
        ptr_deref_1118_data_0,
        ptr_deref_1118_word_address_0,
        "ptr_deref_1118_data_0",
        "ptr_deref_1118_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_902_load_0_req_0,
        ptr_deref_902_load_0_ack_0,
        ptr_deref_902_load_0_req_1,
        ptr_deref_902_load_0_ack_1,
        "ptr_deref_902_load_0",
        "memory_space_13" ,
        ptr_deref_902_data_0,
        ptr_deref_902_word_address_0,
        "ptr_deref_902_data_0",
        "ptr_deref_902_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_919_load_0_req_0,
        ptr_deref_919_load_0_ack_0,
        ptr_deref_919_load_0_req_1,
        ptr_deref_919_load_0_ack_1,
        "ptr_deref_919_load_0",
        "memory_space_13" ,
        ptr_deref_919_data_0,
        ptr_deref_919_word_address_0,
        "ptr_deref_919_data_0",
        "ptr_deref_919_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1118_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_902_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_919_load_0_req_0;
      ptr_deref_1118_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_902_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_919_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1118_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_902_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_919_load_0_req_1;
      ptr_deref_1118_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_902_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_919_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1118_word_address_0 & ptr_deref_902_word_address_0 & ptr_deref_919_word_address_0;
      ptr_deref_1118_data_0 <= data_out(23 downto 16);
      ptr_deref_902_data_0 <= data_out(15 downto 8);
      ptr_deref_919_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_13_lr_req(0),
          mack => memory_space_13_lr_ack(0),
          maddr => memory_space_13_lr_addr(0 downto 0),
          mtag => memory_space_13_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_13_lc_req(0),
          mack => memory_space_13_lc_ack(0),
          mdata => memory_space_13_lc_data(7 downto 0),
          mtag => memory_space_13_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 11
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1135_load_0_req_0,ptr_deref_1135_load_0_ack_0,ptr_deref_1135_load_0_req_1,ptr_deref_1135_load_0_ack_1,sl_one,"ptr_deref_1135_load_0",false,ptr_deref_1135_word_address_0,
    false,ptr_deref_1135_data_0);
    -- shared load operator group (12) : ptr_deref_1135_load_0 
    LoadGroup12: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1135_load_0_req_0,
        ptr_deref_1135_load_0_ack_0,
        ptr_deref_1135_load_0_req_1,
        ptr_deref_1135_load_0_ack_1,
        "ptr_deref_1135_load_0",
        "memory_space_22" ,
        ptr_deref_1135_data_0,
        ptr_deref_1135_word_address_0,
        "ptr_deref_1135_data_0",
        "ptr_deref_1135_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_1135_load_0_req_0;
      ptr_deref_1135_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_1135_load_0_req_1;
      ptr_deref_1135_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1135_word_address_0;
      ptr_deref_1135_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_22_lr_req(0),
          mack => memory_space_22_lr_ack(0),
          maddr => memory_space_22_lr_addr(0 downto 0),
          mtag => memory_space_22_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_22_lc_req(0),
          mack => memory_space_22_lc_ack(0),
          mdata => memory_space_22_lc_data(31 downto 0),
          mtag => memory_space_22_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 12
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1139_load_0_req_0,ptr_deref_1139_load_0_ack_0,ptr_deref_1139_load_0_req_1,ptr_deref_1139_load_0_ack_1,sl_one,"ptr_deref_1139_load_0",false,ptr_deref_1139_word_address_0,
    false,ptr_deref_1139_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_962_load_0_req_0,ptr_deref_962_load_0_ack_0,ptr_deref_962_load_0_req_1,ptr_deref_962_load_0_ack_1,sl_one,"ptr_deref_962_load_0",false,ptr_deref_962_word_address_0,
    false,ptr_deref_962_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_945_load_0_req_0,ptr_deref_945_load_0_ack_0,ptr_deref_945_load_0_req_1,ptr_deref_945_load_0_ack_1,sl_one,"ptr_deref_945_load_0",false,ptr_deref_945_word_address_0,
    false,ptr_deref_945_data_0);
    -- shared load operator group (13) : ptr_deref_1139_load_0 ptr_deref_962_load_0 ptr_deref_945_load_0 
    LoadGroup13: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 2 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 2 downto 0);
      signal guard_vector : std_logic_vector( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1139_load_0_req_0,
        ptr_deref_1139_load_0_ack_0,
        ptr_deref_1139_load_0_req_1,
        ptr_deref_1139_load_0_ack_1,
        "ptr_deref_1139_load_0",
        "memory_space_14" ,
        ptr_deref_1139_data_0,
        ptr_deref_1139_word_address_0,
        "ptr_deref_1139_data_0",
        "ptr_deref_1139_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_962_load_0_req_0,
        ptr_deref_962_load_0_ack_0,
        ptr_deref_962_load_0_req_1,
        ptr_deref_962_load_0_ack_1,
        "ptr_deref_962_load_0",
        "memory_space_14" ,
        ptr_deref_962_data_0,
        ptr_deref_962_word_address_0,
        "ptr_deref_962_data_0",
        "ptr_deref_962_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_945_load_0_req_0,
        ptr_deref_945_load_0_ack_0,
        ptr_deref_945_load_0_req_1,
        ptr_deref_945_load_0_ack_1,
        "ptr_deref_945_load_0",
        "memory_space_14" ,
        ptr_deref_945_data_0,
        ptr_deref_945_word_address_0,
        "ptr_deref_945_data_0",
        "ptr_deref_945_word_address_0" -- 
      );
      reqL_unguarded(2) <= ptr_deref_1139_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_962_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_945_load_0_req_0;
      ptr_deref_1139_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_962_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_945_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(2) <= ptr_deref_1139_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_962_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_945_load_0_req_1;
      ptr_deref_1139_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_962_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_945_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 3) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_1139_word_address_0 & ptr_deref_962_word_address_0 & ptr_deref_945_word_address_0;
      ptr_deref_1139_data_0 <= data_out(23 downto 16);
      ptr_deref_962_data_0 <= data_out(15 downto 8);
      ptr_deref_945_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_14_lr_req(0),
          mack => memory_space_14_lr_ack(0),
          maddr => memory_space_14_lr_addr(0 downto 0),
          mtag => memory_space_14_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_14_lc_req(0),
          mack => memory_space_14_lc_ack(0),
          mdata => memory_space_14_lc_data(7 downto 0),
          mtag => memory_space_14_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 13
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_600_load_0_req_0,ptr_deref_600_load_0_ack_0,ptr_deref_600_load_0_req_1,ptr_deref_600_load_0_ack_1,sl_one,"ptr_deref_600_load_0",false,ptr_deref_600_word_address_0,
    false,ptr_deref_600_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_512_load_0_req_0,ptr_deref_512_load_0_ack_0,ptr_deref_512_load_0_req_1,ptr_deref_512_load_0_ack_1,sl_one,"ptr_deref_512_load_0",false,ptr_deref_512_word_address_0,
    false,ptr_deref_512_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_490_load_0_req_0,ptr_deref_490_load_0_ack_0,ptr_deref_490_load_0_req_1,ptr_deref_490_load_0_ack_1,sl_one,"ptr_deref_490_load_0",false,ptr_deref_490_word_address_0,
    false,ptr_deref_490_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_661_load_0_req_0,ptr_deref_661_load_0_ack_0,ptr_deref_661_load_0_req_1,ptr_deref_661_load_0_ack_1,sl_one,"ptr_deref_661_load_0",false,ptr_deref_661_word_address_0,
    false,ptr_deref_661_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_578_load_0_req_0,ptr_deref_578_load_0_ack_0,ptr_deref_578_load_0_req_1,ptr_deref_578_load_0_ack_1,sl_one,"ptr_deref_578_load_0",false,ptr_deref_578_word_address_0,
    false,ptr_deref_578_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_622_load_0_req_0,ptr_deref_622_load_0_ack_0,ptr_deref_622_load_0_req_1,ptr_deref_622_load_0_ack_1,sl_one,"ptr_deref_622_load_0",false,ptr_deref_622_word_address_0,
    false,ptr_deref_622_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_644_load_0_req_0,ptr_deref_644_load_0_ack_0,ptr_deref_644_load_0_req_1,ptr_deref_644_load_0_ack_1,sl_one,"ptr_deref_644_load_0",false,ptr_deref_644_word_address_0,
    false,ptr_deref_644_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_467_load_0_req_0,ptr_deref_467_load_0_ack_0,ptr_deref_467_load_0_req_1,ptr_deref_467_load_0_ack_1,sl_one,"ptr_deref_467_load_0",false,ptr_deref_467_word_address_0,
    false,ptr_deref_467_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_534_load_0_req_0,ptr_deref_534_load_0_ack_0,ptr_deref_534_load_0_req_1,ptr_deref_534_load_0_ack_1,sl_one,"ptr_deref_534_load_0",false,ptr_deref_534_word_address_0,
    false,ptr_deref_534_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_556_load_0_req_0,ptr_deref_556_load_0_ack_0,ptr_deref_556_load_0_req_1,ptr_deref_556_load_0_ack_1,sl_one,"ptr_deref_556_load_0",false,ptr_deref_556_word_address_0,
    false,ptr_deref_556_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_992_load_0_req_0,ptr_deref_992_load_0_ack_0,ptr_deref_992_load_0_req_1,ptr_deref_992_load_0_ack_1,sl_one,"ptr_deref_992_load_0",false,ptr_deref_992_word_address_0,
    false,ptr_deref_992_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1158_load_0_req_0,ptr_deref_1158_load_0_ack_0,ptr_deref_1158_load_0_req_1,ptr_deref_1158_load_0_ack_1,sl_one,"ptr_deref_1158_load_0",false,ptr_deref_1158_word_address_0,
    false,ptr_deref_1158_data_0);
    -- shared load operator group (14) : ptr_deref_600_load_0 ptr_deref_512_load_0 ptr_deref_490_load_0 ptr_deref_661_load_0 ptr_deref_578_load_0 ptr_deref_622_load_0 ptr_deref_644_load_0 ptr_deref_467_load_0 ptr_deref_534_load_0 ptr_deref_556_load_0 ptr_deref_992_load_0 ptr_deref_1158_load_0 
    LoadGroup14: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 11 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 11 downto 0);
      signal guard_vector : std_logic_vector( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_600_load_0_req_0,
        ptr_deref_600_load_0_ack_0,
        ptr_deref_600_load_0_req_1,
        ptr_deref_600_load_0_ack_1,
        "ptr_deref_600_load_0",
        "memory_space_7" ,
        ptr_deref_600_data_0,
        ptr_deref_600_word_address_0,
        "ptr_deref_600_data_0",
        "ptr_deref_600_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_512_load_0_req_0,
        ptr_deref_512_load_0_ack_0,
        ptr_deref_512_load_0_req_1,
        ptr_deref_512_load_0_ack_1,
        "ptr_deref_512_load_0",
        "memory_space_7" ,
        ptr_deref_512_data_0,
        ptr_deref_512_word_address_0,
        "ptr_deref_512_data_0",
        "ptr_deref_512_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_490_load_0_req_0,
        ptr_deref_490_load_0_ack_0,
        ptr_deref_490_load_0_req_1,
        ptr_deref_490_load_0_ack_1,
        "ptr_deref_490_load_0",
        "memory_space_7" ,
        ptr_deref_490_data_0,
        ptr_deref_490_word_address_0,
        "ptr_deref_490_data_0",
        "ptr_deref_490_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_661_load_0_req_0,
        ptr_deref_661_load_0_ack_0,
        ptr_deref_661_load_0_req_1,
        ptr_deref_661_load_0_ack_1,
        "ptr_deref_661_load_0",
        "memory_space_7" ,
        ptr_deref_661_data_0,
        ptr_deref_661_word_address_0,
        "ptr_deref_661_data_0",
        "ptr_deref_661_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_578_load_0_req_0,
        ptr_deref_578_load_0_ack_0,
        ptr_deref_578_load_0_req_1,
        ptr_deref_578_load_0_ack_1,
        "ptr_deref_578_load_0",
        "memory_space_7" ,
        ptr_deref_578_data_0,
        ptr_deref_578_word_address_0,
        "ptr_deref_578_data_0",
        "ptr_deref_578_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_622_load_0_req_0,
        ptr_deref_622_load_0_ack_0,
        ptr_deref_622_load_0_req_1,
        ptr_deref_622_load_0_ack_1,
        "ptr_deref_622_load_0",
        "memory_space_7" ,
        ptr_deref_622_data_0,
        ptr_deref_622_word_address_0,
        "ptr_deref_622_data_0",
        "ptr_deref_622_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_644_load_0_req_0,
        ptr_deref_644_load_0_ack_0,
        ptr_deref_644_load_0_req_1,
        ptr_deref_644_load_0_ack_1,
        "ptr_deref_644_load_0",
        "memory_space_7" ,
        ptr_deref_644_data_0,
        ptr_deref_644_word_address_0,
        "ptr_deref_644_data_0",
        "ptr_deref_644_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_467_load_0_req_0,
        ptr_deref_467_load_0_ack_0,
        ptr_deref_467_load_0_req_1,
        ptr_deref_467_load_0_ack_1,
        "ptr_deref_467_load_0",
        "memory_space_7" ,
        ptr_deref_467_data_0,
        ptr_deref_467_word_address_0,
        "ptr_deref_467_data_0",
        "ptr_deref_467_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_534_load_0_req_0,
        ptr_deref_534_load_0_ack_0,
        ptr_deref_534_load_0_req_1,
        ptr_deref_534_load_0_ack_1,
        "ptr_deref_534_load_0",
        "memory_space_7" ,
        ptr_deref_534_data_0,
        ptr_deref_534_word_address_0,
        "ptr_deref_534_data_0",
        "ptr_deref_534_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_556_load_0_req_0,
        ptr_deref_556_load_0_ack_0,
        ptr_deref_556_load_0_req_1,
        ptr_deref_556_load_0_ack_1,
        "ptr_deref_556_load_0",
        "memory_space_7" ,
        ptr_deref_556_data_0,
        ptr_deref_556_word_address_0,
        "ptr_deref_556_data_0",
        "ptr_deref_556_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_992_load_0_req_0,
        ptr_deref_992_load_0_ack_0,
        ptr_deref_992_load_0_req_1,
        ptr_deref_992_load_0_ack_1,
        "ptr_deref_992_load_0",
        "memory_space_7" ,
        ptr_deref_992_data_0,
        ptr_deref_992_word_address_0,
        "ptr_deref_992_data_0",
        "ptr_deref_992_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_1158_load_0_req_0,
        ptr_deref_1158_load_0_ack_0,
        ptr_deref_1158_load_0_req_1,
        ptr_deref_1158_load_0_ack_1,
        "ptr_deref_1158_load_0",
        "memory_space_7" ,
        ptr_deref_1158_data_0,
        ptr_deref_1158_word_address_0,
        "ptr_deref_1158_data_0",
        "ptr_deref_1158_word_address_0" -- 
      );
      reqL_unguarded(11) <= ptr_deref_600_load_0_req_0;
      reqL_unguarded(10) <= ptr_deref_512_load_0_req_0;
      reqL_unguarded(9) <= ptr_deref_490_load_0_req_0;
      reqL_unguarded(8) <= ptr_deref_661_load_0_req_0;
      reqL_unguarded(7) <= ptr_deref_578_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_622_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_644_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_467_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_534_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_556_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_992_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1158_load_0_req_0;
      ptr_deref_600_load_0_ack_0 <= ackL_unguarded(11);
      ptr_deref_512_load_0_ack_0 <= ackL_unguarded(10);
      ptr_deref_490_load_0_ack_0 <= ackL_unguarded(9);
      ptr_deref_661_load_0_ack_0 <= ackL_unguarded(8);
      ptr_deref_578_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_622_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_644_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_467_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_534_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_556_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_992_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1158_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(11) <= ptr_deref_600_load_0_req_1;
      reqR_unguarded(10) <= ptr_deref_512_load_0_req_1;
      reqR_unguarded(9) <= ptr_deref_490_load_0_req_1;
      reqR_unguarded(8) <= ptr_deref_661_load_0_req_1;
      reqR_unguarded(7) <= ptr_deref_578_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_622_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_644_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_467_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_534_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_556_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_992_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1158_load_0_req_1;
      ptr_deref_600_load_0_ack_1 <= ackR_unguarded(11);
      ptr_deref_512_load_0_ack_1 <= ackR_unguarded(10);
      ptr_deref_490_load_0_ack_1 <= ackR_unguarded(9);
      ptr_deref_661_load_0_ack_1 <= ackR_unguarded(8);
      ptr_deref_578_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_622_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_644_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_467_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_534_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_556_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_992_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1158_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      guard_vector(8)  <=  '1';
      guard_vector(9)  <=  '1';
      guard_vector(10)  <=  '1';
      guard_vector(11)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 12) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      accessRegulator_8: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(8), -- 
          ack => ackL_unregulated(8),
          regulated_req => reqL(8),
          regulated_ack => ackL(8),
          release_req => reqR(8),
          release_ack => ackR(8),
          clk => clk, reset => reset); -- 
      accessRegulator_9: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(9), -- 
          ack => ackL_unregulated(9),
          regulated_req => reqL(9),
          regulated_ack => ackL(9),
          release_req => reqR(9),
          release_ack => ackR(9),
          clk => clk, reset => reset); -- 
      accessRegulator_10: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(10), -- 
          ack => ackL_unregulated(10),
          regulated_req => reqL(10),
          regulated_ack => ackL(10),
          release_req => reqR(10),
          release_ack => ackR(10),
          clk => clk, reset => reset); -- 
      accessRegulator_11: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(11), -- 
          ack => ackL_unregulated(11),
          regulated_req => reqL(11),
          regulated_ack => ackL(11),
          release_req => reqR(11),
          release_ack => ackR(11),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 12) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_600_word_address_0 & ptr_deref_512_word_address_0 & ptr_deref_490_word_address_0 & ptr_deref_661_word_address_0 & ptr_deref_578_word_address_0 & ptr_deref_622_word_address_0 & ptr_deref_644_word_address_0 & ptr_deref_467_word_address_0 & ptr_deref_534_word_address_0 & ptr_deref_556_word_address_0 & ptr_deref_992_word_address_0 & ptr_deref_1158_word_address_0;
      ptr_deref_600_data_0 <= data_out(95 downto 88);
      ptr_deref_512_data_0 <= data_out(87 downto 80);
      ptr_deref_490_data_0 <= data_out(79 downto 72);
      ptr_deref_661_data_0 <= data_out(71 downto 64);
      ptr_deref_578_data_0 <= data_out(63 downto 56);
      ptr_deref_622_data_0 <= data_out(55 downto 48);
      ptr_deref_644_data_0 <= data_out(47 downto 40);
      ptr_deref_467_data_0 <= data_out(39 downto 32);
      ptr_deref_534_data_0 <= data_out(31 downto 24);
      ptr_deref_556_data_0 <= data_out(23 downto 16);
      ptr_deref_992_data_0 <= data_out(15 downto 8);
      ptr_deref_1158_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 12,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(7 downto 0),
          mtag => memory_space_7_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 14
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_657_load_0_req_0,ptr_deref_657_load_0_ack_0,ptr_deref_657_load_0_req_1,ptr_deref_657_load_0_ack_1,sl_one,"ptr_deref_657_load_0",false,ptr_deref_657_word_address_0,
    false,ptr_deref_657_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_700_load_0_req_0,ptr_deref_700_load_0_ack_0,ptr_deref_700_load_0_req_1,ptr_deref_700_load_0_ack_1,sl_one,"ptr_deref_700_load_0",false,ptr_deref_700_word_address_0,
    false,ptr_deref_700_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_958_load_0_req_0,ptr_deref_958_load_0_ack_0,ptr_deref_958_load_0_req_1,ptr_deref_958_load_0_ack_1,sl_one,"ptr_deref_958_load_0",false,ptr_deref_958_word_address_0,
    false,ptr_deref_958_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_786_load_0_req_0,ptr_deref_786_load_0_ack_0,ptr_deref_786_load_0_req_1,ptr_deref_786_load_0_ack_1,sl_one,"ptr_deref_786_load_0",false,ptr_deref_786_word_address_0,
    false,ptr_deref_786_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_743_load_0_req_0,ptr_deref_743_load_0_ack_0,ptr_deref_743_load_0_req_1,ptr_deref_743_load_0_ack_1,sl_one,"ptr_deref_743_load_0",false,ptr_deref_743_word_address_0,
    false,ptr_deref_743_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_829_load_0_req_0,ptr_deref_829_load_0_ack_0,ptr_deref_829_load_0_req_1,ptr_deref_829_load_0_ack_1,sl_one,"ptr_deref_829_load_0",false,ptr_deref_829_word_address_0,
    false,ptr_deref_829_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_872_load_0_req_0,ptr_deref_872_load_0_ack_0,ptr_deref_872_load_0_req_1,ptr_deref_872_load_0_ack_1,sl_one,"ptr_deref_872_load_0",false,ptr_deref_872_word_address_0,
    false,ptr_deref_872_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_915_load_0_req_0,ptr_deref_915_load_0_ack_0,ptr_deref_915_load_0_req_1,ptr_deref_915_load_0_ack_1,sl_one,"ptr_deref_915_load_0",false,ptr_deref_915_word_address_0,
    false,ptr_deref_915_data_0);
    -- shared load operator group (15) : ptr_deref_657_load_0 ptr_deref_700_load_0 ptr_deref_958_load_0 ptr_deref_786_load_0 ptr_deref_743_load_0 ptr_deref_829_load_0 ptr_deref_872_load_0 ptr_deref_915_load_0 
    LoadGroup15: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_657_load_0_req_0,
        ptr_deref_657_load_0_ack_0,
        ptr_deref_657_load_0_req_1,
        ptr_deref_657_load_0_ack_1,
        "ptr_deref_657_load_0",
        "memory_space_0" ,
        ptr_deref_657_data_0,
        ptr_deref_657_word_address_0,
        "ptr_deref_657_data_0",
        "ptr_deref_657_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_700_load_0_req_0,
        ptr_deref_700_load_0_ack_0,
        ptr_deref_700_load_0_req_1,
        ptr_deref_700_load_0_ack_1,
        "ptr_deref_700_load_0",
        "memory_space_0" ,
        ptr_deref_700_data_0,
        ptr_deref_700_word_address_0,
        "ptr_deref_700_data_0",
        "ptr_deref_700_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_958_load_0_req_0,
        ptr_deref_958_load_0_ack_0,
        ptr_deref_958_load_0_req_1,
        ptr_deref_958_load_0_ack_1,
        "ptr_deref_958_load_0",
        "memory_space_0" ,
        ptr_deref_958_data_0,
        ptr_deref_958_word_address_0,
        "ptr_deref_958_data_0",
        "ptr_deref_958_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_786_load_0_req_0,
        ptr_deref_786_load_0_ack_0,
        ptr_deref_786_load_0_req_1,
        ptr_deref_786_load_0_ack_1,
        "ptr_deref_786_load_0",
        "memory_space_0" ,
        ptr_deref_786_data_0,
        ptr_deref_786_word_address_0,
        "ptr_deref_786_data_0",
        "ptr_deref_786_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_743_load_0_req_0,
        ptr_deref_743_load_0_ack_0,
        ptr_deref_743_load_0_req_1,
        ptr_deref_743_load_0_ack_1,
        "ptr_deref_743_load_0",
        "memory_space_0" ,
        ptr_deref_743_data_0,
        ptr_deref_743_word_address_0,
        "ptr_deref_743_data_0",
        "ptr_deref_743_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_829_load_0_req_0,
        ptr_deref_829_load_0_ack_0,
        ptr_deref_829_load_0_req_1,
        ptr_deref_829_load_0_ack_1,
        "ptr_deref_829_load_0",
        "memory_space_0" ,
        ptr_deref_829_data_0,
        ptr_deref_829_word_address_0,
        "ptr_deref_829_data_0",
        "ptr_deref_829_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_872_load_0_req_0,
        ptr_deref_872_load_0_ack_0,
        ptr_deref_872_load_0_req_1,
        ptr_deref_872_load_0_ack_1,
        "ptr_deref_872_load_0",
        "memory_space_0" ,
        ptr_deref_872_data_0,
        ptr_deref_872_word_address_0,
        "ptr_deref_872_data_0",
        "ptr_deref_872_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_915_load_0_req_0,
        ptr_deref_915_load_0_ack_0,
        ptr_deref_915_load_0_req_1,
        ptr_deref_915_load_0_ack_1,
        "ptr_deref_915_load_0",
        "memory_space_0" ,
        ptr_deref_915_data_0,
        ptr_deref_915_word_address_0,
        "ptr_deref_915_data_0",
        "ptr_deref_915_word_address_0" -- 
      );
      reqL_unguarded(7) <= ptr_deref_657_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_700_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_958_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_786_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_743_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_829_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_872_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_915_load_0_req_0;
      ptr_deref_657_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_700_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_958_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_786_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_743_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_829_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_872_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_915_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_657_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_700_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_958_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_786_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_743_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_829_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_872_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_915_load_0_req_1;
      ptr_deref_657_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_700_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_958_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_786_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_743_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_829_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_872_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_915_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_657_word_address_0 & ptr_deref_700_word_address_0 & ptr_deref_958_word_address_0 & ptr_deref_786_word_address_0 & ptr_deref_743_word_address_0 & ptr_deref_829_word_address_0 & ptr_deref_872_word_address_0 & ptr_deref_915_word_address_0;
      ptr_deref_657_data_0 <= data_out(255 downto 224);
      ptr_deref_700_data_0 <= data_out(223 downto 192);
      ptr_deref_958_data_0 <= data_out(191 downto 160);
      ptr_deref_786_data_0 <= data_out(159 downto 128);
      ptr_deref_743_data_0 <= data_out(127 downto 96);
      ptr_deref_829_data_0 <= data_out(95 downto 64);
      ptr_deref_872_data_0 <= data_out(63 downto 32);
      ptr_deref_915_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 8,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 15
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_717_load_0_req_0,ptr_deref_717_load_0_ack_0,ptr_deref_717_load_0_req_1,ptr_deref_717_load_0_ack_1,sl_one,"ptr_deref_717_load_0",false,ptr_deref_717_word_address_0,
    false,ptr_deref_717_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_674_load_0_req_0,ptr_deref_674_load_0_ack_0,ptr_deref_674_load_0_req_1,ptr_deref_674_load_0_ack_1,sl_one,"ptr_deref_674_load_0",false,ptr_deref_674_word_address_0,
    false,ptr_deref_674_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_975_load_0_req_0,ptr_deref_975_load_0_ack_0,ptr_deref_975_load_0_req_1,ptr_deref_975_load_0_ack_1,sl_one,"ptr_deref_975_load_0",false,ptr_deref_975_word_address_0,
    false,ptr_deref_975_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_760_load_0_req_0,ptr_deref_760_load_0_ack_0,ptr_deref_760_load_0_req_1,ptr_deref_760_load_0_ack_1,sl_one,"ptr_deref_760_load_0",false,ptr_deref_760_word_address_0,
    false,ptr_deref_760_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_803_load_0_req_0,ptr_deref_803_load_0_ack_0,ptr_deref_803_load_0_req_1,ptr_deref_803_load_0_ack_1,sl_one,"ptr_deref_803_load_0",false,ptr_deref_803_word_address_0,
    false,ptr_deref_803_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_846_load_0_req_0,ptr_deref_846_load_0_ack_0,ptr_deref_846_load_0_req_1,ptr_deref_846_load_0_ack_1,sl_one,"ptr_deref_846_load_0",false,ptr_deref_846_word_address_0,
    false,ptr_deref_846_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_889_load_0_req_0,ptr_deref_889_load_0_ack_0,ptr_deref_889_load_0_req_1,ptr_deref_889_load_0_ack_1,sl_one,"ptr_deref_889_load_0",false,ptr_deref_889_word_address_0,
    false,ptr_deref_889_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_932_load_0_req_0,ptr_deref_932_load_0_ack_0,ptr_deref_932_load_0_req_1,ptr_deref_932_load_0_ack_1,sl_one,"ptr_deref_932_load_0",false,ptr_deref_932_word_address_0,
    false,ptr_deref_932_data_0);
    -- shared load operator group (16) : ptr_deref_717_load_0 ptr_deref_674_load_0 ptr_deref_975_load_0 ptr_deref_760_load_0 ptr_deref_803_load_0 ptr_deref_846_load_0 ptr_deref_889_load_0 ptr_deref_932_load_0 
    LoadGroup16: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_717_load_0_req_0,
        ptr_deref_717_load_0_ack_0,
        ptr_deref_717_load_0_req_1,
        ptr_deref_717_load_0_ack_1,
        "ptr_deref_717_load_0",
        "memory_space_1" ,
        ptr_deref_717_data_0,
        ptr_deref_717_word_address_0,
        "ptr_deref_717_data_0",
        "ptr_deref_717_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_674_load_0_req_0,
        ptr_deref_674_load_0_ack_0,
        ptr_deref_674_load_0_req_1,
        ptr_deref_674_load_0_ack_1,
        "ptr_deref_674_load_0",
        "memory_space_1" ,
        ptr_deref_674_data_0,
        ptr_deref_674_word_address_0,
        "ptr_deref_674_data_0",
        "ptr_deref_674_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_975_load_0_req_0,
        ptr_deref_975_load_0_ack_0,
        ptr_deref_975_load_0_req_1,
        ptr_deref_975_load_0_ack_1,
        "ptr_deref_975_load_0",
        "memory_space_1" ,
        ptr_deref_975_data_0,
        ptr_deref_975_word_address_0,
        "ptr_deref_975_data_0",
        "ptr_deref_975_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_760_load_0_req_0,
        ptr_deref_760_load_0_ack_0,
        ptr_deref_760_load_0_req_1,
        ptr_deref_760_load_0_ack_1,
        "ptr_deref_760_load_0",
        "memory_space_1" ,
        ptr_deref_760_data_0,
        ptr_deref_760_word_address_0,
        "ptr_deref_760_data_0",
        "ptr_deref_760_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_803_load_0_req_0,
        ptr_deref_803_load_0_ack_0,
        ptr_deref_803_load_0_req_1,
        ptr_deref_803_load_0_ack_1,
        "ptr_deref_803_load_0",
        "memory_space_1" ,
        ptr_deref_803_data_0,
        ptr_deref_803_word_address_0,
        "ptr_deref_803_data_0",
        "ptr_deref_803_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_846_load_0_req_0,
        ptr_deref_846_load_0_ack_0,
        ptr_deref_846_load_0_req_1,
        ptr_deref_846_load_0_ack_1,
        "ptr_deref_846_load_0",
        "memory_space_1" ,
        ptr_deref_846_data_0,
        ptr_deref_846_word_address_0,
        "ptr_deref_846_data_0",
        "ptr_deref_846_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_889_load_0_req_0,
        ptr_deref_889_load_0_ack_0,
        ptr_deref_889_load_0_req_1,
        ptr_deref_889_load_0_ack_1,
        "ptr_deref_889_load_0",
        "memory_space_1" ,
        ptr_deref_889_data_0,
        ptr_deref_889_word_address_0,
        "ptr_deref_889_data_0",
        "ptr_deref_889_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_932_load_0_req_0,
        ptr_deref_932_load_0_ack_0,
        ptr_deref_932_load_0_req_1,
        ptr_deref_932_load_0_ack_1,
        "ptr_deref_932_load_0",
        "memory_space_1" ,
        ptr_deref_932_data_0,
        ptr_deref_932_word_address_0,
        "ptr_deref_932_data_0",
        "ptr_deref_932_word_address_0" -- 
      );
      reqL_unguarded(7) <= ptr_deref_717_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_674_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_975_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_760_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_803_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_846_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_889_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_932_load_0_req_0;
      ptr_deref_717_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_674_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_975_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_760_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_803_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_846_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_889_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_932_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_717_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_674_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_975_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_760_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_803_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_846_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_889_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_932_load_0_req_1;
      ptr_deref_717_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_674_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_975_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_760_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_803_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_846_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_889_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_932_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_717_word_address_0 & ptr_deref_674_word_address_0 & ptr_deref_975_word_address_0 & ptr_deref_760_word_address_0 & ptr_deref_803_word_address_0 & ptr_deref_846_word_address_0 & ptr_deref_889_word_address_0 & ptr_deref_932_word_address_0;
      ptr_deref_717_data_0 <= data_out(255 downto 224);
      ptr_deref_674_data_0 <= data_out(223 downto 192);
      ptr_deref_975_data_0 <= data_out(191 downto 160);
      ptr_deref_760_data_0 <= data_out(159 downto 128);
      ptr_deref_803_data_0 <= data_out(127 downto 96);
      ptr_deref_846_data_0 <= data_out(95 downto 64);
      ptr_deref_889_data_0 <= data_out(63 downto 32);
      ptr_deref_932_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 8,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 16
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_988_load_0_req_0,ptr_deref_988_load_0_ack_0,ptr_deref_988_load_0_req_1,ptr_deref_988_load_0_ack_1,sl_one,"ptr_deref_988_load_0",false,ptr_deref_988_word_address_0,
    false,ptr_deref_988_data_0);
    -- shared load operator group (17) : ptr_deref_988_load_0 
    LoadGroup17: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_988_load_0_req_0,
        ptr_deref_988_load_0_ack_0,
        ptr_deref_988_load_0_req_1,
        ptr_deref_988_load_0_ack_1,
        "ptr_deref_988_load_0",
        "memory_space_15" ,
        ptr_deref_988_data_0,
        ptr_deref_988_word_address_0,
        "ptr_deref_988_data_0",
        "ptr_deref_988_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_988_load_0_req_0;
      ptr_deref_988_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_988_load_0_req_1;
      ptr_deref_988_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_988_word_address_0;
      ptr_deref_988_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_15_lr_req(0),
          mack => memory_space_15_lr_ack(0),
          maddr => memory_space_15_lr_addr(0 downto 0),
          mtag => memory_space_15_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_15_lc_req(0),
          mack => memory_space_15_lc_ack(0),
          mdata => memory_space_15_lc_data(31 downto 0),
          mtag => memory_space_15_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 17
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1004_store_0_req_0,ptr_deref_1004_store_0_ack_0,ptr_deref_1004_store_0_req_1,ptr_deref_1004_store_0_ack_1,sl_one,"ptr_deref_1004_store_0",false,ptr_deref_1004_word_address_0 & ptr_deref_1004_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1025_store_0_req_0,ptr_deref_1025_store_0_ack_0,ptr_deref_1025_store_0_req_1,ptr_deref_1025_store_0_ack_1,sl_one,"ptr_deref_1025_store_0",false,ptr_deref_1025_word_address_0 & ptr_deref_1025_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1046_store_0_req_0,ptr_deref_1046_store_0_ack_0,ptr_deref_1046_store_0_req_1,ptr_deref_1046_store_0_ack_1,sl_one,"ptr_deref_1046_store_0",false,ptr_deref_1046_word_address_0 & ptr_deref_1046_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1130_store_0_req_0,ptr_deref_1130_store_0_ack_0,ptr_deref_1130_store_0_req_1,ptr_deref_1130_store_0_ack_1,sl_one,"ptr_deref_1130_store_0",false,ptr_deref_1130_word_address_0 & ptr_deref_1130_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1109_store_0_req_0,ptr_deref_1109_store_0_ack_0,ptr_deref_1109_store_0_req_1,ptr_deref_1109_store_0_ack_1,sl_one,"ptr_deref_1109_store_0",false,ptr_deref_1109_word_address_0 & ptr_deref_1109_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1151_store_0_req_0,ptr_deref_1151_store_0_ack_0,ptr_deref_1151_store_0_req_1,ptr_deref_1151_store_0_ack_1,sl_one,"ptr_deref_1151_store_0",false,ptr_deref_1151_word_address_0 & ptr_deref_1151_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1088_store_0_req_0,ptr_deref_1088_store_0_ack_0,ptr_deref_1088_store_0_req_1,ptr_deref_1088_store_0_ack_1,sl_one,"ptr_deref_1088_store_0",false,ptr_deref_1088_word_address_0 & ptr_deref_1088_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1067_store_0_req_0,ptr_deref_1067_store_0_ack_0,ptr_deref_1067_store_0_req_1,ptr_deref_1067_store_0_ack_1,sl_one,"ptr_deref_1067_store_0",false,ptr_deref_1067_word_address_0 & ptr_deref_1067_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1004_store_0_req_0,
      ptr_deref_1004_store_0_ack_0,
      ptr_deref_1004_store_0_req_1,
      ptr_deref_1004_store_0_ack_1,
      "ptr_deref_1004_store_0",
      "memory_space_2" ,
      ptr_deref_1004_data_0,
      ptr_deref_1004_word_address_0,
      "ptr_deref_1004_data_0",
      "ptr_deref_1004_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1025_store_0_req_0,
      ptr_deref_1025_store_0_ack_0,
      ptr_deref_1025_store_0_req_1,
      ptr_deref_1025_store_0_ack_1,
      "ptr_deref_1025_store_0",
      "memory_space_2" ,
      ptr_deref_1025_data_0,
      ptr_deref_1025_word_address_0,
      "ptr_deref_1025_data_0",
      "ptr_deref_1025_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1046_store_0_req_0,
      ptr_deref_1046_store_0_ack_0,
      ptr_deref_1046_store_0_req_1,
      ptr_deref_1046_store_0_ack_1,
      "ptr_deref_1046_store_0",
      "memory_space_2" ,
      ptr_deref_1046_data_0,
      ptr_deref_1046_word_address_0,
      "ptr_deref_1046_data_0",
      "ptr_deref_1046_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1130_store_0_req_0,
      ptr_deref_1130_store_0_ack_0,
      ptr_deref_1130_store_0_req_1,
      ptr_deref_1130_store_0_ack_1,
      "ptr_deref_1130_store_0",
      "memory_space_2" ,
      ptr_deref_1130_data_0,
      ptr_deref_1130_word_address_0,
      "ptr_deref_1130_data_0",
      "ptr_deref_1130_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1109_store_0_req_0,
      ptr_deref_1109_store_0_ack_0,
      ptr_deref_1109_store_0_req_1,
      ptr_deref_1109_store_0_ack_1,
      "ptr_deref_1109_store_0",
      "memory_space_2" ,
      ptr_deref_1109_data_0,
      ptr_deref_1109_word_address_0,
      "ptr_deref_1109_data_0",
      "ptr_deref_1109_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1151_store_0_req_0,
      ptr_deref_1151_store_0_ack_0,
      ptr_deref_1151_store_0_req_1,
      ptr_deref_1151_store_0_ack_1,
      "ptr_deref_1151_store_0",
      "memory_space_2" ,
      ptr_deref_1151_data_0,
      ptr_deref_1151_word_address_0,
      "ptr_deref_1151_data_0",
      "ptr_deref_1151_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1088_store_0_req_0,
      ptr_deref_1088_store_0_ack_0,
      ptr_deref_1088_store_0_req_1,
      ptr_deref_1088_store_0_ack_1,
      "ptr_deref_1088_store_0",
      "memory_space_2" ,
      ptr_deref_1088_data_0,
      ptr_deref_1088_word_address_0,
      "ptr_deref_1088_data_0",
      "ptr_deref_1088_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1067_store_0_req_0,
      ptr_deref_1067_store_0_ack_0,
      ptr_deref_1067_store_0_req_1,
      ptr_deref_1067_store_0_ack_1,
      "ptr_deref_1067_store_0",
      "memory_space_2" ,
      ptr_deref_1067_data_0,
      ptr_deref_1067_word_address_0,
      "ptr_deref_1067_data_0",
      "ptr_deref_1067_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_1004_store_0 ptr_deref_1025_store_0 ptr_deref_1046_store_0 ptr_deref_1130_store_0 ptr_deref_1109_store_0 ptr_deref_1151_store_0 ptr_deref_1088_store_0 ptr_deref_1067_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_1004_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_1025_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_1046_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_1130_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_1109_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_1151_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_1088_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1067_store_0_req_0;
      ptr_deref_1004_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_1025_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_1046_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_1130_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_1109_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_1151_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_1088_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1067_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_1004_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_1025_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_1046_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_1130_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_1109_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_1151_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_1088_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1067_store_0_req_1;
      ptr_deref_1004_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_1025_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_1046_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_1130_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_1109_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_1151_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_1088_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1067_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_1004_word_address_0 & ptr_deref_1025_word_address_0 & ptr_deref_1046_word_address_0 & ptr_deref_1130_word_address_0 & ptr_deref_1109_word_address_0 & ptr_deref_1151_word_address_0 & ptr_deref_1088_word_address_0 & ptr_deref_1067_word_address_0;
      data_in <= ptr_deref_1004_data_0 & ptr_deref_1025_data_0 & ptr_deref_1046_data_0 & ptr_deref_1130_data_0 & ptr_deref_1109_data_0 & ptr_deref_1151_data_0 & ptr_deref_1088_data_0 & ptr_deref_1067_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_459_store_0_req_0,ptr_deref_459_store_0_ack_0,ptr_deref_459_store_0_req_1,ptr_deref_459_store_0_ack_1,sl_one,"ptr_deref_459_store_0",false,ptr_deref_459_word_address_0 & ptr_deref_459_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_1175_store_0_req_0,ptr_deref_1175_store_0_ack_0,ptr_deref_1175_store_0_req_1,ptr_deref_1175_store_0_ack_1,sl_one,"ptr_deref_1175_store_0",false,ptr_deref_1175_word_address_0 & ptr_deref_1175_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_459_store_0_req_0,
      ptr_deref_459_store_0_ack_0,
      ptr_deref_459_store_0_req_1,
      ptr_deref_459_store_0_ack_1,
      "ptr_deref_459_store_0",
      "memory_space_7" ,
      ptr_deref_459_data_0,
      ptr_deref_459_word_address_0,
      "ptr_deref_459_data_0",
      "ptr_deref_459_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_1175_store_0_req_0,
      ptr_deref_1175_store_0_ack_0,
      ptr_deref_1175_store_0_req_1,
      ptr_deref_1175_store_0_ack_1,
      "ptr_deref_1175_store_0",
      "memory_space_7" ,
      ptr_deref_1175_data_0,
      ptr_deref_1175_word_address_0,
      "ptr_deref_1175_data_0",
      "ptr_deref_1175_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_459_store_0 ptr_deref_1175_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      -- 
    begin -- 
      reqL_unguarded(1) <= ptr_deref_459_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_1175_store_0_req_0;
      ptr_deref_459_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_1175_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= ptr_deref_459_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_1175_store_0_req_1;
      ptr_deref_459_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_1175_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 2) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_459_word_address_0 & ptr_deref_1175_word_address_0;
      data_in <= ptr_deref_459_data_0 & ptr_deref_1175_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 2,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(7 downto 0),
          mtag => memory_space_7_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_507_store_0_req_0,ptr_deref_507_store_0_ack_0,ptr_deref_507_store_0_req_1,ptr_deref_507_store_0_ack_1,sl_one,"ptr_deref_507_store_0",false,ptr_deref_507_word_address_0 & ptr_deref_507_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_507_store_0_req_0,
      ptr_deref_507_store_0_ack_0,
      ptr_deref_507_store_0_req_1,
      ptr_deref_507_store_0_ack_1,
      "ptr_deref_507_store_0",
      "memory_space_8" ,
      ptr_deref_507_data_0,
      ptr_deref_507_word_address_0,
      "ptr_deref_507_data_0",
      "ptr_deref_507_word_address_0" -- 
    );
    -- shared store operator group (2) : ptr_deref_507_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_507_store_0_req_0;
      ptr_deref_507_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_507_store_0_req_1;
      ptr_deref_507_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_507_word_address_0;
      data_in <= ptr_deref_507_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(7 downto 0),
          mtag => memory_space_8_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_529_store_0_req_0,ptr_deref_529_store_0_ack_0,ptr_deref_529_store_0_req_1,ptr_deref_529_store_0_ack_1,sl_one,"ptr_deref_529_store_0",false,ptr_deref_529_word_address_0 & ptr_deref_529_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_529_store_0_req_0,
      ptr_deref_529_store_0_ack_0,
      ptr_deref_529_store_0_req_1,
      ptr_deref_529_store_0_ack_1,
      "ptr_deref_529_store_0",
      "memory_space_9" ,
      ptr_deref_529_data_0,
      ptr_deref_529_word_address_0,
      "ptr_deref_529_data_0",
      "ptr_deref_529_word_address_0" -- 
    );
    -- shared store operator group (3) : ptr_deref_529_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_529_store_0_req_0;
      ptr_deref_529_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_529_store_0_req_1;
      ptr_deref_529_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_529_word_address_0;
      data_in <= ptr_deref_529_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(0 downto 0),
          mdata => memory_space_9_sr_data(7 downto 0),
          mtag => memory_space_9_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_551_store_0_req_0,ptr_deref_551_store_0_ack_0,ptr_deref_551_store_0_req_1,ptr_deref_551_store_0_ack_1,sl_one,"ptr_deref_551_store_0",false,ptr_deref_551_word_address_0 & ptr_deref_551_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_551_store_0_req_0,
      ptr_deref_551_store_0_ack_0,
      ptr_deref_551_store_0_req_1,
      ptr_deref_551_store_0_ack_1,
      "ptr_deref_551_store_0",
      "memory_space_10" ,
      ptr_deref_551_data_0,
      ptr_deref_551_word_address_0,
      "ptr_deref_551_data_0",
      "ptr_deref_551_word_address_0" -- 
    );
    -- shared store operator group (4) : ptr_deref_551_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_551_store_0_req_0;
      ptr_deref_551_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_551_store_0_req_1;
      ptr_deref_551_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_551_word_address_0;
      data_in <= ptr_deref_551_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_10_sr_req(0),
          mack => memory_space_10_sr_ack(0),
          maddr => memory_space_10_sr_addr(0 downto 0),
          mdata => memory_space_10_sr_data(7 downto 0),
          mtag => memory_space_10_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_10_sc_req(0),
          mack => memory_space_10_sc_ack(0),
          mtag => memory_space_10_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_573_store_0_req_0,ptr_deref_573_store_0_ack_0,ptr_deref_573_store_0_req_1,ptr_deref_573_store_0_ack_1,sl_one,"ptr_deref_573_store_0",false,ptr_deref_573_word_address_0 & ptr_deref_573_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_573_store_0_req_0,
      ptr_deref_573_store_0_ack_0,
      ptr_deref_573_store_0_req_1,
      ptr_deref_573_store_0_ack_1,
      "ptr_deref_573_store_0",
      "memory_space_11" ,
      ptr_deref_573_data_0,
      ptr_deref_573_word_address_0,
      "ptr_deref_573_data_0",
      "ptr_deref_573_word_address_0" -- 
    );
    -- shared store operator group (5) : ptr_deref_573_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_573_store_0_req_0;
      ptr_deref_573_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_573_store_0_req_1;
      ptr_deref_573_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_573_word_address_0;
      data_in <= ptr_deref_573_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_11_sr_req(0),
          mack => memory_space_11_sr_ack(0),
          maddr => memory_space_11_sr_addr(0 downto 0),
          mdata => memory_space_11_sr_data(7 downto 0),
          mtag => memory_space_11_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_11_sc_req(0),
          mack => memory_space_11_sc_ack(0),
          mtag => memory_space_11_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_595_store_0_req_0,ptr_deref_595_store_0_ack_0,ptr_deref_595_store_0_req_1,ptr_deref_595_store_0_ack_1,sl_one,"ptr_deref_595_store_0",false,ptr_deref_595_word_address_0 & ptr_deref_595_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_595_store_0_req_0,
      ptr_deref_595_store_0_ack_0,
      ptr_deref_595_store_0_req_1,
      ptr_deref_595_store_0_ack_1,
      "ptr_deref_595_store_0",
      "memory_space_12" ,
      ptr_deref_595_data_0,
      ptr_deref_595_word_address_0,
      "ptr_deref_595_data_0",
      "ptr_deref_595_word_address_0" -- 
    );
    -- shared store operator group (6) : ptr_deref_595_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_595_store_0_req_0;
      ptr_deref_595_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_595_store_0_req_1;
      ptr_deref_595_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_595_word_address_0;
      data_in <= ptr_deref_595_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_12_sr_req(0),
          mack => memory_space_12_sr_ack(0),
          maddr => memory_space_12_sr_addr(0 downto 0),
          mdata => memory_space_12_sr_data(7 downto 0),
          mtag => memory_space_12_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_12_sc_req(0),
          mack => memory_space_12_sc_ack(0),
          mtag => memory_space_12_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_617_store_0_req_0,ptr_deref_617_store_0_ack_0,ptr_deref_617_store_0_req_1,ptr_deref_617_store_0_ack_1,sl_one,"ptr_deref_617_store_0",false,ptr_deref_617_word_address_0 & ptr_deref_617_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_617_store_0_req_0,
      ptr_deref_617_store_0_ack_0,
      ptr_deref_617_store_0_req_1,
      ptr_deref_617_store_0_ack_1,
      "ptr_deref_617_store_0",
      "memory_space_13" ,
      ptr_deref_617_data_0,
      ptr_deref_617_word_address_0,
      "ptr_deref_617_data_0",
      "ptr_deref_617_word_address_0" -- 
    );
    -- shared store operator group (7) : ptr_deref_617_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_617_store_0_req_0;
      ptr_deref_617_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_617_store_0_req_1;
      ptr_deref_617_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_617_word_address_0;
      data_in <= ptr_deref_617_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_13_sr_req(0),
          mack => memory_space_13_sr_ack(0),
          maddr => memory_space_13_sr_addr(0 downto 0),
          mdata => memory_space_13_sr_data(7 downto 0),
          mtag => memory_space_13_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_13_sc_req(0),
          mack => memory_space_13_sc_ack(0),
          mtag => memory_space_13_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_639_store_0_req_0,ptr_deref_639_store_0_ack_0,ptr_deref_639_store_0_req_1,ptr_deref_639_store_0_ack_1,sl_one,"ptr_deref_639_store_0",false,ptr_deref_639_word_address_0 & ptr_deref_639_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_639_store_0_req_0,
      ptr_deref_639_store_0_ack_0,
      ptr_deref_639_store_0_req_1,
      ptr_deref_639_store_0_ack_1,
      "ptr_deref_639_store_0",
      "memory_space_14" ,
      ptr_deref_639_data_0,
      ptr_deref_639_word_address_0,
      "ptr_deref_639_data_0",
      "ptr_deref_639_word_address_0" -- 
    );
    -- shared store operator group (8) : ptr_deref_639_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_639_store_0_req_0;
      ptr_deref_639_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_639_store_0_req_1;
      ptr_deref_639_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_639_word_address_0;
      data_in <= ptr_deref_639_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_14_sr_req(0),
          mack => memory_space_14_sr_ack(0),
          maddr => memory_space_14_sr_addr(0 downto 0),
          mdata => memory_space_14_sr_data(7 downto 0),
          mtag => memory_space_14_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_14_sc_req(0),
          mack => memory_space_14_sc_ack(0),
          mtag => memory_space_14_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_682_store_0_req_0,ptr_deref_682_store_0_ack_0,ptr_deref_682_store_0_req_1,ptr_deref_682_store_0_ack_1,sl_one,"ptr_deref_682_store_0",false,ptr_deref_682_word_address_0 & ptr_deref_682_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_682_store_0_req_0,
      ptr_deref_682_store_0_ack_0,
      ptr_deref_682_store_0_req_1,
      ptr_deref_682_store_0_ack_1,
      "ptr_deref_682_store_0",
      "memory_space_15" ,
      ptr_deref_682_data_0,
      ptr_deref_682_word_address_0,
      "ptr_deref_682_data_0",
      "ptr_deref_682_word_address_0" -- 
    );
    -- shared store operator group (9) : ptr_deref_682_store_0 
    StoreGroup9: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_682_store_0_req_0;
      ptr_deref_682_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_682_store_0_req_1;
      ptr_deref_682_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_682_word_address_0;
      data_in <= ptr_deref_682_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_15_sr_req(0),
          mack => memory_space_15_sr_ack(0),
          maddr => memory_space_15_sr_addr(0 downto 0),
          mdata => memory_space_15_sr_data(31 downto 0),
          mtag => memory_space_15_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_15_sc_req(0),
          mack => memory_space_15_sc_ack(0),
          mtag => memory_space_15_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 9
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_725_store_0_req_0,ptr_deref_725_store_0_ack_0,ptr_deref_725_store_0_req_1,ptr_deref_725_store_0_ack_1,sl_one,"ptr_deref_725_store_0",false,ptr_deref_725_word_address_0 & ptr_deref_725_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_725_store_0_req_0,
      ptr_deref_725_store_0_ack_0,
      ptr_deref_725_store_0_req_1,
      ptr_deref_725_store_0_ack_1,
      "ptr_deref_725_store_0",
      "memory_space_16" ,
      ptr_deref_725_data_0,
      ptr_deref_725_word_address_0,
      "ptr_deref_725_data_0",
      "ptr_deref_725_word_address_0" -- 
    );
    -- shared store operator group (10) : ptr_deref_725_store_0 
    StoreGroup10: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_725_store_0_req_0;
      ptr_deref_725_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_725_store_0_req_1;
      ptr_deref_725_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_725_word_address_0;
      data_in <= ptr_deref_725_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_16_sr_req(0),
          mack => memory_space_16_sr_ack(0),
          maddr => memory_space_16_sr_addr(0 downto 0),
          mdata => memory_space_16_sr_data(31 downto 0),
          mtag => memory_space_16_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_16_sc_req(0),
          mack => memory_space_16_sc_ack(0),
          mtag => memory_space_16_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 10
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_768_store_0_req_0,ptr_deref_768_store_0_ack_0,ptr_deref_768_store_0_req_1,ptr_deref_768_store_0_ack_1,sl_one,"ptr_deref_768_store_0",false,ptr_deref_768_word_address_0 & ptr_deref_768_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_768_store_0_req_0,
      ptr_deref_768_store_0_ack_0,
      ptr_deref_768_store_0_req_1,
      ptr_deref_768_store_0_ack_1,
      "ptr_deref_768_store_0",
      "memory_space_17" ,
      ptr_deref_768_data_0,
      ptr_deref_768_word_address_0,
      "ptr_deref_768_data_0",
      "ptr_deref_768_word_address_0" -- 
    );
    -- shared store operator group (11) : ptr_deref_768_store_0 
    StoreGroup11: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_768_store_0_req_0;
      ptr_deref_768_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_768_store_0_req_1;
      ptr_deref_768_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_768_word_address_0;
      data_in <= ptr_deref_768_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_17_sr_req(0),
          mack => memory_space_17_sr_ack(0),
          maddr => memory_space_17_sr_addr(0 downto 0),
          mdata => memory_space_17_sr_data(31 downto 0),
          mtag => memory_space_17_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_17_sc_req(0),
          mack => memory_space_17_sc_ack(0),
          mtag => memory_space_17_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 11
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_811_store_0_req_0,ptr_deref_811_store_0_ack_0,ptr_deref_811_store_0_req_1,ptr_deref_811_store_0_ack_1,sl_one,"ptr_deref_811_store_0",false,ptr_deref_811_word_address_0 & ptr_deref_811_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_811_store_0_req_0,
      ptr_deref_811_store_0_ack_0,
      ptr_deref_811_store_0_req_1,
      ptr_deref_811_store_0_ack_1,
      "ptr_deref_811_store_0",
      "memory_space_18" ,
      ptr_deref_811_data_0,
      ptr_deref_811_word_address_0,
      "ptr_deref_811_data_0",
      "ptr_deref_811_word_address_0" -- 
    );
    -- shared store operator group (12) : ptr_deref_811_store_0 
    StoreGroup12: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_811_store_0_req_0;
      ptr_deref_811_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_811_store_0_req_1;
      ptr_deref_811_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_811_word_address_0;
      data_in <= ptr_deref_811_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_18_sr_req(0),
          mack => memory_space_18_sr_ack(0),
          maddr => memory_space_18_sr_addr(0 downto 0),
          mdata => memory_space_18_sr_data(31 downto 0),
          mtag => memory_space_18_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_18_sc_req(0),
          mack => memory_space_18_sc_ack(0),
          mtag => memory_space_18_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 12
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_854_store_0_req_0,ptr_deref_854_store_0_ack_0,ptr_deref_854_store_0_req_1,ptr_deref_854_store_0_ack_1,sl_one,"ptr_deref_854_store_0",false,ptr_deref_854_word_address_0 & ptr_deref_854_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_854_store_0_req_0,
      ptr_deref_854_store_0_ack_0,
      ptr_deref_854_store_0_req_1,
      ptr_deref_854_store_0_ack_1,
      "ptr_deref_854_store_0",
      "memory_space_19" ,
      ptr_deref_854_data_0,
      ptr_deref_854_word_address_0,
      "ptr_deref_854_data_0",
      "ptr_deref_854_word_address_0" -- 
    );
    -- shared store operator group (13) : ptr_deref_854_store_0 
    StoreGroup13: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_854_store_0_req_0;
      ptr_deref_854_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_854_store_0_req_1;
      ptr_deref_854_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_854_word_address_0;
      data_in <= ptr_deref_854_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_19_sr_req(0),
          mack => memory_space_19_sr_ack(0),
          maddr => memory_space_19_sr_addr(0 downto 0),
          mdata => memory_space_19_sr_data(31 downto 0),
          mtag => memory_space_19_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_19_sc_req(0),
          mack => memory_space_19_sc_ack(0),
          mtag => memory_space_19_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 13
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_897_store_0_req_0,ptr_deref_897_store_0_ack_0,ptr_deref_897_store_0_req_1,ptr_deref_897_store_0_ack_1,sl_one,"ptr_deref_897_store_0",false,ptr_deref_897_word_address_0 & ptr_deref_897_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_897_store_0_req_0,
      ptr_deref_897_store_0_ack_0,
      ptr_deref_897_store_0_req_1,
      ptr_deref_897_store_0_ack_1,
      "ptr_deref_897_store_0",
      "memory_space_20" ,
      ptr_deref_897_data_0,
      ptr_deref_897_word_address_0,
      "ptr_deref_897_data_0",
      "ptr_deref_897_word_address_0" -- 
    );
    -- shared store operator group (14) : ptr_deref_897_store_0 
    StoreGroup14: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_897_store_0_req_0;
      ptr_deref_897_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_897_store_0_req_1;
      ptr_deref_897_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_897_word_address_0;
      data_in <= ptr_deref_897_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_20_sr_req(0),
          mack => memory_space_20_sr_ack(0),
          maddr => memory_space_20_sr_addr(0 downto 0),
          mdata => memory_space_20_sr_data(31 downto 0),
          mtag => memory_space_20_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_20_sc_req(0),
          mack => memory_space_20_sc_ack(0),
          mtag => memory_space_20_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 14
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_940_store_0_req_0,ptr_deref_940_store_0_ack_0,ptr_deref_940_store_0_req_1,ptr_deref_940_store_0_ack_1,sl_one,"ptr_deref_940_store_0",false,ptr_deref_940_word_address_0 & ptr_deref_940_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_940_store_0_req_0,
      ptr_deref_940_store_0_ack_0,
      ptr_deref_940_store_0_req_1,
      ptr_deref_940_store_0_ack_1,
      "ptr_deref_940_store_0",
      "memory_space_21" ,
      ptr_deref_940_data_0,
      ptr_deref_940_word_address_0,
      "ptr_deref_940_data_0",
      "ptr_deref_940_word_address_0" -- 
    );
    -- shared store operator group (15) : ptr_deref_940_store_0 
    StoreGroup15: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_940_store_0_req_0;
      ptr_deref_940_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_940_store_0_req_1;
      ptr_deref_940_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_940_word_address_0;
      data_in <= ptr_deref_940_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_21_sr_req(0),
          mack => memory_space_21_sr_ack(0),
          maddr => memory_space_21_sr_addr(0 downto 0),
          mdata => memory_space_21_sr_data(31 downto 0),
          mtag => memory_space_21_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_21_sc_req(0),
          mack => memory_space_21_sc_ack(0),
          mtag => memory_space_21_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 15
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_983_store_0_req_0,ptr_deref_983_store_0_ack_0,ptr_deref_983_store_0_req_1,ptr_deref_983_store_0_ack_1,sl_one,"ptr_deref_983_store_0",false,ptr_deref_983_word_address_0 & ptr_deref_983_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_983_store_0_req_0,
      ptr_deref_983_store_0_ack_0,
      ptr_deref_983_store_0_req_1,
      ptr_deref_983_store_0_ack_1,
      "ptr_deref_983_store_0",
      "memory_space_22" ,
      ptr_deref_983_data_0,
      ptr_deref_983_word_address_0,
      "ptr_deref_983_data_0",
      "ptr_deref_983_word_address_0" -- 
    );
    -- shared store operator group (16) : ptr_deref_983_store_0 
    StoreGroup16: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_983_store_0_req_0;
      ptr_deref_983_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_983_store_0_req_1;
      ptr_deref_983_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_983_word_address_0;
      data_in <= ptr_deref_983_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_22_sr_req(0),
          mack => memory_space_22_sr_ack(0),
          maddr => memory_space_22_sr_addr(0 downto 0),
          mdata => memory_space_22_sr_data(31 downto 0),
          mtag => memory_space_22_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_22_sc_req(0),
          mack => memory_space_22_sc_ack(0),
          mtag => memory_space_22_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 16
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_10: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_10_lr_addr,
      lr_req_in => memory_space_10_lr_req,
      lr_ack_out => memory_space_10_lr_ack,
      lr_tag_in => memory_space_10_lr_tag,
      lc_req_in => memory_space_10_lc_req,
      lc_ack_out => memory_space_10_lc_ack,
      lc_data_out => memory_space_10_lc_data,
      lc_tag_out => memory_space_10_lc_tag,
      sr_addr_in => memory_space_10_sr_addr,
      sr_data_in => memory_space_10_sr_data,
      sr_req_in => memory_space_10_sr_req,
      sr_ack_out => memory_space_10_sr_ack,
      sr_tag_in => memory_space_10_sr_tag,
      sc_req_in=> memory_space_10_sc_req,
      sc_ack_out => memory_space_10_sc_ack,
      sc_tag_out => memory_space_10_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_11: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_11_lr_addr,
      lr_req_in => memory_space_11_lr_req,
      lr_ack_out => memory_space_11_lr_ack,
      lr_tag_in => memory_space_11_lr_tag,
      lc_req_in => memory_space_11_lc_req,
      lc_ack_out => memory_space_11_lc_ack,
      lc_data_out => memory_space_11_lc_data,
      lc_tag_out => memory_space_11_lc_tag,
      sr_addr_in => memory_space_11_sr_addr,
      sr_data_in => memory_space_11_sr_data,
      sr_req_in => memory_space_11_sr_req,
      sr_ack_out => memory_space_11_sr_ack,
      sr_tag_in => memory_space_11_sr_tag,
      sc_req_in=> memory_space_11_sc_req,
      sc_ack_out => memory_space_11_sc_ack,
      sc_tag_out => memory_space_11_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_12: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_12_lr_addr,
      lr_req_in => memory_space_12_lr_req,
      lr_ack_out => memory_space_12_lr_ack,
      lr_tag_in => memory_space_12_lr_tag,
      lc_req_in => memory_space_12_lc_req,
      lc_ack_out => memory_space_12_lc_ack,
      lc_data_out => memory_space_12_lc_data,
      lc_tag_out => memory_space_12_lc_tag,
      sr_addr_in => memory_space_12_sr_addr,
      sr_data_in => memory_space_12_sr_data,
      sr_req_in => memory_space_12_sr_req,
      sr_ack_out => memory_space_12_sr_ack,
      sr_tag_in => memory_space_12_sr_tag,
      sc_req_in=> memory_space_12_sc_req,
      sc_ack_out => memory_space_12_sc_ack,
      sc_tag_out => memory_space_12_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_13: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_13_lr_addr,
      lr_req_in => memory_space_13_lr_req,
      lr_ack_out => memory_space_13_lr_ack,
      lr_tag_in => memory_space_13_lr_tag,
      lc_req_in => memory_space_13_lc_req,
      lc_ack_out => memory_space_13_lc_ack,
      lc_data_out => memory_space_13_lc_data,
      lc_tag_out => memory_space_13_lc_tag,
      sr_addr_in => memory_space_13_sr_addr,
      sr_data_in => memory_space_13_sr_data,
      sr_req_in => memory_space_13_sr_req,
      sr_ack_out => memory_space_13_sr_ack,
      sr_tag_in => memory_space_13_sr_tag,
      sc_req_in=> memory_space_13_sc_req,
      sc_ack_out => memory_space_13_sc_ack,
      sc_tag_out => memory_space_13_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_14: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_14_lr_addr,
      lr_req_in => memory_space_14_lr_req,
      lr_ack_out => memory_space_14_lr_ack,
      lr_tag_in => memory_space_14_lr_tag,
      lc_req_in => memory_space_14_lc_req,
      lc_ack_out => memory_space_14_lc_ack,
      lc_data_out => memory_space_14_lc_data,
      lc_tag_out => memory_space_14_lc_tag,
      sr_addr_in => memory_space_14_sr_addr,
      sr_data_in => memory_space_14_sr_data,
      sr_req_in => memory_space_14_sr_req,
      sr_ack_out => memory_space_14_sr_ack,
      sr_tag_in => memory_space_14_sr_tag,
      sc_req_in=> memory_space_14_sc_req,
      sc_ack_out => memory_space_14_sc_ack,
      sc_tag_out => memory_space_14_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_15: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_15_lr_addr,
      lr_req_in => memory_space_15_lr_req,
      lr_ack_out => memory_space_15_lr_ack,
      lr_tag_in => memory_space_15_lr_tag,
      lc_req_in => memory_space_15_lc_req,
      lc_ack_out => memory_space_15_lc_ack,
      lc_data_out => memory_space_15_lc_data,
      lc_tag_out => memory_space_15_lc_tag,
      sr_addr_in => memory_space_15_sr_addr,
      sr_data_in => memory_space_15_sr_data,
      sr_req_in => memory_space_15_sr_req,
      sr_ack_out => memory_space_15_sr_ack,
      sr_tag_in => memory_space_15_sr_tag,
      sc_req_in=> memory_space_15_sc_req,
      sc_ack_out => memory_space_15_sc_ack,
      sc_tag_out => memory_space_15_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_16: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_16_lr_addr,
      lr_req_in => memory_space_16_lr_req,
      lr_ack_out => memory_space_16_lr_ack,
      lr_tag_in => memory_space_16_lr_tag,
      lc_req_in => memory_space_16_lc_req,
      lc_ack_out => memory_space_16_lc_ack,
      lc_data_out => memory_space_16_lc_data,
      lc_tag_out => memory_space_16_lc_tag,
      sr_addr_in => memory_space_16_sr_addr,
      sr_data_in => memory_space_16_sr_data,
      sr_req_in => memory_space_16_sr_req,
      sr_ack_out => memory_space_16_sr_ack,
      sr_tag_in => memory_space_16_sr_tag,
      sc_req_in=> memory_space_16_sc_req,
      sc_ack_out => memory_space_16_sc_ack,
      sc_tag_out => memory_space_16_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_17: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_17_lr_addr,
      lr_req_in => memory_space_17_lr_req,
      lr_ack_out => memory_space_17_lr_ack,
      lr_tag_in => memory_space_17_lr_tag,
      lc_req_in => memory_space_17_lc_req,
      lc_ack_out => memory_space_17_lc_ack,
      lc_data_out => memory_space_17_lc_data,
      lc_tag_out => memory_space_17_lc_tag,
      sr_addr_in => memory_space_17_sr_addr,
      sr_data_in => memory_space_17_sr_data,
      sr_req_in => memory_space_17_sr_req,
      sr_ack_out => memory_space_17_sr_ack,
      sr_tag_in => memory_space_17_sr_tag,
      sc_req_in=> memory_space_17_sc_req,
      sc_ack_out => memory_space_17_sc_ack,
      sc_tag_out => memory_space_17_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_18: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_18_lr_addr,
      lr_req_in => memory_space_18_lr_req,
      lr_ack_out => memory_space_18_lr_ack,
      lr_tag_in => memory_space_18_lr_tag,
      lc_req_in => memory_space_18_lc_req,
      lc_ack_out => memory_space_18_lc_ack,
      lc_data_out => memory_space_18_lc_data,
      lc_tag_out => memory_space_18_lc_tag,
      sr_addr_in => memory_space_18_sr_addr,
      sr_data_in => memory_space_18_sr_data,
      sr_req_in => memory_space_18_sr_req,
      sr_ack_out => memory_space_18_sr_ack,
      sr_tag_in => memory_space_18_sr_tag,
      sc_req_in=> memory_space_18_sc_req,
      sc_ack_out => memory_space_18_sc_ack,
      sc_tag_out => memory_space_18_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_19: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_19_lr_addr,
      lr_req_in => memory_space_19_lr_req,
      lr_ack_out => memory_space_19_lr_ack,
      lr_tag_in => memory_space_19_lr_tag,
      lc_req_in => memory_space_19_lc_req,
      lc_ack_out => memory_space_19_lc_ack,
      lc_data_out => memory_space_19_lc_data,
      lc_tag_out => memory_space_19_lc_tag,
      sr_addr_in => memory_space_19_sr_addr,
      sr_data_in => memory_space_19_sr_data,
      sr_req_in => memory_space_19_sr_req,
      sr_ack_out => memory_space_19_sr_ack,
      sr_tag_in => memory_space_19_sr_tag,
      sc_req_in=> memory_space_19_sc_req,
      sc_ack_out => memory_space_19_sc_ack,
      sc_tag_out => memory_space_19_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_20: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_20_lr_addr,
      lr_req_in => memory_space_20_lr_req,
      lr_ack_out => memory_space_20_lr_ack,
      lr_tag_in => memory_space_20_lr_tag,
      lc_req_in => memory_space_20_lc_req,
      lc_ack_out => memory_space_20_lc_ack,
      lc_data_out => memory_space_20_lc_data,
      lc_tag_out => memory_space_20_lc_tag,
      sr_addr_in => memory_space_20_sr_addr,
      sr_data_in => memory_space_20_sr_data,
      sr_req_in => memory_space_20_sr_req,
      sr_ack_out => memory_space_20_sr_ack,
      sr_tag_in => memory_space_20_sr_tag,
      sc_req_in=> memory_space_20_sc_req,
      sc_ack_out => memory_space_20_sc_ack,
      sc_tag_out => memory_space_20_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_21: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_21_lr_addr,
      lr_req_in => memory_space_21_lr_req,
      lr_ack_out => memory_space_21_lr_ack,
      lr_tag_in => memory_space_21_lr_tag,
      lc_req_in => memory_space_21_lc_req,
      lc_ack_out => memory_space_21_lc_ack,
      lc_data_out => memory_space_21_lc_data,
      lc_tag_out => memory_space_21_lc_tag,
      sr_addr_in => memory_space_21_sr_addr,
      sr_data_in => memory_space_21_sr_data,
      sr_req_in => memory_space_21_sr_req,
      sr_ack_out => memory_space_21_sr_ack,
      sr_tag_in => memory_space_21_sr_tag,
      sc_req_in=> memory_space_21_sc_req,
      sc_ack_out => memory_space_21_sc_ack,
      sc_tag_out => memory_space_21_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_22: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_22_lr_addr,
      lr_req_in => memory_space_22_lr_req,
      lr_ack_out => memory_space_22_lr_ack,
      lr_tag_in => memory_space_22_lr_tag,
      lc_req_in => memory_space_22_lc_req,
      lc_ack_out => memory_space_22_lc_ack,
      lc_data_out => memory_space_22_lc_data,
      lc_tag_out => memory_space_22_lc_tag,
      sr_addr_in => memory_space_22_sr_addr,
      sr_data_in => memory_space_22_sr_data,
      sr_req_in => memory_space_22_sr_req,
      sr_ack_out => memory_space_22_sr_ack,
      sr_tag_in => memory_space_22_sr_tag,
      sc_req_in=> memory_space_22_sc_req,
      sc_ack_out => memory_space_22_sc_ack,
      sc_tag_out => memory_space_22_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 8,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module getData
  component getData is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(3 downto 0);
      in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module getData
  signal getData_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getData_tag_out   : std_logic_vector(1 downto 0);
  signal getData_start_req : std_logic;
  signal getData_start_ack : std_logic;
  signal getData_fin_req   : std_logic;
  signal getData_fin_ack : std_logic;
  -- caller side aggregated signals for module getData
  signal getData_call_reqs: std_logic_vector(0 downto 0);
  signal getData_call_acks: std_logic_vector(0 downto 0);
  signal getData_return_reqs: std_logic_vector(0 downto 0);
  signal getData_return_acks: std_logic_vector(0 downto 0);
  signal getData_call_tag: std_logic_vector(0 downto 0);
  signal getData_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module sendResult
  component sendResult is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      out_data_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module sendResult
  signal sendResult_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal sendResult_tag_out   : std_logic_vector(1 downto 0);
  signal sendResult_start_req : std_logic;
  signal sendResult_start_ack : std_logic;
  signal sendResult_fin_req   : std_logic;
  signal sendResult_fin_ack : std_logic;
  -- caller side aggregated signals for module sendResult
  signal sendResult_call_reqs: std_logic_vector(0 downto 0);
  signal sendResult_call_acks: std_logic_vector(0 downto 0);
  signal sendResult_return_reqs: std_logic_vector(0 downto 0);
  signal sendResult_return_acks: std_logic_vector(0 downto 0);
  signal sendResult_call_tag: std_logic_vector(0 downto 0);
  signal sendResult_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module vectorSum
  component vectorSum is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      x_vectorSum_x_call_reqs : out  std_logic_vector(0 downto 0);
      x_vectorSum_x_call_acks : in   std_logic_vector(0 downto 0);
      x_vectorSum_x_call_tag  :  out  std_logic_vector(0 downto 0);
      x_vectorSum_x_return_reqs : out  std_logic_vector(0 downto 0);
      x_vectorSum_x_return_acks : in   std_logic_vector(0 downto 0);
      x_vectorSum_x_return_tag :  in   std_logic_vector(0 downto 0);
      getData_call_reqs : out  std_logic_vector(0 downto 0);
      getData_call_acks : in   std_logic_vector(0 downto 0);
      getData_call_tag  :  out  std_logic_vector(0 downto 0);
      getData_return_reqs : out  std_logic_vector(0 downto 0);
      getData_return_acks : in   std_logic_vector(0 downto 0);
      getData_return_tag :  in   std_logic_vector(0 downto 0);
      sendResult_call_reqs : out  std_logic_vector(0 downto 0);
      sendResult_call_acks : in   std_logic_vector(0 downto 0);
      sendResult_call_tag  :  out  std_logic_vector(0 downto 0);
      sendResult_return_reqs : out  std_logic_vector(0 downto 0);
      sendResult_return_acks : in   std_logic_vector(0 downto 0);
      sendResult_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module vectorSum
  signal vectorSum_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal vectorSum_tag_out   : std_logic_vector(1 downto 0);
  signal vectorSum_start_req : std_logic;
  signal vectorSum_start_ack : std_logic;
  signal vectorSum_fin_req   : std_logic;
  signal vectorSum_fin_ack : std_logic;
  -- declarations related to module x_vectorSum_x
  component x_vectorSum_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module x_vectorSum_x
  signal x_vectorSum_x_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal x_vectorSum_x_tag_out   : std_logic_vector(1 downto 0);
  signal x_vectorSum_x_start_req : std_logic;
  signal x_vectorSum_x_start_ack : std_logic;
  signal x_vectorSum_x_fin_req   : std_logic;
  signal x_vectorSum_x_fin_ack : std_logic;
  -- caller side aggregated signals for module x_vectorSum_x
  signal x_vectorSum_x_call_reqs: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_call_acks: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_reqs: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_acks: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_call_tag: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_pipe
  signal in_data_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_pipe
  signal out_data_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module getData
  -- call arbiter for module getData
  getData_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getData_call_reqs,
      call_acks => getData_call_acks,
      return_reqs => getData_return_reqs,
      return_acks => getData_return_acks,
      call_tag  => getData_call_tag,
      return_tag  => getData_return_tag,
      call_mtag => getData_tag_in,
      return_mtag => getData_tag_out,
      call_mreq => getData_start_req,
      call_mack => getData_start_ack,
      return_mreq => getData_fin_req,
      return_mack => getData_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  getData_instance:getData-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => getData_start_req,
      start_ack => getData_start_ack,
      fin_req => getData_fin_req,
      fin_ack => getData_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(6 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(6 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      in_data_pipe_pipe_read_req => in_data_pipe_pipe_read_req(0 downto 0),
      in_data_pipe_pipe_read_ack => in_data_pipe_pipe_read_ack(0 downto 0),
      in_data_pipe_pipe_read_data => in_data_pipe_pipe_read_data(31 downto 0),
      tag_in => getData_tag_in,
      tag_out => getData_tag_out-- 
    ); -- 
  -- module sendResult
  -- call arbiter for module sendResult
  sendResult_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => sendResult_call_reqs,
      call_acks => sendResult_call_acks,
      return_reqs => sendResult_return_reqs,
      return_acks => sendResult_return_acks,
      call_tag  => sendResult_call_tag,
      return_tag  => sendResult_return_tag,
      call_mtag => sendResult_tag_in,
      return_mtag => sendResult_tag_out,
      call_mreq => sendResult_start_req,
      call_mack => sendResult_start_ack,
      return_mreq => sendResult_fin_req,
      return_mack => sendResult_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  sendResult_instance:sendResult-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => sendResult_start_req,
      start_ack => sendResult_start_ack,
      fin_req => sendResult_fin_req,
      fin_ack => sendResult_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(6 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      out_data_pipe_pipe_write_req => out_data_pipe_pipe_write_req(0 downto 0),
      out_data_pipe_pipe_write_ack => out_data_pipe_pipe_write_ack(0 downto 0),
      out_data_pipe_pipe_write_data => out_data_pipe_pipe_write_data(31 downto 0),
      tag_in => sendResult_tag_in,
      tag_out => sendResult_tag_out-- 
    ); -- 
  -- module vectorSum
  vectorSum_instance:vectorSum-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => vectorSum_start_req,
      start_ack => vectorSum_start_ack,
      fin_req => vectorSum_fin_req,
      fin_ack => vectorSum_fin_ack,
      clk => clk,
      reset => reset,
      getData_call_reqs => getData_call_reqs(0 downto 0),
      getData_call_acks => getData_call_acks(0 downto 0),
      getData_call_tag => getData_call_tag(0 downto 0),
      getData_return_reqs => getData_return_reqs(0 downto 0),
      getData_return_acks => getData_return_acks(0 downto 0),
      getData_return_tag => getData_return_tag(0 downto 0),
      sendResult_call_reqs => sendResult_call_reqs(0 downto 0),
      sendResult_call_acks => sendResult_call_acks(0 downto 0),
      sendResult_call_tag => sendResult_call_tag(0 downto 0),
      sendResult_return_reqs => sendResult_return_reqs(0 downto 0),
      sendResult_return_acks => sendResult_return_acks(0 downto 0),
      sendResult_return_tag => sendResult_return_tag(0 downto 0),
      x_vectorSum_x_call_reqs => x_vectorSum_x_call_reqs(0 downto 0),
      x_vectorSum_x_call_acks => x_vectorSum_x_call_acks(0 downto 0),
      x_vectorSum_x_call_tag => x_vectorSum_x_call_tag(0 downto 0),
      x_vectorSum_x_return_reqs => x_vectorSum_x_return_reqs(0 downto 0),
      x_vectorSum_x_return_acks => x_vectorSum_x_return_acks(0 downto 0),
      x_vectorSum_x_return_tag => x_vectorSum_x_return_tag(0 downto 0),
      tag_in => vectorSum_tag_in,
      tag_out => vectorSum_tag_out-- 
    ); -- 
  -- module will be run forever 
  vectorSum_tag_in <= (others => '0');
  vectorSum_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => vectorSum_start_req, start_ack => vectorSum_start_ack,  fin_req => vectorSum_fin_req,  fin_ack => vectorSum_fin_ack);
  -- module x_vectorSum_x
  -- call arbiter for module x_vectorSum_x
  x_vectorSum_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => x_vectorSum_x_call_reqs,
      call_acks => x_vectorSum_x_call_acks,
      return_reqs => x_vectorSum_x_return_reqs,
      return_acks => x_vectorSum_x_return_acks,
      call_tag  => x_vectorSum_x_call_tag,
      return_tag  => x_vectorSum_x_return_tag,
      call_mtag => x_vectorSum_x_tag_in,
      return_mtag => x_vectorSum_x_tag_out,
      call_mreq => x_vectorSum_x_start_req,
      call_mack => x_vectorSum_x_start_ack,
      return_mreq => x_vectorSum_x_fin_req,
      return_mack => x_vectorSum_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  x_vectorSum_x_instance:x_vectorSum_x-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => x_vectorSum_x_start_req,
      start_ack => x_vectorSum_x_start_ack,
      fin_req => x_vectorSum_x_fin_req,
      fin_ack => x_vectorSum_x_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(6 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(6 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(6 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      tag_in => x_vectorSum_x_tag_in,
      tag_out => x_vectorSum_x_tag_out-- 
    ); -- 
  in_data_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_pipe_read_req,
      read_ack => in_data_pipe_pipe_read_ack,
      read_data => in_data_pipe_pipe_read_data,
      write_req => in_data_pipe_pipe_write_req,
      write_ack => in_data_pipe_pipe_write_ack,
      write_data => in_data_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_pipe_read_req,
      read_ack => out_data_pipe_pipe_read_ack,
      read_data => out_data_pipe_pipe_read_data,
      write_req => out_data_pipe_pipe_write_req,
      write_ack => out_data_pipe_pipe_write_ack,
      write_data => out_data_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
