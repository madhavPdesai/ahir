 library ieee;        
 use ieee.std_logic_1164.all;        
 use ieee.numeric_std.all;        
         
 library ahir;        
 use ahir.Types.all;        
 use ahir.Subprograms.all;        
 use ahir.Utilities.all;        
 use ahir.BaseComponents.all;        
  
 entity TB_wrapper is        
   port        
     (all_tests_succeeded : out boolean;        
      all_tests_evaluated : out boolean);        
 end TB_wrapper;        
 
 architecture Behave of TB_wrapper is        
   signal done_flag    : BooleanArray(122 downto 0);        
   signal success_flag : BooleanArray(122 downto 0);        
         
 begin        
  
   tb0 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNot",        
                               tb_id               => "ApIntNot num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(0),        
      all_tests_evaluated => done_flag(0));        
         
   tb1 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNot",        
                               tb_id               => "ApIntNot num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(1),        
      all_tests_evaluated => done_flag(1));        
         
   tb2 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNot",        
                               tb_id               => "ApIntNot num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(2),        
      all_tests_evaluated => done_flag(2));        
  
   tb3 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntSigned",        
                               tb_id               => "ApIntToApIntSigned num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(3),        
      all_tests_evaluated => done_flag(3));        
         
   tb4 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntSigned",        
                               tb_id               => "ApIntToApIntSigned num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(4),        
      all_tests_evaluated => done_flag(4));        
         
   tb5 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntSigned",        
                               tb_id               => "ApIntToApIntSigned num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(5),        
      all_tests_evaluated => done_flag(5));        
  
   tb6 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntUnsigned",        
                               tb_id               => "ApIntToApIntUnsigned num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(6),        
      all_tests_evaluated => done_flag(6));        
         
   tb7 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntUnsigned",        
                               tb_id               => "ApIntToApIntUnsigned num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(7),        
      all_tests_evaluated => done_flag(7));        
         
   tb8 : ApInt_S_1_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntToApIntUnsigned",        
                               tb_id               => "ApIntToApIntUnsigned num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(8),        
      all_tests_evaluated => done_flag(8));        
  
   tb9 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAdd num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(9),        
      all_tests_evaluated => done_flag(9));        
         
   tb10 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAdd num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(10),        
      all_tests_evaluated => done_flag(10));        
         
   tb11 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAdd num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(11),        
      all_tests_evaluated => done_flag(11));        
  
   tb12 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSub num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(12),        
      all_tests_evaluated => done_flag(12));        
         
   tb13 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSub num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(13),        
      all_tests_evaluated => done_flag(13));        
         
   tb14 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSub num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(14),        
      all_tests_evaluated => done_flag(14));        
  
   tb15 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAnd num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(15),        
      all_tests_evaluated => done_flag(15));        
         
   tb16 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAnd num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(16),        
      all_tests_evaluated => done_flag(16));        
         
   tb17 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAnd num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(17),        
      all_tests_evaluated => done_flag(17));        
  
   tb18 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOr num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(18),        
      all_tests_evaluated => done_flag(18));        
         
   tb19 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOr num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(19),        
      all_tests_evaluated => done_flag(19));        
         
   tb20 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOr num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(20),        
      all_tests_evaluated => done_flag(20));        
  
   tb21 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXor num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(21),        
      all_tests_evaluated => done_flag(21));        
         
   tb22 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXor num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(22),        
      all_tests_evaluated => done_flag(22));        
         
   tb23 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXor num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(23),        
      all_tests_evaluated => done_flag(23));        
  
   tb24 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMul num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(24),        
      all_tests_evaluated => done_flag(24));        
         
   tb25 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMul num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(25),        
      all_tests_evaluated => done_flag(25));        
         
   tb26 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMul num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(26),        
      all_tests_evaluated => done_flag(26));        
  
   tb27 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHL num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(27),        
      all_tests_evaluated => done_flag(27));        
         
   tb28 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHL num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(28),        
      all_tests_evaluated => done_flag(28));        
         
   tb29 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHL num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(29),        
      all_tests_evaluated => done_flag(29));        
  
   tb30 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHR num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(30),        
      all_tests_evaluated => done_flag(30));        
         
   tb31 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHR num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(31),        
      all_tests_evaluated => done_flag(31));        
         
   tb32 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHR num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(32),        
      all_tests_evaluated => done_flag(32));        
  
   tb33 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHR num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(33),        
      all_tests_evaluated => done_flag(33));        
         
   tb34 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHR num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(34),        
      all_tests_evaluated => done_flag(34));        
         
   tb35 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHR num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(35),        
      all_tests_evaluated => done_flag(35));        
  
   tb36 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEq num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(36),        
      all_tests_evaluated => done_flag(36));        
         
   tb37 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEq num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(37),        
      all_tests_evaluated => done_flag(37));        
         
   tb38 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEq num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(38),        
      all_tests_evaluated => done_flag(38));        
  
   tb39 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNe num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(39),        
      all_tests_evaluated => done_flag(39));        
         
   tb40 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNe num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(40),        
      all_tests_evaluated => done_flag(40));        
         
   tb41 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNe num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(41),        
      all_tests_evaluated => done_flag(41));        
  
   tb42 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgt num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(42),        
      all_tests_evaluated => done_flag(42));        
         
   tb43 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgt num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(43),        
      all_tests_evaluated => done_flag(43));        
         
   tb44 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgt num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(44),        
      all_tests_evaluated => done_flag(44));        
  
   tb45 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUge num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(45),        
      all_tests_evaluated => done_flag(45));        
         
   tb46 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUge num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(46),        
      all_tests_evaluated => done_flag(46));        
         
   tb47 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUge num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(47),        
      all_tests_evaluated => done_flag(47));        
  
   tb48 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUlt num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(48),        
      all_tests_evaluated => done_flag(48));        
         
   tb49 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUlt num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(49),        
      all_tests_evaluated => done_flag(49));        
         
   tb50 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUlt num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(50),        
      all_tests_evaluated => done_flag(50));        
  
   tb51 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUle num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(51),        
      all_tests_evaluated => done_flag(51));        
         
   tb52 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUle num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(52),        
      all_tests_evaluated => done_flag(52));        
         
   tb53 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUle num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(53),        
      all_tests_evaluated => done_flag(53));        
  
   tb54 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgt num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(54),        
      all_tests_evaluated => done_flag(54));        
         
   tb55 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgt num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(55),        
      all_tests_evaluated => done_flag(55));        
         
   tb56 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgt num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(56),        
      all_tests_evaluated => done_flag(56));        
  
   tb57 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSge num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(57),        
      all_tests_evaluated => done_flag(57));        
         
   tb58 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSge num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(58),        
      all_tests_evaluated => done_flag(58));        
         
   tb59 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSge num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(59),        
      all_tests_evaluated => done_flag(59));        
  
   tb60 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSlt num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(60),        
      all_tests_evaluated => done_flag(60));        
         
   tb61 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSlt num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(61),        
      all_tests_evaluated => done_flag(61));        
         
   tb62 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSlt num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(62),        
      all_tests_evaluated => done_flag(62));        
  
   tb63 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSle num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(63),        
      all_tests_evaluated => done_flag(63));        
         
   tb64 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSle num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(64),        
      all_tests_evaluated => done_flag(64));        
         
   tb65 : ApInt_S_2_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSle num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(65),        
      all_tests_evaluated => done_flag(65));        
  
   tb66 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAddC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(66),        
      all_tests_evaluated => done_flag(66));        
         
   tb67 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAddC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(67),        
      all_tests_evaluated => done_flag(67));        
         
   tb68 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAdd",        
                               tb_id               => "ApIntAddC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(68),        
      all_tests_evaluated => done_flag(68));        
  
   tb69 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSubC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(69),        
      all_tests_evaluated => done_flag(69));        
         
   tb70 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSubC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(70),        
      all_tests_evaluated => done_flag(70));        
         
   tb71 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSub",        
                               tb_id               => "ApIntSubC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(71),        
      all_tests_evaluated => done_flag(71));        
  
   tb72 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAndC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(72),        
      all_tests_evaluated => done_flag(72));        
         
   tb73 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAndC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(73),        
      all_tests_evaluated => done_flag(73));        
         
   tb74 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntAnd",        
                               tb_id               => "ApIntAndC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(74),        
      all_tests_evaluated => done_flag(74));        
  
   tb75 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOrC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(75),        
      all_tests_evaluated => done_flag(75));        
         
   tb76 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOrC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(76),        
      all_tests_evaluated => done_flag(76));        
         
   tb77 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntOr",        
                               tb_id               => "ApIntOrC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(77),        
      all_tests_evaluated => done_flag(77));        
  
   tb78 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXorC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(78),        
      all_tests_evaluated => done_flag(78));        
         
   tb79 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXorC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(79),        
      all_tests_evaluated => done_flag(79));        
         
   tb80 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntXor",        
                               tb_id               => "ApIntXorC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(80),        
      all_tests_evaluated => done_flag(80));        
  
   tb81 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMulC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(81),        
      all_tests_evaluated => done_flag(81));        
         
   tb82 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMulC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(82),        
      all_tests_evaluated => done_flag(82));        
         
   tb83 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntMul",        
                               tb_id               => "ApIntMulC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(83),        
      all_tests_evaluated => done_flag(83));        
  
   tb84 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHLC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(84),        
      all_tests_evaluated => done_flag(84));        
         
   tb85 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHLC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(85),        
      all_tests_evaluated => done_flag(85));        
         
   tb86 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSHL",        
                               tb_id               => "ApIntSHLC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(86),        
      all_tests_evaluated => done_flag(86));        
  
   tb87 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHRC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(87),        
      all_tests_evaluated => done_flag(87));        
         
   tb88 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHRC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(88),        
      all_tests_evaluated => done_flag(88));        
         
   tb89 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntLSHR",        
                               tb_id               => "ApIntLSHRC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(89),        
      all_tests_evaluated => done_flag(89));        
  
   tb90 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHRC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(90),        
      all_tests_evaluated => done_flag(90));        
         
   tb91 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHRC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(91),        
      all_tests_evaluated => done_flag(91));        
         
   tb92 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 8,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntASHR",        
                               tb_id               => "ApIntASHRC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(92),        
      all_tests_evaluated => done_flag(92));        
  
   tb93 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEqC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(93),        
      all_tests_evaluated => done_flag(93));        
         
   tb94 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEqC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(94),        
      all_tests_evaluated => done_flag(94));        
         
   tb95 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntEq",        
                               tb_id               => "ApIntEqC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(95),        
      all_tests_evaluated => done_flag(95));        
  
   tb96 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNeC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(96),        
      all_tests_evaluated => done_flag(96));        
         
   tb97 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNeC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(97),        
      all_tests_evaluated => done_flag(97));        
         
   tb98 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntNe",        
                               tb_id               => "ApIntNeC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(98),        
      all_tests_evaluated => done_flag(98));        
  
   tb99 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgtC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(99),        
      all_tests_evaluated => done_flag(99));        
         
   tb100 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgtC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(100),        
      all_tests_evaluated => done_flag(100));        
         
   tb101 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUgt",        
                               tb_id               => "ApIntUgtC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(101),        
      all_tests_evaluated => done_flag(101));        
  
   tb102 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUgeC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(102),        
      all_tests_evaluated => done_flag(102));        
         
   tb103 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUgeC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(103),        
      all_tests_evaluated => done_flag(103));        
         
   tb104 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUge",        
                               tb_id               => "ApIntUgeC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(104),        
      all_tests_evaluated => done_flag(104));        
  
   tb105 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUltC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(105),        
      all_tests_evaluated => done_flag(105));        
         
   tb106 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUltC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(106),        
      all_tests_evaluated => done_flag(106));        
         
   tb107 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUlt",        
                               tb_id               => "ApIntUltC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(107),        
      all_tests_evaluated => done_flag(107));        
  
   tb108 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUleC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(108),        
      all_tests_evaluated => done_flag(108));        
         
   tb109 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUleC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(109),        
      all_tests_evaluated => done_flag(109));        
         
   tb110 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntUle",        
                               tb_id               => "ApIntUleC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(110),        
      all_tests_evaluated => done_flag(110));        
  
   tb111 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgtC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(111),        
      all_tests_evaluated => done_flag(111));        
         
   tb112 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgtC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(112),        
      all_tests_evaluated => done_flag(112));        
         
   tb113 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSgt",        
                               tb_id               => "ApIntSgtC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(113),        
      all_tests_evaluated => done_flag(113));        
  
   tb114 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSgeC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(114),        
      all_tests_evaluated => done_flag(114));        
         
   tb115 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSgeC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(115),        
      all_tests_evaluated => done_flag(115));        
         
   tb116 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSge",        
                               tb_id               => "ApIntSgeC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(116),        
      all_tests_evaluated => done_flag(116));        
  
   tb117 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSltC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(117),        
      all_tests_evaluated => done_flag(117));        
         
   tb118 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSltC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(118),        
      all_tests_evaluated => done_flag(118));        
         
   tb119 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSlt",        
                               tb_id               => "ApIntSltC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(119),        
      all_tests_evaluated => done_flag(119));        
  
   tb120 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSleC num_req=1"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(120),        
      all_tests_evaluated => done_flag(120));        
         
   tb121 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSleC num_req=2"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(121),        
      all_tests_evaluated => done_flag(121));        
         
   tb122 : ApInt_S_2_C_TB generic map(g_num_req           => 5,        
                               g_input_data_width  => 8,        
                               g_output_data_width => 1,        
                               verbose_mode        => false,        
                               operator_id         => "ApIntSle",        
                               tb_id               => "ApIntSleC num_req=5"        
                               )        
     port map        
     (all_tests_succeeded => success_flag(122),        
      all_tests_evaluated => done_flag(122));        
  
   process(done_flag)        
   begin        
     if(AndReduce(done_flag))then        
       all_tests_evaluated <= true;        
       if(AndReduce(success_flag)) then        
      assert false report "All Tests Have Passed  " severity note;        
      all_tests_succeeded <= true;        
       else        
      assert false report "Some Tests Have Failed " severity error;        
      all_tests_succeeded <= false;        
       end if;        
     else        
       all_tests_evaluated <= false;        
     end if;        
   end process;        
         
 end Behave;        
         
 -------------------------------------------------------        
 configuration conf_TB of TB_wrapper is        
         
   for Behave 
     for tb0 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntNot;        
         end for;        
       end for;        
     end for;	
     for tb1 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntNot;        
         end for;        
       end for;        
     end for; 	
     for tb2 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntNot;        
         end for;        
       end for;        
     end for; 
     for tb3 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntSigned;        
         end for;        
       end for;        
     end for;	
     for tb4 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntSigned;        
         end for;        
       end for;        
     end for; 	
     for tb5 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntSigned;        
         end for;        
       end for;        
     end for; 
     for tb6 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntUnsigned;        
         end for;        
       end for;        
     end for;	
     for tb7 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntUnsigned;        
         end for;        
       end for;        
     end for; 	
     for tb8 : ApInt_S_1_TB        
       for Behave        
         for op2 : ApInt_S_1        
           use configuration ahir.ApIntToApIntUnsigned;        
         end for;        
       end for;        
     end for; 
     for tb9 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAdd;        
         end for;        
       end for;        
     end for;	
     for tb10 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAdd;        
         end for;        
       end for;        
     end for; 	
     for tb11 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAdd;        
         end for;        
       end for;        
     end for; 
     for tb12 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSub;        
         end for;        
       end for;        
     end for;	
     for tb13 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSub;        
         end for;        
       end for;        
     end for; 	
     for tb14 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSub;        
         end for;        
       end for;        
     end for; 
     for tb15 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAnd;        
         end for;        
       end for;        
     end for;	
     for tb16 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAnd;        
         end for;        
       end for;        
     end for; 	
     for tb17 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntAnd;        
         end for;        
       end for;        
     end for; 
     for tb18 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntOr;        
         end for;        
       end for;        
     end for;	
     for tb19 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntOr;        
         end for;        
       end for;        
     end for; 	
     for tb20 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntOr;        
         end for;        
       end for;        
     end for; 
     for tb21 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntXor;        
         end for;        
       end for;        
     end for;	
     for tb22 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntXor;        
         end for;        
       end for;        
     end for; 	
     for tb23 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntXor;        
         end for;        
       end for;        
     end for; 
     for tb24 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntMul;        
         end for;        
       end for;        
     end for;	
     for tb25 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntMul;        
         end for;        
       end for;        
     end for; 	
     for tb26 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntMul;        
         end for;        
       end for;        
     end for; 
     for tb27 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSHL;        
         end for;        
       end for;        
     end for;	
     for tb28 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSHL;        
         end for;        
       end for;        
     end for; 	
     for tb29 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSHL;        
         end for;        
       end for;        
     end for; 
     for tb30 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntLSHR;        
         end for;        
       end for;        
     end for;	
     for tb31 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntLSHR;        
         end for;        
       end for;        
     end for; 	
     for tb32 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntLSHR;        
         end for;        
       end for;        
     end for; 
     for tb33 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntASHR;        
         end for;        
       end for;        
     end for;	
     for tb34 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntASHR;        
         end for;        
       end for;        
     end for; 	
     for tb35 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntASHR;        
         end for;        
       end for;        
     end for; 
     for tb36 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntEq;        
         end for;        
       end for;        
     end for;	
     for tb37 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntEq;        
         end for;        
       end for;        
     end for; 	
     for tb38 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntEq;        
         end for;        
       end for;        
     end for; 
     for tb39 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntNe;        
         end for;        
       end for;        
     end for;	
     for tb40 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntNe;        
         end for;        
       end for;        
     end for; 	
     for tb41 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntNe;        
         end for;        
       end for;        
     end for; 
     for tb42 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUgt;        
         end for;        
       end for;        
     end for;	
     for tb43 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUgt;        
         end for;        
       end for;        
     end for; 	
     for tb44 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUgt;        
         end for;        
       end for;        
     end for; 
     for tb45 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUge;        
         end for;        
       end for;        
     end for;	
     for tb46 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUge;        
         end for;        
       end for;        
     end for; 	
     for tb47 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUge;        
         end for;        
       end for;        
     end for; 
     for tb48 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUlt;        
         end for;        
       end for;        
     end for;	
     for tb49 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUlt;        
         end for;        
       end for;        
     end for; 	
     for tb50 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUlt;        
         end for;        
       end for;        
     end for; 
     for tb51 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUle;        
         end for;        
       end for;        
     end for;	
     for tb52 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUle;        
         end for;        
       end for;        
     end for; 	
     for tb53 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntUle;        
         end for;        
       end for;        
     end for; 
     for tb54 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSgt;        
         end for;        
       end for;        
     end for;	
     for tb55 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSgt;        
         end for;        
       end for;        
     end for; 	
     for tb56 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSgt;        
         end for;        
       end for;        
     end for; 
     for tb57 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSge;        
         end for;        
       end for;        
     end for;	
     for tb58 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSge;        
         end for;        
       end for;        
     end for; 	
     for tb59 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSge;        
         end for;        
       end for;        
     end for; 
     for tb60 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSlt;        
         end for;        
       end for;        
     end for;	
     for tb61 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSlt;        
         end for;        
       end for;        
     end for; 	
     for tb62 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSlt;        
         end for;        
       end for;        
     end for; 
     for tb63 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSle;        
         end for;        
       end for;        
     end for;	
     for tb64 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSle;        
         end for;        
       end for;        
     end for; 	
     for tb65 : ApInt_S_2_TB        
       for Behave        
         for op2 : ApInt_S_2        
           use configuration ahir.ApIntSle;        
         end for;        
       end for;        
     end for; 
     for tb66 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAddC;        
         end for;        
       end for;        
     end for;	
     for tb67 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAddC;        
         end for;        
       end for;        
     end for; 	
     for tb68 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAddC;        
         end for;        
       end for;        
     end for; 
     for tb69 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSubC;        
         end for;        
       end for;        
     end for;	
     for tb70 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSubC;        
         end for;        
       end for;        
     end for; 	
     for tb71 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSubC;        
         end for;        
       end for;        
     end for; 
     for tb72 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAndC;        
         end for;        
       end for;        
     end for;	
     for tb73 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAndC;        
         end for;        
       end for;        
     end for; 	
     for tb74 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntAndC;        
         end for;        
       end for;        
     end for; 
     for tb75 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntOrC;        
         end for;        
       end for;        
     end for;	
     for tb76 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntOrC;        
         end for;        
       end for;        
     end for; 	
     for tb77 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntOrC;        
         end for;        
       end for;        
     end for; 
     for tb78 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntXorC;        
         end for;        
       end for;        
     end for;	
     for tb79 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntXorC;        
         end for;        
       end for;        
     end for; 	
     for tb80 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntXorC;        
         end for;        
       end for;        
     end for; 
     for tb81 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntMulC;        
         end for;        
       end for;        
     end for;	
     for tb82 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntMulC;        
         end for;        
       end for;        
     end for; 	
     for tb83 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntMulC;        
         end for;        
       end for;        
     end for; 
     for tb84 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSHLC;        
         end for;        
       end for;        
     end for;	
     for tb85 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSHLC;        
         end for;        
       end for;        
     end for; 	
     for tb86 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSHLC;        
         end for;        
       end for;        
     end for; 
     for tb87 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntLSHRC;        
         end for;        
       end for;        
     end for;	
     for tb88 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntLSHRC;        
         end for;        
       end for;        
     end for; 	
     for tb89 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntLSHRC;        
         end for;        
       end for;        
     end for; 
     for tb90 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntASHRC;        
         end for;        
       end for;        
     end for;	
     for tb91 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntASHRC;        
         end for;        
       end for;        
     end for; 	
     for tb92 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntASHRC;        
         end for;        
       end for;        
     end for; 
     for tb93 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntEqC;        
         end for;        
       end for;        
     end for;	
     for tb94 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntEqC;        
         end for;        
       end for;        
     end for; 	
     for tb95 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntEqC;        
         end for;        
       end for;        
     end for; 
     for tb96 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntNeC;        
         end for;        
       end for;        
     end for;	
     for tb97 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntNeC;        
         end for;        
       end for;        
     end for; 	
     for tb98 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntNeC;        
         end for;        
       end for;        
     end for; 
     for tb99 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgtC;        
         end for;        
       end for;        
     end for;	
     for tb100 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgtC;        
         end for;        
       end for;        
     end for; 	
     for tb101 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgtC;        
         end for;        
       end for;        
     end for; 
     for tb102 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgeC;        
         end for;        
       end for;        
     end for;	
     for tb103 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgeC;        
         end for;        
       end for;        
     end for; 	
     for tb104 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUgeC;        
         end for;        
       end for;        
     end for; 
     for tb105 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUltC;        
         end for;        
       end for;        
     end for;	
     for tb106 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUltC;        
         end for;        
       end for;        
     end for; 	
     for tb107 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUltC;        
         end for;        
       end for;        
     end for; 
     for tb108 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUleC;        
         end for;        
       end for;        
     end for;	
     for tb109 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUleC;        
         end for;        
       end for;        
     end for; 	
     for tb110 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntUleC;        
         end for;        
       end for;        
     end for; 
     for tb111 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgtC;        
         end for;        
       end for;        
     end for;	
     for tb112 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgtC;        
         end for;        
       end for;        
     end for; 	
     for tb113 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgtC;        
         end for;        
       end for;        
     end for; 
     for tb114 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgeC;        
         end for;        
       end for;        
     end for;	
     for tb115 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgeC;        
         end for;        
       end for;        
     end for; 	
     for tb116 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSgeC;        
         end for;        
       end for;        
     end for; 
     for tb117 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSltC;        
         end for;        
       end for;        
     end for;	
     for tb118 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSltC;        
         end for;        
       end for;        
     end for; 	
     for tb119 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSltC;        
         end for;        
       end for;        
     end for; 
     for tb120 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSleC;        
         end for;        
       end for;        
     end for;	
     for tb121 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSleC;        
         end for;        
       end for;        
     end for; 	
     for tb122 : ApInt_S_2_C_TB        
       for Behave        
         for op2 : ApInt_S_2_C        
           use configuration ahir.ApIntSleC;        
         end for;        
       end for;        
     end for;
   end for;        
         
 end conf_TB;
