------------------------------------------------------------------------------------------------
--
-- Copyright (C) 2010-: Madhav P. Desai
-- All Rights Reserved.
--  
-- Permission is hereby granted, free of charge, to any person obtaining a
-- copy of this software and associated documentation files (the
-- "Software"), to deal with the Software without restriction, including
-- without limitation the rights to use, copy, modify, merge, publish,
-- distribute, sublicense, and/or sell copies of the Software, and to
-- permit persons to whom the Software is furnished to do so, subject to
-- the following conditions:
-- 
--  * Redistributions of source code must retain the above copyright
--    notice, this list of conditions and the following disclaimers.
--  * Redistributions in binary form must reproduce the above
--    copyright notice, this list of conditions and the following
--    disclaimers in the documentation and/or other materials provided
--    with the distribution.
--  * Neither the names of the AHIR Team, the Indian Institute of
--    Technology Bombay, nor the names of its contributors may be used
--    to endorse or promote products derived from this Software
--    without specific prior written permission.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
-- OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
library work;
use work.vc_system_package.all;
entity foo is -- 
  port ( -- 
    a : in  std_logic_vector(31 downto 0);
    b : in  std_logic_vector(31 downto 0);
    c : out  std_logic_vector(31 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start : in std_logic;
    fin   : out std_logic;
    tag_in: in std_logic_vector(0 downto 0);
    tag_out: out std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity foo;
architecture Default of foo is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  -- links between control-path and data-path
  signal a_gt_b_ack_0 : boolean;
  signal a_gt_b_req_1 : boolean;
  signal branch_req_0 : boolean;
  signal a_gt_b_req_0 : boolean;
  signal sub1_ack_0 : boolean;
  signal sub1_req_1 : boolean;
  signal a_gt_b_ack_1 : boolean;
  signal branch_ack_0 : boolean;
  signal sub0_ack_1 : boolean;
  signal sub0_req_0 : boolean;
  signal sub0_ack_0 : boolean;
  signal sub0_req_1 : boolean;
  signal branch_ack_1 : boolean;
  signal sub1_ack_1 : boolean;
  signal sub1_req_0 : boolean;
  signal resolve_ack_0 : boolean;
  -- 
begin --  
  -- tag register
  process(clk) 
  begin -- 
    if clk'event and clk = '1' then -- 
      if start='1' then -- 
        tag_out <= tag_in; -- 
      end if; -- 
    end if; -- 
  end process;
  -- the control path
  always_true_symbol <= true; 
  foo_CP_0: Block -- control-path 
    signal cp_elements: BooleanArray(10 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= true when start = '1' else false;
    fin <= '1' when cp_elements(10) else '0';
    a_gt_b_req_0 <= cp_elements(0);
    cp_elements(1) <= a_gt_b_ack_0;
    a_gt_b_req_1 <= cp_elements(1);
    cp_elements(2) <= a_gt_b_ack_1;
    branch_req_0 <= cp_elements(2);
    cp_elements(3) <= branch_ack_0;
    sub0_req_0 <= cp_elements(3);
    cp_elements(4) <= sub0_ack_0;
    sub0_req_1 <= cp_elements(4);
    cp_elements(5) <= sub0_ack_1;
    resolve_req_0 <= cp_elements(5);
    cp_elements(6) <= branch_ack_1;
    sub1_req_0 <= cp_elements(6);
    cp_elements(7) <= sub1_ack_0;
    sub1_req_1 <= cp_elements(7);
    cp_elements(8) <= sub1_ack_1;
    resolve_req_1 <= cp_elements(8);
    cp_elements(9) <= OrReduce(cp_elements(8) & cp_elements(5));
    cp_elements(10) <= resolve_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal p : std_logic_vector(0 downto 0);
    signal q : std_logic_vector(31 downto 0);
    signal r : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    resolve: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= q & r;
      req <= resolve_req_0 & resolve_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => resolve_ack_0,
          idata => idata,
          odata => c,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator resolve
    branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(31 downto 0);
      begin 
      condition_sig <= a;
      branch_instance: BranchBase -- 
        generic map( condition_width => 32)
        port map( -- 
          condition => condition_sig,
          req => branch_req_0,
          ack0 => branch_ack_0,
          ack1 => branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : a_gt_b 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a & b;
      p <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => a_gt_b_req_0,
          ackL => a_gt_b_ack_0,
          reqR => a_gt_b_req_1,
          ackR => a_gt_b_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : sub1 sub0 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= a & b & b & a;
      q <= data_out(63 downto 32);
      r <= data_out(31 downto 0);
      reqL(1) <= sub1_req_0;
      reqL(0) <= sub0_req_0;
      sub1_ack_0 <= ackL(1);
      sub0_ack_0 <= ackL(0);
      reqR(1) <= sub1_req_1;
      reqR(0) <= sub0_req_1;
      sub1_ack_1 <= ackR(1);
      sub0_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true, 
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
library work;
use work.vc_system_package.all;
entity test_system is  -- system 
  port (-- 
    foo_a : in  std_logic_vector(31 downto 0);
    foo_b : in  std_logic_vector(31 downto 0);
    foo_c : out  std_logic_vector(31 downto 0);
    foo_tag_in: in std_logic_vector(0 downto 0);
    foo_tag_out: out std_logic_vector(0 downto 0);
    foo_start : in std_logic;
    foo_fin   : out std_logic;
    clk : in std_logic;
    reset : in std_logic); -- 
  -- 
end entity; 
architecture Default of test_system is -- system-architecture 
  -- declarations related to module foo
  component foo is -- 
    port ( -- 
      a : in  std_logic_vector(31 downto 0);
      b : in  std_logic_vector(31 downto 0);
      c : out  std_logic_vector(31 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start : in std_logic;
      fin   : out std_logic;
      tag_in: in std_logic_vector(0 downto 0);
      tag_out: out std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component;
  -- 
begin -- 
  -- module foo
  foo_instance:foo-- 
    port map(-- 
      a => foo_a,
      b => foo_b,
      c => foo_c,
      start => foo_start,
      fin => foo_fin,
      clk => clk,
      reset => reset,
      tag_in => foo_tag_in,
      tag_out => foo_tag_out-- 
    ); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
library work;
use work.vc_system_package.all;
entity test_system_Test_Bench is -- 
  -- 
end entity;
architecture Default of test_system_Test_Bench is -- 
  component test_system is -- 
    port (-- 
      foo_a : in  std_logic_vector(31 downto 0);
      foo_b : in  std_logic_vector(31 downto 0);
      foo_c : out  std_logic_vector(31 downto 0);
      foo_tag_in: in std_logic_vector(0 downto 0);
      foo_tag_out: out std_logic_vector(0 downto 0);
      foo_start : in std_logic;
      foo_fin   : out std_logic;
      clk : in std_logic;
      reset : in std_logic); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal foo_a :  std_logic_vector(31 downto 0) := (others => '0');
  signal foo_b :  std_logic_vector(31 downto 0) := (others => '0');
  signal foo_c :   std_logic_vector(31 downto 0);
  signal foo_tag_in: std_logic_vector(0 downto 0);
  signal foo_tag_out: std_logic_vector(0 downto 0);
  signal foo_start : std_logic := '0';
  signal foo_fin   : std_logic := '0';
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  process
  begin --
    wait until clk = '1';
    reset <= '0';
    wait;
    --
  end process;
  -- a rudimentary tb.. will start all the top-level modules ..
  process
  begin --
    wait until clk = '1';
    foo_start <= '1';
    wait until clk = '1';
    foo_start <= '0';
    while foo_fin /= '1' loop -- 
      wait until clk = '1';
      -- 
    end loop;
    wait;
    --
  end process;
  test_system_instance: test_system -- 
    port map ( -- 
      foo_a => foo_a,
      foo_b => foo_b,
      foo_c => foo_c,
      foo_tag_in => foo_tag_in,
      foo_tag_out => foo_tag_out,
      foo_start => foo_start,
      foo_fin  => foo_fin ,
      clk => clk,
      reset => reset); -- 
  -- 
end Default;
