
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;
use ahir.components.all;

entity start_cp is
  port(
    LambdaIn : in BooleanArray(292 downto 1);
    LambdaOut : out BooleanArray(294 downto 1);
    clk : in std_logic;
    reset : in std_logic);
end start_cp;

architecture default_arch of start_cp is
  signal place_0_preds : BooleanArray(0 downto 0);
  signal place_0_succs : BooleanArray(0 downto 0);
  signal place_0_token : boolean;
  signal place_6_preds : BooleanArray(0 downto 0);
  signal place_6_succs : BooleanArray(1 downto 0);
  signal place_6_token : boolean;
  signal place_13_preds : BooleanArray(0 downto 0);
  signal place_13_succs : BooleanArray(1 downto 0);
  signal place_13_token : boolean;
  signal place_18_preds : BooleanArray(0 downto 0);
  signal place_18_succs : BooleanArray(0 downto 0);
  signal place_18_token : boolean;
  signal place_24_preds : BooleanArray(1 downto 0);
  signal place_24_succs : BooleanArray(0 downto 0);
  signal place_24_token : boolean;
  signal place_28_preds : BooleanArray(1 downto 0);
  signal place_28_succs : BooleanArray(0 downto 0);
  signal place_28_token : boolean;
  signal place_36_preds : BooleanArray(0 downto 0);
  signal place_36_succs : BooleanArray(0 downto 0);
  signal place_36_token : boolean;
  signal place_37_preds : BooleanArray(0 downto 0);
  signal place_37_succs : BooleanArray(0 downto 0);
  signal place_37_token : boolean;
  signal place_38_preds : BooleanArray(0 downto 0);
  signal place_38_succs : BooleanArray(0 downto 0);
  signal place_38_token : boolean;
  signal place_43_preds : BooleanArray(0 downto 0);
  signal place_43_succs : BooleanArray(0 downto 0);
  signal place_43_token : boolean;
  signal place_44_preds : BooleanArray(0 downto 0);
  signal place_44_succs : BooleanArray(0 downto 0);
  signal place_44_token : boolean;
  signal place_45_preds : BooleanArray(0 downto 0);
  signal place_45_succs : BooleanArray(0 downto 0);
  signal place_45_token : boolean;
  signal place_50_preds : BooleanArray(0 downto 0);
  signal place_50_succs : BooleanArray(0 downto 0);
  signal place_50_token : boolean;
  signal place_51_preds : BooleanArray(0 downto 0);
  signal place_51_succs : BooleanArray(0 downto 0);
  signal place_51_token : boolean;
  signal place_52_preds : BooleanArray(0 downto 0);
  signal place_52_succs : BooleanArray(0 downto 0);
  signal place_52_token : boolean;
  signal place_58_preds : BooleanArray(0 downto 0);
  signal place_58_succs : BooleanArray(0 downto 0);
  signal place_58_token : boolean;
  signal place_59_preds : BooleanArray(0 downto 0);
  signal place_59_succs : BooleanArray(0 downto 0);
  signal place_59_token : boolean;
  signal place_60_preds : BooleanArray(0 downto 0);
  signal place_60_succs : BooleanArray(0 downto 0);
  signal place_60_token : boolean;
  signal place_65_preds : BooleanArray(0 downto 0);
  signal place_65_succs : BooleanArray(0 downto 0);
  signal place_65_token : boolean;
  signal place_66_preds : BooleanArray(0 downto 0);
  signal place_66_succs : BooleanArray(0 downto 0);
  signal place_66_token : boolean;
  signal place_67_preds : BooleanArray(0 downto 0);
  signal place_67_succs : BooleanArray(0 downto 0);
  signal place_67_token : boolean;
  signal place_73_preds : BooleanArray(0 downto 0);
  signal place_73_succs : BooleanArray(0 downto 0);
  signal place_73_token : boolean;
  signal place_74_preds : BooleanArray(0 downto 0);
  signal place_74_succs : BooleanArray(0 downto 0);
  signal place_74_token : boolean;
  signal place_75_preds : BooleanArray(0 downto 0);
  signal place_75_succs : BooleanArray(0 downto 0);
  signal place_75_token : boolean;
  signal place_80_preds : BooleanArray(0 downto 0);
  signal place_80_succs : BooleanArray(0 downto 0);
  signal place_80_token : boolean;
  signal place_81_preds : BooleanArray(0 downto 0);
  signal place_81_succs : BooleanArray(0 downto 0);
  signal place_81_token : boolean;
  signal place_82_preds : BooleanArray(0 downto 0);
  signal place_82_succs : BooleanArray(0 downto 0);
  signal place_82_token : boolean;
  signal place_87_preds : BooleanArray(0 downto 0);
  signal place_87_succs : BooleanArray(0 downto 0);
  signal place_87_token : boolean;
  signal place_88_preds : BooleanArray(0 downto 0);
  signal place_88_succs : BooleanArray(0 downto 0);
  signal place_88_token : boolean;
  signal place_89_preds : BooleanArray(0 downto 0);
  signal place_89_succs : BooleanArray(0 downto 0);
  signal place_89_token : boolean;
  signal place_94_preds : BooleanArray(0 downto 0);
  signal place_94_succs : BooleanArray(0 downto 0);
  signal place_94_token : boolean;
  signal place_95_preds : BooleanArray(0 downto 0);
  signal place_95_succs : BooleanArray(0 downto 0);
  signal place_95_token : boolean;
  signal place_96_preds : BooleanArray(0 downto 0);
  signal place_96_succs : BooleanArray(0 downto 0);
  signal place_96_token : boolean;
  signal place_102_preds : BooleanArray(0 downto 0);
  signal place_102_succs : BooleanArray(0 downto 0);
  signal place_102_token : boolean;
  signal place_103_preds : BooleanArray(0 downto 0);
  signal place_103_succs : BooleanArray(0 downto 0);
  signal place_103_token : boolean;
  signal place_104_preds : BooleanArray(0 downto 0);
  signal place_104_succs : BooleanArray(0 downto 0);
  signal place_104_token : boolean;
  signal place_109_preds : BooleanArray(0 downto 0);
  signal place_109_succs : BooleanArray(0 downto 0);
  signal place_109_token : boolean;
  signal place_110_preds : BooleanArray(0 downto 0);
  signal place_110_succs : BooleanArray(0 downto 0);
  signal place_110_token : boolean;
  signal place_111_preds : BooleanArray(0 downto 0);
  signal place_111_succs : BooleanArray(0 downto 0);
  signal place_111_token : boolean;
  signal place_117_preds : BooleanArray(0 downto 0);
  signal place_117_succs : BooleanArray(0 downto 0);
  signal place_117_token : boolean;
  signal place_118_preds : BooleanArray(0 downto 0);
  signal place_118_succs : BooleanArray(0 downto 0);
  signal place_118_token : boolean;
  signal place_119_preds : BooleanArray(0 downto 0);
  signal place_119_succs : BooleanArray(0 downto 0);
  signal place_119_token : boolean;
  signal place_124_preds : BooleanArray(0 downto 0);
  signal place_124_succs : BooleanArray(0 downto 0);
  signal place_124_token : boolean;
  signal place_125_preds : BooleanArray(0 downto 0);
  signal place_125_succs : BooleanArray(0 downto 0);
  signal place_125_token : boolean;
  signal place_126_preds : BooleanArray(0 downto 0);
  signal place_126_succs : BooleanArray(0 downto 0);
  signal place_126_token : boolean;
  signal place_131_preds : BooleanArray(0 downto 0);
  signal place_131_succs : BooleanArray(0 downto 0);
  signal place_131_token : boolean;
  signal place_132_preds : BooleanArray(0 downto 0);
  signal place_132_succs : BooleanArray(0 downto 0);
  signal place_132_token : boolean;
  signal place_133_preds : BooleanArray(0 downto 0);
  signal place_133_succs : BooleanArray(0 downto 0);
  signal place_133_token : boolean;
  signal place_138_preds : BooleanArray(0 downto 0);
  signal place_138_succs : BooleanArray(0 downto 0);
  signal place_138_token : boolean;
  signal place_139_preds : BooleanArray(0 downto 0);
  signal place_139_succs : BooleanArray(0 downto 0);
  signal place_139_token : boolean;
  signal place_140_preds : BooleanArray(0 downto 0);
  signal place_140_succs : BooleanArray(0 downto 0);
  signal place_140_token : boolean;
  signal place_146_preds : BooleanArray(0 downto 0);
  signal place_146_succs : BooleanArray(0 downto 0);
  signal place_146_token : boolean;
  signal place_147_preds : BooleanArray(0 downto 0);
  signal place_147_succs : BooleanArray(0 downto 0);
  signal place_147_token : boolean;
  signal place_148_preds : BooleanArray(0 downto 0);
  signal place_148_succs : BooleanArray(0 downto 0);
  signal place_148_token : boolean;
  signal place_153_preds : BooleanArray(0 downto 0);
  signal place_153_succs : BooleanArray(0 downto 0);
  signal place_153_token : boolean;
  signal place_154_preds : BooleanArray(0 downto 0);
  signal place_154_succs : BooleanArray(0 downto 0);
  signal place_154_token : boolean;
  signal place_155_preds : BooleanArray(0 downto 0);
  signal place_155_succs : BooleanArray(0 downto 0);
  signal place_155_token : boolean;
  signal place_160_preds : BooleanArray(0 downto 0);
  signal place_160_succs : BooleanArray(0 downto 0);
  signal place_160_token : boolean;
  signal place_161_preds : BooleanArray(0 downto 0);
  signal place_161_succs : BooleanArray(0 downto 0);
  signal place_161_token : boolean;
  signal place_162_preds : BooleanArray(0 downto 0);
  signal place_162_succs : BooleanArray(0 downto 0);
  signal place_162_token : boolean;
  signal place_165_preds : BooleanArray(0 downto 0);
  signal place_165_succs : BooleanArray(0 downto 0);
  signal place_165_token : boolean;
  signal place_173_preds : BooleanArray(0 downto 0);
  signal place_173_succs : BooleanArray(0 downto 0);
  signal place_173_token : boolean;
  signal place_174_preds : BooleanArray(0 downto 0);
  signal place_174_succs : BooleanArray(0 downto 0);
  signal place_174_token : boolean;
  signal place_175_preds : BooleanArray(0 downto 0);
  signal place_175_succs : BooleanArray(0 downto 0);
  signal place_175_token : boolean;
  signal place_180_preds : BooleanArray(0 downto 0);
  signal place_180_succs : BooleanArray(0 downto 0);
  signal place_180_token : boolean;
  signal place_181_preds : BooleanArray(0 downto 0);
  signal place_181_succs : BooleanArray(0 downto 0);
  signal place_181_token : boolean;
  signal place_182_preds : BooleanArray(0 downto 0);
  signal place_182_succs : BooleanArray(0 downto 0);
  signal place_182_token : boolean;
  signal place_187_preds : BooleanArray(0 downto 0);
  signal place_187_succs : BooleanArray(0 downto 0);
  signal place_187_token : boolean;
  signal place_188_preds : BooleanArray(0 downto 0);
  signal place_188_succs : BooleanArray(0 downto 0);
  signal place_188_token : boolean;
  signal place_189_preds : BooleanArray(0 downto 0);
  signal place_189_succs : BooleanArray(0 downto 0);
  signal place_189_token : boolean;
  signal place_195_preds : BooleanArray(0 downto 0);
  signal place_195_succs : BooleanArray(0 downto 0);
  signal place_195_token : boolean;
  signal place_196_preds : BooleanArray(0 downto 0);
  signal place_196_succs : BooleanArray(0 downto 0);
  signal place_196_token : boolean;
  signal place_197_preds : BooleanArray(0 downto 0);
  signal place_197_succs : BooleanArray(0 downto 0);
  signal place_197_token : boolean;
  signal place_202_preds : BooleanArray(0 downto 0);
  signal place_202_succs : BooleanArray(0 downto 0);
  signal place_202_token : boolean;
  signal place_203_preds : BooleanArray(0 downto 0);
  signal place_203_succs : BooleanArray(0 downto 0);
  signal place_203_token : boolean;
  signal place_204_preds : BooleanArray(0 downto 0);
  signal place_204_succs : BooleanArray(0 downto 0);
  signal place_204_token : boolean;
  signal place_209_preds : BooleanArray(0 downto 0);
  signal place_209_succs : BooleanArray(0 downto 0);
  signal place_209_token : boolean;
  signal place_210_preds : BooleanArray(0 downto 0);
  signal place_210_succs : BooleanArray(0 downto 0);
  signal place_210_token : boolean;
  signal place_211_preds : BooleanArray(0 downto 0);
  signal place_211_succs : BooleanArray(0 downto 0);
  signal place_211_token : boolean;
  signal place_213_preds : BooleanArray(0 downto 0);
  signal place_213_succs : BooleanArray(0 downto 0);
  signal place_213_token : boolean;
  signal place_221_preds : BooleanArray(0 downto 0);
  signal place_221_succs : BooleanArray(0 downto 0);
  signal place_221_token : boolean;
  signal place_222_preds : BooleanArray(0 downto 0);
  signal place_222_succs : BooleanArray(0 downto 0);
  signal place_222_token : boolean;
  signal place_223_preds : BooleanArray(0 downto 0);
  signal place_223_succs : BooleanArray(0 downto 0);
  signal place_223_token : boolean;
  signal place_228_preds : BooleanArray(0 downto 0);
  signal place_228_succs : BooleanArray(0 downto 0);
  signal place_228_token : boolean;
  signal place_229_preds : BooleanArray(0 downto 0);
  signal place_229_succs : BooleanArray(0 downto 0);
  signal place_229_token : boolean;
  signal place_230_preds : BooleanArray(0 downto 0);
  signal place_230_succs : BooleanArray(0 downto 0);
  signal place_230_token : boolean;
  signal place_232_preds : BooleanArray(1 downto 0);
  signal place_232_succs : BooleanArray(0 downto 0);
  signal place_232_token : boolean;
  signal place_236_preds : BooleanArray(1 downto 0);
  signal place_236_succs : BooleanArray(0 downto 0);
  signal place_236_token : boolean;
  signal place_244_preds : BooleanArray(0 downto 0);
  signal place_244_succs : BooleanArray(0 downto 0);
  signal place_244_token : boolean;
  signal place_245_preds : BooleanArray(0 downto 0);
  signal place_245_succs : BooleanArray(0 downto 0);
  signal place_245_token : boolean;
  signal place_246_preds : BooleanArray(0 downto 0);
  signal place_246_succs : BooleanArray(0 downto 0);
  signal place_246_token : boolean;
  signal place_251_preds : BooleanArray(0 downto 0);
  signal place_251_succs : BooleanArray(0 downto 0);
  signal place_251_token : boolean;
  signal place_252_preds : BooleanArray(0 downto 0);
  signal place_252_succs : BooleanArray(0 downto 0);
  signal place_252_token : boolean;
  signal place_253_preds : BooleanArray(0 downto 0);
  signal place_253_succs : BooleanArray(0 downto 0);
  signal place_253_token : boolean;
  signal place_258_preds : BooleanArray(0 downto 0);
  signal place_258_succs : BooleanArray(0 downto 0);
  signal place_258_token : boolean;
  signal place_259_preds : BooleanArray(0 downto 0);
  signal place_259_succs : BooleanArray(0 downto 0);
  signal place_259_token : boolean;
  signal place_260_preds : BooleanArray(0 downto 0);
  signal place_260_succs : BooleanArray(0 downto 0);
  signal place_260_token : boolean;
  signal place_266_preds : BooleanArray(0 downto 0);
  signal place_266_succs : BooleanArray(0 downto 0);
  signal place_266_token : boolean;
  signal place_267_preds : BooleanArray(0 downto 0);
  signal place_267_succs : BooleanArray(0 downto 0);
  signal place_267_token : boolean;
  signal place_268_preds : BooleanArray(0 downto 0);
  signal place_268_succs : BooleanArray(0 downto 0);
  signal place_268_token : boolean;
  signal place_273_preds : BooleanArray(0 downto 0);
  signal place_273_succs : BooleanArray(0 downto 0);
  signal place_273_token : boolean;
  signal place_274_preds : BooleanArray(0 downto 0);
  signal place_274_succs : BooleanArray(0 downto 0);
  signal place_274_token : boolean;
  signal place_275_preds : BooleanArray(0 downto 0);
  signal place_275_succs : BooleanArray(0 downto 0);
  signal place_275_token : boolean;
  signal place_281_preds : BooleanArray(0 downto 0);
  signal place_281_succs : BooleanArray(0 downto 0);
  signal place_281_token : boolean;
  signal place_282_preds : BooleanArray(0 downto 0);
  signal place_282_succs : BooleanArray(0 downto 0);
  signal place_282_token : boolean;
  signal place_283_preds : BooleanArray(0 downto 0);
  signal place_283_succs : BooleanArray(0 downto 0);
  signal place_283_token : boolean;
  signal place_288_preds : BooleanArray(0 downto 0);
  signal place_288_succs : BooleanArray(0 downto 0);
  signal place_288_token : boolean;
  signal place_289_preds : BooleanArray(0 downto 0);
  signal place_289_succs : BooleanArray(0 downto 0);
  signal place_289_token : boolean;
  signal place_290_preds : BooleanArray(0 downto 0);
  signal place_290_succs : BooleanArray(0 downto 0);
  signal place_290_token : boolean;
  signal place_295_preds : BooleanArray(0 downto 0);
  signal place_295_succs : BooleanArray(0 downto 0);
  signal place_295_token : boolean;
  signal place_296_preds : BooleanArray(0 downto 0);
  signal place_296_succs : BooleanArray(0 downto 0);
  signal place_296_token : boolean;
  signal place_297_preds : BooleanArray(0 downto 0);
  signal place_297_succs : BooleanArray(0 downto 0);
  signal place_297_token : boolean;
  signal place_302_preds : BooleanArray(0 downto 0);
  signal place_302_succs : BooleanArray(0 downto 0);
  signal place_302_token : boolean;
  signal place_303_preds : BooleanArray(0 downto 0);
  signal place_303_succs : BooleanArray(0 downto 0);
  signal place_303_token : boolean;
  signal place_304_preds : BooleanArray(0 downto 0);
  signal place_304_succs : BooleanArray(0 downto 0);
  signal place_304_token : boolean;
  signal place_310_preds : BooleanArray(0 downto 0);
  signal place_310_succs : BooleanArray(0 downto 0);
  signal place_310_token : boolean;
  signal place_311_preds : BooleanArray(0 downto 0);
  signal place_311_succs : BooleanArray(0 downto 0);
  signal place_311_token : boolean;
  signal place_312_preds : BooleanArray(0 downto 0);
  signal place_312_succs : BooleanArray(0 downto 0);
  signal place_312_token : boolean;
  signal place_317_preds : BooleanArray(0 downto 0);
  signal place_317_succs : BooleanArray(0 downto 0);
  signal place_317_token : boolean;
  signal place_318_preds : BooleanArray(0 downto 0);
  signal place_318_succs : BooleanArray(0 downto 0);
  signal place_318_token : boolean;
  signal place_319_preds : BooleanArray(0 downto 0);
  signal place_319_succs : BooleanArray(0 downto 0);
  signal place_319_token : boolean;
  signal place_325_preds : BooleanArray(0 downto 0);
  signal place_325_succs : BooleanArray(0 downto 0);
  signal place_325_token : boolean;
  signal place_326_preds : BooleanArray(0 downto 0);
  signal place_326_succs : BooleanArray(0 downto 0);
  signal place_326_token : boolean;
  signal place_327_preds : BooleanArray(0 downto 0);
  signal place_327_succs : BooleanArray(0 downto 0);
  signal place_327_token : boolean;
  signal place_332_preds : BooleanArray(0 downto 0);
  signal place_332_succs : BooleanArray(0 downto 0);
  signal place_332_token : boolean;
  signal place_333_preds : BooleanArray(0 downto 0);
  signal place_333_succs : BooleanArray(0 downto 0);
  signal place_333_token : boolean;
  signal place_334_preds : BooleanArray(0 downto 0);
  signal place_334_succs : BooleanArray(0 downto 0);
  signal place_334_token : boolean;
  signal place_339_preds : BooleanArray(0 downto 0);
  signal place_339_succs : BooleanArray(0 downto 0);
  signal place_339_token : boolean;
  signal place_340_preds : BooleanArray(0 downto 0);
  signal place_340_succs : BooleanArray(0 downto 0);
  signal place_340_token : boolean;
  signal place_341_preds : BooleanArray(0 downto 0);
  signal place_341_succs : BooleanArray(0 downto 0);
  signal place_341_token : boolean;
  signal place_346_preds : BooleanArray(0 downto 0);
  signal place_346_succs : BooleanArray(0 downto 0);
  signal place_346_token : boolean;
  signal place_347_preds : BooleanArray(0 downto 0);
  signal place_347_succs : BooleanArray(0 downto 0);
  signal place_347_token : boolean;
  signal place_348_preds : BooleanArray(0 downto 0);
  signal place_348_succs : BooleanArray(0 downto 0);
  signal place_348_token : boolean;
  signal place_354_preds : BooleanArray(0 downto 0);
  signal place_354_succs : BooleanArray(0 downto 0);
  signal place_354_token : boolean;
  signal place_355_preds : BooleanArray(0 downto 0);
  signal place_355_succs : BooleanArray(0 downto 0);
  signal place_355_token : boolean;
  signal place_356_preds : BooleanArray(0 downto 0);
  signal place_356_succs : BooleanArray(0 downto 0);
  signal place_356_token : boolean;
  signal place_361_preds : BooleanArray(0 downto 0);
  signal place_361_succs : BooleanArray(0 downto 0);
  signal place_361_token : boolean;
  signal place_362_preds : BooleanArray(0 downto 0);
  signal place_362_succs : BooleanArray(0 downto 0);
  signal place_362_token : boolean;
  signal place_363_preds : BooleanArray(0 downto 0);
  signal place_363_succs : BooleanArray(0 downto 0);
  signal place_363_token : boolean;
  signal place_368_preds : BooleanArray(0 downto 0);
  signal place_368_succs : BooleanArray(0 downto 0);
  signal place_368_token : boolean;
  signal place_369_preds : BooleanArray(0 downto 0);
  signal place_369_succs : BooleanArray(0 downto 0);
  signal place_369_token : boolean;
  signal place_370_preds : BooleanArray(0 downto 0);
  signal place_370_succs : BooleanArray(0 downto 0);
  signal place_370_token : boolean;
  signal place_377_preds : BooleanArray(0 downto 0);
  signal place_377_succs : BooleanArray(0 downto 0);
  signal place_377_token : boolean;
  signal place_378_preds : BooleanArray(0 downto 0);
  signal place_378_succs : BooleanArray(0 downto 0);
  signal place_378_token : boolean;
  signal place_379_preds : BooleanArray(0 downto 0);
  signal place_379_succs : BooleanArray(0 downto 0);
  signal place_379_token : boolean;
  signal place_380_preds : BooleanArray(0 downto 0);
  signal place_380_succs : BooleanArray(0 downto 0);
  signal place_380_token : boolean;
  signal place_388_preds : BooleanArray(0 downto 0);
  signal place_388_succs : BooleanArray(0 downto 0);
  signal place_388_token : boolean;
  signal place_389_preds : BooleanArray(0 downto 0);
  signal place_389_succs : BooleanArray(0 downto 0);
  signal place_389_token : boolean;
  signal place_390_preds : BooleanArray(0 downto 0);
  signal place_390_succs : BooleanArray(0 downto 0);
  signal place_390_token : boolean;
  signal place_395_preds : BooleanArray(0 downto 0);
  signal place_395_succs : BooleanArray(0 downto 0);
  signal place_395_token : boolean;
  signal place_396_preds : BooleanArray(0 downto 0);
  signal place_396_succs : BooleanArray(0 downto 0);
  signal place_396_token : boolean;
  signal place_397_preds : BooleanArray(0 downto 0);
  signal place_397_succs : BooleanArray(0 downto 0);
  signal place_397_token : boolean;
  signal place_402_preds : BooleanArray(0 downto 0);
  signal place_402_succs : BooleanArray(0 downto 0);
  signal place_402_token : boolean;
  signal place_403_preds : BooleanArray(0 downto 0);
  signal place_403_succs : BooleanArray(0 downto 0);
  signal place_403_token : boolean;
  signal place_404_preds : BooleanArray(0 downto 0);
  signal place_404_succs : BooleanArray(0 downto 0);
  signal place_404_token : boolean;
  signal place_410_preds : BooleanArray(0 downto 0);
  signal place_410_succs : BooleanArray(0 downto 0);
  signal place_410_token : boolean;
  signal place_411_preds : BooleanArray(0 downto 0);
  signal place_411_succs : BooleanArray(0 downto 0);
  signal place_411_token : boolean;
  signal place_412_preds : BooleanArray(0 downto 0);
  signal place_412_succs : BooleanArray(0 downto 0);
  signal place_412_token : boolean;
  signal place_417_preds : BooleanArray(0 downto 0);
  signal place_417_succs : BooleanArray(0 downto 0);
  signal place_417_token : boolean;
  signal place_418_preds : BooleanArray(0 downto 0);
  signal place_418_succs : BooleanArray(0 downto 0);
  signal place_418_token : boolean;
  signal place_419_preds : BooleanArray(0 downto 0);
  signal place_419_succs : BooleanArray(0 downto 0);
  signal place_419_token : boolean;
  signal place_424_preds : BooleanArray(0 downto 0);
  signal place_424_succs : BooleanArray(0 downto 0);
  signal place_424_token : boolean;
  signal place_425_preds : BooleanArray(0 downto 0);
  signal place_425_succs : BooleanArray(0 downto 0);
  signal place_425_token : boolean;
  signal place_426_preds : BooleanArray(0 downto 0);
  signal place_426_succs : BooleanArray(0 downto 0);
  signal place_426_token : boolean;
  signal place_432_preds : BooleanArray(0 downto 0);
  signal place_432_succs : BooleanArray(0 downto 0);
  signal place_432_token : boolean;
  signal place_433_preds : BooleanArray(0 downto 0);
  signal place_433_succs : BooleanArray(0 downto 0);
  signal place_433_token : boolean;
  signal place_434_preds : BooleanArray(0 downto 0);
  signal place_434_succs : BooleanArray(0 downto 0);
  signal place_434_token : boolean;
  signal place_435_preds : BooleanArray(0 downto 0);
  signal place_435_succs : BooleanArray(0 downto 0);
  signal place_435_token : boolean;
  signal place_443_preds : BooleanArray(0 downto 0);
  signal place_443_succs : BooleanArray(0 downto 0);
  signal place_443_token : boolean;
  signal place_444_preds : BooleanArray(0 downto 0);
  signal place_444_succs : BooleanArray(0 downto 0);
  signal place_444_token : boolean;
  signal place_445_preds : BooleanArray(0 downto 0);
  signal place_445_succs : BooleanArray(0 downto 0);
  signal place_445_token : boolean;
  signal place_450_preds : BooleanArray(0 downto 0);
  signal place_450_succs : BooleanArray(0 downto 0);
  signal place_450_token : boolean;
  signal place_451_preds : BooleanArray(0 downto 0);
  signal place_451_succs : BooleanArray(0 downto 0);
  signal place_451_token : boolean;
  signal place_452_preds : BooleanArray(0 downto 0);
  signal place_452_succs : BooleanArray(0 downto 0);
  signal place_452_token : boolean;
  signal place_457_preds : BooleanArray(0 downto 0);
  signal place_457_succs : BooleanArray(0 downto 0);
  signal place_457_token : boolean;
  signal place_458_preds : BooleanArray(0 downto 0);
  signal place_458_succs : BooleanArray(0 downto 0);
  signal place_458_token : boolean;
  signal place_459_preds : BooleanArray(0 downto 0);
  signal place_459_succs : BooleanArray(0 downto 0);
  signal place_459_token : boolean;
  signal place_464_preds : BooleanArray(0 downto 0);
  signal place_464_succs : BooleanArray(0 downto 0);
  signal place_464_token : boolean;
  signal place_465_preds : BooleanArray(0 downto 0);
  signal place_465_succs : BooleanArray(0 downto 0);
  signal place_465_token : boolean;
  signal place_466_preds : BooleanArray(0 downto 0);
  signal place_466_succs : BooleanArray(0 downto 0);
  signal place_466_token : boolean;
  signal place_471_preds : BooleanArray(0 downto 0);
  signal place_471_succs : BooleanArray(0 downto 0);
  signal place_471_token : boolean;
  signal place_472_preds : BooleanArray(0 downto 0);
  signal place_472_succs : BooleanArray(0 downto 0);
  signal place_472_token : boolean;
  signal place_473_preds : BooleanArray(0 downto 0);
  signal place_473_succs : BooleanArray(0 downto 0);
  signal place_473_token : boolean;
  signal place_479_preds : BooleanArray(0 downto 0);
  signal place_479_succs : BooleanArray(0 downto 0);
  signal place_479_token : boolean;
  signal place_480_preds : BooleanArray(0 downto 0);
  signal place_480_succs : BooleanArray(0 downto 0);
  signal place_480_token : boolean;
  signal place_481_preds : BooleanArray(0 downto 0);
  signal place_481_succs : BooleanArray(0 downto 0);
  signal place_481_token : boolean;
  signal place_486_preds : BooleanArray(0 downto 0);
  signal place_486_succs : BooleanArray(0 downto 0);
  signal place_486_token : boolean;
  signal place_487_preds : BooleanArray(0 downto 0);
  signal place_487_succs : BooleanArray(0 downto 0);
  signal place_487_token : boolean;
  signal place_488_preds : BooleanArray(0 downto 0);
  signal place_488_succs : BooleanArray(0 downto 0);
  signal place_488_token : boolean;
  signal place_494_preds : BooleanArray(0 downto 0);
  signal place_494_succs : BooleanArray(0 downto 0);
  signal place_494_token : boolean;
  signal place_495_preds : BooleanArray(0 downto 0);
  signal place_495_succs : BooleanArray(0 downto 0);
  signal place_495_token : boolean;
  signal place_496_preds : BooleanArray(0 downto 0);
  signal place_496_succs : BooleanArray(0 downto 0);
  signal place_496_token : boolean;
  signal place_497_preds : BooleanArray(0 downto 0);
  signal place_497_succs : BooleanArray(0 downto 0);
  signal place_497_token : boolean;
  signal place_505_preds : BooleanArray(0 downto 0);
  signal place_505_succs : BooleanArray(0 downto 0);
  signal place_505_token : boolean;
  signal place_506_preds : BooleanArray(0 downto 0);
  signal place_506_succs : BooleanArray(0 downto 0);
  signal place_506_token : boolean;
  signal place_507_preds : BooleanArray(0 downto 0);
  signal place_507_succs : BooleanArray(0 downto 0);
  signal place_507_token : boolean;
  signal place_512_preds : BooleanArray(0 downto 0);
  signal place_512_succs : BooleanArray(0 downto 0);
  signal place_512_token : boolean;
  signal place_513_preds : BooleanArray(0 downto 0);
  signal place_513_succs : BooleanArray(0 downto 0);
  signal place_513_token : boolean;
  signal place_514_preds : BooleanArray(0 downto 0);
  signal place_514_succs : BooleanArray(0 downto 0);
  signal place_514_token : boolean;
  signal place_519_preds : BooleanArray(0 downto 0);
  signal place_519_succs : BooleanArray(0 downto 0);
  signal place_519_token : boolean;
  signal place_520_preds : BooleanArray(0 downto 0);
  signal place_520_succs : BooleanArray(0 downto 0);
  signal place_520_token : boolean;
  signal place_521_preds : BooleanArray(0 downto 0);
  signal place_521_succs : BooleanArray(0 downto 0);
  signal place_521_token : boolean;
  signal place_527_preds : BooleanArray(0 downto 0);
  signal place_527_succs : BooleanArray(0 downto 0);
  signal place_527_token : boolean;
  signal place_528_preds : BooleanArray(0 downto 0);
  signal place_528_succs : BooleanArray(0 downto 0);
  signal place_528_token : boolean;
  signal place_529_preds : BooleanArray(0 downto 0);
  signal place_529_succs : BooleanArray(0 downto 0);
  signal place_529_token : boolean;
  signal place_534_preds : BooleanArray(0 downto 0);
  signal place_534_succs : BooleanArray(0 downto 0);
  signal place_534_token : boolean;
  signal place_535_preds : BooleanArray(0 downto 0);
  signal place_535_succs : BooleanArray(0 downto 0);
  signal place_535_token : boolean;
  signal place_536_preds : BooleanArray(0 downto 0);
  signal place_536_succs : BooleanArray(0 downto 0);
  signal place_536_token : boolean;
  signal place_542_preds : BooleanArray(0 downto 0);
  signal place_542_succs : BooleanArray(0 downto 0);
  signal place_542_token : boolean;
  signal place_543_preds : BooleanArray(0 downto 0);
  signal place_543_succs : BooleanArray(0 downto 0);
  signal place_543_token : boolean;
  signal place_544_preds : BooleanArray(0 downto 0);
  signal place_544_succs : BooleanArray(0 downto 0);
  signal place_544_token : boolean;
  signal place_545_preds : BooleanArray(0 downto 0);
  signal place_545_succs : BooleanArray(0 downto 0);
  signal place_545_token : boolean;
  signal place_553_preds : BooleanArray(0 downto 0);
  signal place_553_succs : BooleanArray(0 downto 0);
  signal place_553_token : boolean;
  signal place_554_preds : BooleanArray(0 downto 0);
  signal place_554_succs : BooleanArray(0 downto 0);
  signal place_554_token : boolean;
  signal place_555_preds : BooleanArray(0 downto 0);
  signal place_555_succs : BooleanArray(0 downto 0);
  signal place_555_token : boolean;
  signal place_560_preds : BooleanArray(0 downto 0);
  signal place_560_succs : BooleanArray(0 downto 0);
  signal place_560_token : boolean;
  signal place_561_preds : BooleanArray(0 downto 0);
  signal place_561_succs : BooleanArray(0 downto 0);
  signal place_561_token : boolean;
  signal place_562_preds : BooleanArray(0 downto 0);
  signal place_562_succs : BooleanArray(0 downto 0);
  signal place_562_token : boolean;
  signal place_567_preds : BooleanArray(0 downto 0);
  signal place_567_succs : BooleanArray(0 downto 0);
  signal place_567_token : boolean;
  signal place_568_preds : BooleanArray(0 downto 0);
  signal place_568_succs : BooleanArray(0 downto 0);
  signal place_568_token : boolean;
  signal place_569_preds : BooleanArray(0 downto 0);
  signal place_569_succs : BooleanArray(0 downto 0);
  signal place_569_token : boolean;
  signal place_575_preds : BooleanArray(0 downto 0);
  signal place_575_succs : BooleanArray(0 downto 0);
  signal place_575_token : boolean;
  signal place_576_preds : BooleanArray(0 downto 0);
  signal place_576_succs : BooleanArray(0 downto 0);
  signal place_576_token : boolean;
  signal place_577_preds : BooleanArray(0 downto 0);
  signal place_577_succs : BooleanArray(0 downto 0);
  signal place_577_token : boolean;
  signal place_582_preds : BooleanArray(0 downto 0);
  signal place_582_succs : BooleanArray(0 downto 0);
  signal place_582_token : boolean;
  signal place_583_preds : BooleanArray(0 downto 0);
  signal place_583_succs : BooleanArray(0 downto 0);
  signal place_583_token : boolean;
  signal place_584_preds : BooleanArray(0 downto 0);
  signal place_584_succs : BooleanArray(0 downto 0);
  signal place_584_token : boolean;
  signal place_590_preds : BooleanArray(0 downto 0);
  signal place_590_succs : BooleanArray(0 downto 0);
  signal place_590_token : boolean;
  signal place_591_preds : BooleanArray(0 downto 0);
  signal place_591_succs : BooleanArray(0 downto 0);
  signal place_591_token : boolean;
  signal place_592_preds : BooleanArray(0 downto 0);
  signal place_592_succs : BooleanArray(0 downto 0);
  signal place_592_token : boolean;
  signal place_593_preds : BooleanArray(0 downto 0);
  signal place_593_succs : BooleanArray(0 downto 0);
  signal place_593_token : boolean;
  signal place_601_preds : BooleanArray(0 downto 0);
  signal place_601_succs : BooleanArray(0 downto 0);
  signal place_601_token : boolean;
  signal place_602_preds : BooleanArray(0 downto 0);
  signal place_602_succs : BooleanArray(0 downto 0);
  signal place_602_token : boolean;
  signal place_603_preds : BooleanArray(0 downto 0);
  signal place_603_succs : BooleanArray(0 downto 0);
  signal place_603_token : boolean;
  signal place_608_preds : BooleanArray(0 downto 0);
  signal place_608_succs : BooleanArray(0 downto 0);
  signal place_608_token : boolean;
  signal place_609_preds : BooleanArray(0 downto 0);
  signal place_609_succs : BooleanArray(0 downto 0);
  signal place_609_token : boolean;
  signal place_610_preds : BooleanArray(0 downto 0);
  signal place_610_succs : BooleanArray(0 downto 0);
  signal place_610_token : boolean;
  signal place_615_preds : BooleanArray(0 downto 0);
  signal place_615_succs : BooleanArray(0 downto 0);
  signal place_615_token : boolean;
  signal place_616_preds : BooleanArray(0 downto 0);
  signal place_616_succs : BooleanArray(0 downto 0);
  signal place_616_token : boolean;
  signal place_617_preds : BooleanArray(0 downto 0);
  signal place_617_succs : BooleanArray(0 downto 0);
  signal place_617_token : boolean;
  signal place_623_preds : BooleanArray(0 downto 0);
  signal place_623_succs : BooleanArray(0 downto 0);
  signal place_623_token : boolean;
  signal place_624_preds : BooleanArray(0 downto 0);
  signal place_624_succs : BooleanArray(0 downto 0);
  signal place_624_token : boolean;
  signal place_625_preds : BooleanArray(0 downto 0);
  signal place_625_succs : BooleanArray(0 downto 0);
  signal place_625_token : boolean;
  signal place_630_preds : BooleanArray(0 downto 0);
  signal place_630_succs : BooleanArray(0 downto 0);
  signal place_630_token : boolean;
  signal place_631_preds : BooleanArray(0 downto 0);
  signal place_631_succs : BooleanArray(0 downto 0);
  signal place_631_token : boolean;
  signal place_632_preds : BooleanArray(0 downto 0);
  signal place_632_succs : BooleanArray(0 downto 0);
  signal place_632_token : boolean;
  signal place_638_preds : BooleanArray(0 downto 0);
  signal place_638_succs : BooleanArray(0 downto 0);
  signal place_638_token : boolean;
  signal place_639_preds : BooleanArray(0 downto 0);
  signal place_639_succs : BooleanArray(0 downto 0);
  signal place_639_token : boolean;
  signal place_640_preds : BooleanArray(0 downto 0);
  signal place_640_succs : BooleanArray(0 downto 0);
  signal place_640_token : boolean;
  signal place_641_preds : BooleanArray(0 downto 0);
  signal place_641_succs : BooleanArray(0 downto 0);
  signal place_641_token : boolean;
  signal place_649_preds : BooleanArray(0 downto 0);
  signal place_649_succs : BooleanArray(0 downto 0);
  signal place_649_token : boolean;
  signal place_650_preds : BooleanArray(0 downto 0);
  signal place_650_succs : BooleanArray(0 downto 0);
  signal place_650_token : boolean;
  signal place_651_preds : BooleanArray(0 downto 0);
  signal place_651_succs : BooleanArray(0 downto 0);
  signal place_651_token : boolean;
  signal place_656_preds : BooleanArray(0 downto 0);
  signal place_656_succs : BooleanArray(0 downto 0);
  signal place_656_token : boolean;
  signal place_657_preds : BooleanArray(0 downto 0);
  signal place_657_succs : BooleanArray(0 downto 0);
  signal place_657_token : boolean;
  signal place_658_preds : BooleanArray(0 downto 0);
  signal place_658_succs : BooleanArray(0 downto 0);
  signal place_658_token : boolean;
  signal place_663_preds : BooleanArray(0 downto 0);
  signal place_663_succs : BooleanArray(0 downto 0);
  signal place_663_token : boolean;
  signal place_664_preds : BooleanArray(0 downto 0);
  signal place_664_succs : BooleanArray(0 downto 0);
  signal place_664_token : boolean;
  signal place_665_preds : BooleanArray(0 downto 0);
  signal place_665_succs : BooleanArray(0 downto 0);
  signal place_665_token : boolean;
  signal place_671_preds : BooleanArray(0 downto 0);
  signal place_671_succs : BooleanArray(0 downto 0);
  signal place_671_token : boolean;
  signal place_672_preds : BooleanArray(0 downto 0);
  signal place_672_succs : BooleanArray(0 downto 0);
  signal place_672_token : boolean;
  signal place_673_preds : BooleanArray(0 downto 0);
  signal place_673_succs : BooleanArray(0 downto 0);
  signal place_673_token : boolean;
  signal place_678_preds : BooleanArray(0 downto 0);
  signal place_678_succs : BooleanArray(0 downto 0);
  signal place_678_token : boolean;
  signal place_679_preds : BooleanArray(0 downto 0);
  signal place_679_succs : BooleanArray(0 downto 0);
  signal place_679_token : boolean;
  signal place_680_preds : BooleanArray(0 downto 0);
  signal place_680_succs : BooleanArray(0 downto 0);
  signal place_680_token : boolean;
  signal place_686_preds : BooleanArray(0 downto 0);
  signal place_686_succs : BooleanArray(0 downto 0);
  signal place_686_token : boolean;
  signal place_687_preds : BooleanArray(0 downto 0);
  signal place_687_succs : BooleanArray(0 downto 0);
  signal place_687_token : boolean;
  signal place_688_preds : BooleanArray(0 downto 0);
  signal place_688_succs : BooleanArray(0 downto 0);
  signal place_688_token : boolean;
  signal place_689_preds : BooleanArray(0 downto 0);
  signal place_689_succs : BooleanArray(0 downto 0);
  signal place_689_token : boolean;
  signal place_697_preds : BooleanArray(0 downto 0);
  signal place_697_succs : BooleanArray(0 downto 0);
  signal place_697_token : boolean;
  signal place_698_preds : BooleanArray(0 downto 0);
  signal place_698_succs : BooleanArray(0 downto 0);
  signal place_698_token : boolean;
  signal place_699_preds : BooleanArray(0 downto 0);
  signal place_699_succs : BooleanArray(0 downto 0);
  signal place_699_token : boolean;
  signal place_704_preds : BooleanArray(0 downto 0);
  signal place_704_succs : BooleanArray(0 downto 0);
  signal place_704_token : boolean;
  signal place_705_preds : BooleanArray(0 downto 0);
  signal place_705_succs : BooleanArray(0 downto 0);
  signal place_705_token : boolean;
  signal place_706_preds : BooleanArray(0 downto 0);
  signal place_706_succs : BooleanArray(0 downto 0);
  signal place_706_token : boolean;
  signal place_711_preds : BooleanArray(0 downto 0);
  signal place_711_succs : BooleanArray(0 downto 0);
  signal place_711_token : boolean;
  signal place_712_preds : BooleanArray(0 downto 0);
  signal place_712_succs : BooleanArray(0 downto 0);
  signal place_712_token : boolean;
  signal place_713_preds : BooleanArray(0 downto 0);
  signal place_713_succs : BooleanArray(0 downto 0);
  signal place_713_token : boolean;
  signal place_719_preds : BooleanArray(0 downto 0);
  signal place_719_succs : BooleanArray(0 downto 0);
  signal place_719_token : boolean;
  signal place_720_preds : BooleanArray(0 downto 0);
  signal place_720_succs : BooleanArray(0 downto 0);
  signal place_720_token : boolean;
  signal place_721_preds : BooleanArray(0 downto 0);
  signal place_721_succs : BooleanArray(0 downto 0);
  signal place_721_token : boolean;
  signal place_726_preds : BooleanArray(0 downto 0);
  signal place_726_succs : BooleanArray(0 downto 0);
  signal place_726_token : boolean;
  signal place_727_preds : BooleanArray(0 downto 0);
  signal place_727_succs : BooleanArray(0 downto 0);
  signal place_727_token : boolean;
  signal place_728_preds : BooleanArray(0 downto 0);
  signal place_728_succs : BooleanArray(0 downto 0);
  signal place_728_token : boolean;
  signal place_734_preds : BooleanArray(0 downto 0);
  signal place_734_succs : BooleanArray(0 downto 0);
  signal place_734_token : boolean;
  signal place_735_preds : BooleanArray(0 downto 0);
  signal place_735_succs : BooleanArray(0 downto 0);
  signal place_735_token : boolean;
  signal place_736_preds : BooleanArray(0 downto 0);
  signal place_736_succs : BooleanArray(0 downto 0);
  signal place_736_token : boolean;
  signal place_737_preds : BooleanArray(0 downto 0);
  signal place_737_succs : BooleanArray(0 downto 0);
  signal place_737_token : boolean;
  signal place_745_preds : BooleanArray(0 downto 0);
  signal place_745_succs : BooleanArray(0 downto 0);
  signal place_745_token : boolean;
  signal place_746_preds : BooleanArray(0 downto 0);
  signal place_746_succs : BooleanArray(0 downto 0);
  signal place_746_token : boolean;
  signal place_747_preds : BooleanArray(0 downto 0);
  signal place_747_succs : BooleanArray(0 downto 0);
  signal place_747_token : boolean;
  signal place_752_preds : BooleanArray(0 downto 0);
  signal place_752_succs : BooleanArray(0 downto 0);
  signal place_752_token : boolean;
  signal place_753_preds : BooleanArray(0 downto 0);
  signal place_753_succs : BooleanArray(0 downto 0);
  signal place_753_token : boolean;
  signal place_754_preds : BooleanArray(0 downto 0);
  signal place_754_succs : BooleanArray(0 downto 0);
  signal place_754_token : boolean;
  signal place_759_preds : BooleanArray(0 downto 0);
  signal place_759_succs : BooleanArray(0 downto 0);
  signal place_759_token : boolean;
  signal place_760_preds : BooleanArray(0 downto 0);
  signal place_760_succs : BooleanArray(0 downto 0);
  signal place_760_token : boolean;
  signal place_761_preds : BooleanArray(0 downto 0);
  signal place_761_succs : BooleanArray(0 downto 0);
  signal place_761_token : boolean;
  signal place_767_preds : BooleanArray(0 downto 0);
  signal place_767_succs : BooleanArray(0 downto 0);
  signal place_767_token : boolean;
  signal place_768_preds : BooleanArray(0 downto 0);
  signal place_768_succs : BooleanArray(0 downto 0);
  signal place_768_token : boolean;
  signal place_769_preds : BooleanArray(0 downto 0);
  signal place_769_succs : BooleanArray(0 downto 0);
  signal place_769_token : boolean;
  signal place_774_preds : BooleanArray(0 downto 0);
  signal place_774_succs : BooleanArray(0 downto 0);
  signal place_774_token : boolean;
  signal place_775_preds : BooleanArray(0 downto 0);
  signal place_775_succs : BooleanArray(0 downto 0);
  signal place_775_token : boolean;
  signal place_776_preds : BooleanArray(0 downto 0);
  signal place_776_succs : BooleanArray(0 downto 0);
  signal place_776_token : boolean;
  signal place_782_preds : BooleanArray(0 downto 0);
  signal place_782_succs : BooleanArray(0 downto 0);
  signal place_782_token : boolean;
  signal place_783_preds : BooleanArray(0 downto 0);
  signal place_783_succs : BooleanArray(0 downto 0);
  signal place_783_token : boolean;
  signal place_784_preds : BooleanArray(0 downto 0);
  signal place_784_succs : BooleanArray(0 downto 0);
  signal place_784_token : boolean;
  signal place_785_preds : BooleanArray(0 downto 0);
  signal place_785_succs : BooleanArray(0 downto 0);
  signal place_785_token : boolean;
  signal place_793_preds : BooleanArray(0 downto 0);
  signal place_793_succs : BooleanArray(0 downto 0);
  signal place_793_token : boolean;
  signal place_794_preds : BooleanArray(0 downto 0);
  signal place_794_succs : BooleanArray(0 downto 0);
  signal place_794_token : boolean;
  signal place_795_preds : BooleanArray(0 downto 0);
  signal place_795_succs : BooleanArray(0 downto 0);
  signal place_795_token : boolean;
  signal place_800_preds : BooleanArray(0 downto 0);
  signal place_800_succs : BooleanArray(0 downto 0);
  signal place_800_token : boolean;
  signal place_801_preds : BooleanArray(0 downto 0);
  signal place_801_succs : BooleanArray(0 downto 0);
  signal place_801_token : boolean;
  signal place_802_preds : BooleanArray(0 downto 0);
  signal place_802_succs : BooleanArray(0 downto 0);
  signal place_802_token : boolean;
  signal place_807_preds : BooleanArray(0 downto 0);
  signal place_807_succs : BooleanArray(0 downto 0);
  signal place_807_token : boolean;
  signal place_808_preds : BooleanArray(0 downto 0);
  signal place_808_succs : BooleanArray(0 downto 0);
  signal place_808_token : boolean;
  signal place_809_preds : BooleanArray(0 downto 0);
  signal place_809_succs : BooleanArray(0 downto 0);
  signal place_809_token : boolean;
  signal place_815_preds : BooleanArray(0 downto 0);
  signal place_815_succs : BooleanArray(0 downto 0);
  signal place_815_token : boolean;
  signal place_816_preds : BooleanArray(0 downto 0);
  signal place_816_succs : BooleanArray(0 downto 0);
  signal place_816_token : boolean;
  signal place_817_preds : BooleanArray(0 downto 0);
  signal place_817_succs : BooleanArray(0 downto 0);
  signal place_817_token : boolean;
  signal place_822_preds : BooleanArray(0 downto 0);
  signal place_822_succs : BooleanArray(0 downto 0);
  signal place_822_token : boolean;
  signal place_823_preds : BooleanArray(0 downto 0);
  signal place_823_succs : BooleanArray(0 downto 0);
  signal place_823_token : boolean;
  signal place_824_preds : BooleanArray(0 downto 0);
  signal place_824_succs : BooleanArray(0 downto 0);
  signal place_824_token : boolean;
  signal place_830_preds : BooleanArray(0 downto 0);
  signal place_830_succs : BooleanArray(0 downto 0);
  signal place_830_token : boolean;
  signal place_831_preds : BooleanArray(0 downto 0);
  signal place_831_succs : BooleanArray(0 downto 0);
  signal place_831_token : boolean;
  signal place_832_preds : BooleanArray(0 downto 0);
  signal place_832_succs : BooleanArray(0 downto 0);
  signal place_832_token : boolean;
  signal place_833_preds : BooleanArray(0 downto 0);
  signal place_833_succs : BooleanArray(0 downto 0);
  signal place_833_token : boolean;
  signal place_841_preds : BooleanArray(0 downto 0);
  signal place_841_succs : BooleanArray(0 downto 0);
  signal place_841_token : boolean;
  signal place_842_preds : BooleanArray(0 downto 0);
  signal place_842_succs : BooleanArray(0 downto 0);
  signal place_842_token : boolean;
  signal place_843_preds : BooleanArray(0 downto 0);
  signal place_843_succs : BooleanArray(0 downto 0);
  signal place_843_token : boolean;
  signal place_848_preds : BooleanArray(0 downto 0);
  signal place_848_succs : BooleanArray(0 downto 0);
  signal place_848_token : boolean;
  signal place_849_preds : BooleanArray(0 downto 0);
  signal place_849_succs : BooleanArray(0 downto 0);
  signal place_849_token : boolean;
  signal place_850_preds : BooleanArray(0 downto 0);
  signal place_850_succs : BooleanArray(0 downto 0);
  signal place_850_token : boolean;
  signal place_855_preds : BooleanArray(0 downto 0);
  signal place_855_succs : BooleanArray(0 downto 0);
  signal place_855_token : boolean;
  signal place_856_preds : BooleanArray(0 downto 0);
  signal place_856_succs : BooleanArray(0 downto 0);
  signal place_856_token : boolean;
  signal place_857_preds : BooleanArray(0 downto 0);
  signal place_857_succs : BooleanArray(0 downto 0);
  signal place_857_token : boolean;
  signal place_863_preds : BooleanArray(0 downto 0);
  signal place_863_succs : BooleanArray(0 downto 0);
  signal place_863_token : boolean;
  signal place_864_preds : BooleanArray(0 downto 0);
  signal place_864_succs : BooleanArray(0 downto 0);
  signal place_864_token : boolean;
  signal place_865_preds : BooleanArray(0 downto 0);
  signal place_865_succs : BooleanArray(0 downto 0);
  signal place_865_token : boolean;
  signal place_870_preds : BooleanArray(0 downto 0);
  signal place_870_succs : BooleanArray(0 downto 0);
  signal place_870_token : boolean;
  signal place_871_preds : BooleanArray(0 downto 0);
  signal place_871_succs : BooleanArray(0 downto 0);
  signal place_871_token : boolean;
  signal place_872_preds : BooleanArray(0 downto 0);
  signal place_872_succs : BooleanArray(0 downto 0);
  signal place_872_token : boolean;
  signal place_878_preds : BooleanArray(0 downto 0);
  signal place_878_succs : BooleanArray(0 downto 0);
  signal place_878_token : boolean;
  signal place_879_preds : BooleanArray(0 downto 0);
  signal place_879_succs : BooleanArray(0 downto 0);
  signal place_879_token : boolean;
  signal place_880_preds : BooleanArray(0 downto 0);
  signal place_880_succs : BooleanArray(0 downto 0);
  signal place_880_token : boolean;
  signal place_881_preds : BooleanArray(0 downto 0);
  signal place_881_succs : BooleanArray(0 downto 0);
  signal place_881_token : boolean;
  signal place_889_preds : BooleanArray(0 downto 0);
  signal place_889_succs : BooleanArray(0 downto 0);
  signal place_889_token : boolean;
  signal place_890_preds : BooleanArray(0 downto 0);
  signal place_890_succs : BooleanArray(0 downto 0);
  signal place_890_token : boolean;
  signal place_891_preds : BooleanArray(0 downto 0);
  signal place_891_succs : BooleanArray(0 downto 0);
  signal place_891_token : boolean;
  signal place_896_preds : BooleanArray(0 downto 0);
  signal place_896_succs : BooleanArray(0 downto 0);
  signal place_896_token : boolean;
  signal place_897_preds : BooleanArray(0 downto 0);
  signal place_897_succs : BooleanArray(0 downto 0);
  signal place_897_token : boolean;
  signal place_898_preds : BooleanArray(0 downto 0);
  signal place_898_succs : BooleanArray(0 downto 0);
  signal place_898_token : boolean;
  signal place_903_preds : BooleanArray(0 downto 0);
  signal place_903_succs : BooleanArray(0 downto 0);
  signal place_903_token : boolean;
  signal place_904_preds : BooleanArray(0 downto 0);
  signal place_904_succs : BooleanArray(0 downto 0);
  signal place_904_token : boolean;
  signal place_905_preds : BooleanArray(0 downto 0);
  signal place_905_succs : BooleanArray(0 downto 0);
  signal place_905_token : boolean;
  signal place_911_preds : BooleanArray(0 downto 0);
  signal place_911_succs : BooleanArray(0 downto 0);
  signal place_911_token : boolean;
  signal place_912_preds : BooleanArray(0 downto 0);
  signal place_912_succs : BooleanArray(0 downto 0);
  signal place_912_token : boolean;
  signal place_913_preds : BooleanArray(0 downto 0);
  signal place_913_succs : BooleanArray(0 downto 0);
  signal place_913_token : boolean;
  signal place_918_preds : BooleanArray(0 downto 0);
  signal place_918_succs : BooleanArray(0 downto 0);
  signal place_918_token : boolean;
  signal place_919_preds : BooleanArray(0 downto 0);
  signal place_919_succs : BooleanArray(0 downto 0);
  signal place_919_token : boolean;
  signal place_920_preds : BooleanArray(0 downto 0);
  signal place_920_succs : BooleanArray(0 downto 0);
  signal place_920_token : boolean;
  signal place_926_preds : BooleanArray(0 downto 0);
  signal place_926_succs : BooleanArray(0 downto 0);
  signal place_926_token : boolean;
  signal place_927_preds : BooleanArray(0 downto 0);
  signal place_927_succs : BooleanArray(0 downto 0);
  signal place_927_token : boolean;
  signal place_928_preds : BooleanArray(0 downto 0);
  signal place_928_succs : BooleanArray(0 downto 0);
  signal place_928_token : boolean;
  signal place_929_preds : BooleanArray(0 downto 0);
  signal place_929_succs : BooleanArray(0 downto 0);
  signal place_929_token : boolean;
  signal place_937_preds : BooleanArray(0 downto 0);
  signal place_937_succs : BooleanArray(0 downto 0);
  signal place_937_token : boolean;
  signal place_938_preds : BooleanArray(0 downto 0);
  signal place_938_succs : BooleanArray(0 downto 0);
  signal place_938_token : boolean;
  signal place_939_preds : BooleanArray(0 downto 0);
  signal place_939_succs : BooleanArray(0 downto 0);
  signal place_939_token : boolean;
  signal place_944_preds : BooleanArray(0 downto 0);
  signal place_944_succs : BooleanArray(0 downto 0);
  signal place_944_token : boolean;
  signal place_945_preds : BooleanArray(0 downto 0);
  signal place_945_succs : BooleanArray(0 downto 0);
  signal place_945_token : boolean;
  signal place_946_preds : BooleanArray(0 downto 0);
  signal place_946_succs : BooleanArray(0 downto 0);
  signal place_946_token : boolean;
  signal place_951_preds : BooleanArray(0 downto 0);
  signal place_951_succs : BooleanArray(0 downto 0);
  signal place_951_token : boolean;
  signal place_952_preds : BooleanArray(0 downto 0);
  signal place_952_succs : BooleanArray(0 downto 0);
  signal place_952_token : boolean;
  signal place_953_preds : BooleanArray(0 downto 0);
  signal place_953_succs : BooleanArray(0 downto 0);
  signal place_953_token : boolean;
  signal place_959_preds : BooleanArray(0 downto 0);
  signal place_959_succs : BooleanArray(0 downto 0);
  signal place_959_token : boolean;
  signal place_960_preds : BooleanArray(0 downto 0);
  signal place_960_succs : BooleanArray(0 downto 0);
  signal place_960_token : boolean;
  signal place_961_preds : BooleanArray(0 downto 0);
  signal place_961_succs : BooleanArray(0 downto 0);
  signal place_961_token : boolean;
  signal place_966_preds : BooleanArray(0 downto 0);
  signal place_966_succs : BooleanArray(0 downto 0);
  signal place_966_token : boolean;
  signal place_967_preds : BooleanArray(0 downto 0);
  signal place_967_succs : BooleanArray(0 downto 0);
  signal place_967_token : boolean;
  signal place_968_preds : BooleanArray(0 downto 0);
  signal place_968_succs : BooleanArray(0 downto 0);
  signal place_968_token : boolean;
  signal place_974_preds : BooleanArray(0 downto 0);
  signal place_974_succs : BooleanArray(0 downto 0);
  signal place_974_token : boolean;
  signal place_975_preds : BooleanArray(0 downto 0);
  signal place_975_succs : BooleanArray(0 downto 0);
  signal place_975_token : boolean;
  signal place_976_preds : BooleanArray(0 downto 0);
  signal place_976_succs : BooleanArray(0 downto 0);
  signal place_976_token : boolean;
  signal place_977_preds : BooleanArray(0 downto 0);
  signal place_977_succs : BooleanArray(0 downto 0);
  signal place_977_token : boolean;
  signal place_985_preds : BooleanArray(0 downto 0);
  signal place_985_succs : BooleanArray(0 downto 0);
  signal place_985_token : boolean;
  signal place_986_preds : BooleanArray(0 downto 0);
  signal place_986_succs : BooleanArray(0 downto 0);
  signal place_986_token : boolean;
  signal place_987_preds : BooleanArray(0 downto 0);
  signal place_987_succs : BooleanArray(0 downto 0);
  signal place_987_token : boolean;
  signal place_992_preds : BooleanArray(0 downto 0);
  signal place_992_succs : BooleanArray(0 downto 0);
  signal place_992_token : boolean;
  signal place_993_preds : BooleanArray(0 downto 0);
  signal place_993_succs : BooleanArray(0 downto 0);
  signal place_993_token : boolean;
  signal place_994_preds : BooleanArray(0 downto 0);
  signal place_994_succs : BooleanArray(0 downto 0);
  signal place_994_token : boolean;
  signal place_999_preds : BooleanArray(0 downto 0);
  signal place_999_succs : BooleanArray(0 downto 0);
  signal place_999_token : boolean;
  signal place_1000_preds : BooleanArray(0 downto 0);
  signal place_1000_succs : BooleanArray(0 downto 0);
  signal place_1000_token : boolean;
  signal place_1001_preds : BooleanArray(0 downto 0);
  signal place_1001_succs : BooleanArray(0 downto 0);
  signal place_1001_token : boolean;
  signal place_1007_preds : BooleanArray(0 downto 0);
  signal place_1007_succs : BooleanArray(0 downto 0);
  signal place_1007_token : boolean;
  signal place_1008_preds : BooleanArray(0 downto 0);
  signal place_1008_succs : BooleanArray(0 downto 0);
  signal place_1008_token : boolean;
  signal place_1009_preds : BooleanArray(0 downto 0);
  signal place_1009_succs : BooleanArray(0 downto 0);
  signal place_1009_token : boolean;
  signal place_1014_preds : BooleanArray(0 downto 0);
  signal place_1014_succs : BooleanArray(0 downto 0);
  signal place_1014_token : boolean;
  signal place_1015_preds : BooleanArray(0 downto 0);
  signal place_1015_succs : BooleanArray(0 downto 0);
  signal place_1015_token : boolean;
  signal place_1016_preds : BooleanArray(0 downto 0);
  signal place_1016_succs : BooleanArray(0 downto 0);
  signal place_1016_token : boolean;
  signal place_1022_preds : BooleanArray(0 downto 0);
  signal place_1022_succs : BooleanArray(0 downto 0);
  signal place_1022_token : boolean;
  signal place_1023_preds : BooleanArray(0 downto 0);
  signal place_1023_succs : BooleanArray(0 downto 0);
  signal place_1023_token : boolean;
  signal place_1024_preds : BooleanArray(0 downto 0);
  signal place_1024_succs : BooleanArray(0 downto 0);
  signal place_1024_token : boolean;
  signal place_1025_preds : BooleanArray(0 downto 0);
  signal place_1025_succs : BooleanArray(0 downto 0);
  signal place_1025_token : boolean;
  signal place_1029_preds : BooleanArray(0 downto 0);
  signal place_1029_succs : BooleanArray(0 downto 0);
  signal place_1029_token : boolean;
  signal place_1032_preds : BooleanArray(0 downto 0);
  signal place_1032_succs : BooleanArray(0 downto 0);
  signal place_1032_token : boolean;
  signal place_1036_preds : BooleanArray(0 downto 0);
  signal place_1036_succs : BooleanArray(0 downto 0);
  signal place_1036_token : boolean;
  signal place_1039_preds : BooleanArray(0 downto 0);
  signal place_1039_succs : BooleanArray(0 downto 0);
  signal place_1039_token : boolean;
  signal place_1047_preds : BooleanArray(0 downto 0);
  signal place_1047_succs : BooleanArray(0 downto 0);
  signal place_1047_token : boolean;
  signal place_1048_preds : BooleanArray(0 downto 0);
  signal place_1048_succs : BooleanArray(0 downto 0);
  signal place_1048_token : boolean;
  signal place_1049_preds : BooleanArray(0 downto 0);
  signal place_1049_succs : BooleanArray(0 downto 0);
  signal place_1049_token : boolean;
  signal place_1050_preds : BooleanArray(0 downto 0);
  signal place_1050_succs : BooleanArray(0 downto 0);
  signal place_1050_token : boolean;
  signal place_1053_preds : BooleanArray(0 downto 0);
  signal place_1053_succs : BooleanArray(0 downto 0);
  signal place_1053_token : boolean;
  signal place_1060_preds : BooleanArray(0 downto 0);
  signal place_1060_succs : BooleanArray(0 downto 0);
  signal place_1060_token : boolean;
  signal place_1061_preds : BooleanArray(0 downto 0);
  signal place_1061_succs : BooleanArray(0 downto 0);
  signal place_1061_token : boolean;
  signal place_1062_preds : BooleanArray(0 downto 0);
  signal place_1062_succs : BooleanArray(0 downto 0);
  signal place_1062_token : boolean;
  signal place_1067_preds : BooleanArray(0 downto 0);
  signal place_1067_succs : BooleanArray(0 downto 0);
  signal place_1067_token : boolean;
  signal place_1068_preds : BooleanArray(0 downto 0);
  signal place_1068_succs : BooleanArray(0 downto 0);
  signal place_1068_token : boolean;
  signal place_1069_preds : BooleanArray(0 downto 0);
  signal place_1069_succs : BooleanArray(0 downto 0);
  signal place_1069_token : boolean;
  signal place_1075_preds : BooleanArray(0 downto 0);
  signal place_1075_succs : BooleanArray(0 downto 0);
  signal place_1075_token : boolean;
  signal place_1076_preds : BooleanArray(0 downto 0);
  signal place_1076_succs : BooleanArray(0 downto 0);
  signal place_1076_token : boolean;
  signal place_1077_preds : BooleanArray(0 downto 0);
  signal place_1077_succs : BooleanArray(0 downto 0);
  signal place_1077_token : boolean;
  signal place_1079_preds : BooleanArray(0 downto 0);
  signal place_1079_succs : BooleanArray(0 downto 0);
  signal place_1079_token : boolean;
  signal place_1082_preds : BooleanArray(0 downto 0);
  signal place_1082_succs : BooleanArray(0 downto 0);
  signal place_1082_token : boolean;
  signal place_1083_preds : BooleanArray(0 downto 0);
  signal place_1083_succs : BooleanArray(0 downto 0);
  signal place_1083_token : boolean;
  signal place_1084_preds : BooleanArray(0 downto 0);
  signal place_1084_succs : BooleanArray(0 downto 0);
  signal place_1084_token : boolean;
  signal place_1085_preds : BooleanArray(0 downto 0);
  signal place_1085_succs : BooleanArray(0 downto 0);
  signal place_1085_token : boolean;
  signal place_1086_preds : BooleanArray(0 downto 0);
  signal place_1086_succs : BooleanArray(0 downto 0);
  signal place_1086_token : boolean;
  signal place_1087_preds : BooleanArray(0 downto 0);
  signal place_1087_succs : BooleanArray(0 downto 0);
  signal place_1087_token : boolean;
  signal place_1088_preds : BooleanArray(0 downto 0);
  signal place_1088_succs : BooleanArray(0 downto 0);
  signal place_1088_token : boolean;
  signal place_1089_preds : BooleanArray(0 downto 0);
  signal place_1089_succs : BooleanArray(0 downto 0);
  signal place_1089_token : boolean;
  signal place_1090_preds : BooleanArray(0 downto 0);
  signal place_1090_succs : BooleanArray(0 downto 0);
  signal place_1090_token : boolean;
  signal place_1091_preds : BooleanArray(0 downto 0);
  signal place_1091_succs : BooleanArray(0 downto 0);
  signal place_1091_token : boolean;
  signal place_1092_preds : BooleanArray(0 downto 0);
  signal place_1092_succs : BooleanArray(0 downto 0);
  signal place_1092_token : boolean;
  signal place_1093_preds : BooleanArray(0 downto 0);
  signal place_1093_succs : BooleanArray(0 downto 0);
  signal place_1093_token : boolean;
  signal place_1094_preds : BooleanArray(0 downto 0);
  signal place_1094_succs : BooleanArray(0 downto 0);
  signal place_1094_token : boolean;
  signal place_1095_preds : BooleanArray(0 downto 0);
  signal place_1095_succs : BooleanArray(0 downto 0);
  signal place_1095_token : boolean;
  signal place_1096_preds : BooleanArray(0 downto 0);
  signal place_1096_succs : BooleanArray(0 downto 0);
  signal place_1096_token : boolean;
  signal place_1097_preds : BooleanArray(0 downto 0);
  signal place_1097_succs : BooleanArray(0 downto 0);
  signal place_1097_token : boolean;
  signal place_1098_preds : BooleanArray(0 downto 0);
  signal place_1098_succs : BooleanArray(0 downto 0);
  signal place_1098_token : boolean;
  signal place_1099_preds : BooleanArray(0 downto 0);
  signal place_1099_succs : BooleanArray(0 downto 0);
  signal place_1099_token : boolean;
  signal place_1100_preds : BooleanArray(0 downto 0);
  signal place_1100_succs : BooleanArray(0 downto 0);
  signal place_1100_token : boolean;
  signal place_1101_preds : BooleanArray(0 downto 0);
  signal place_1101_succs : BooleanArray(0 downto 0);
  signal place_1101_token : boolean;
  signal place_1102_preds : BooleanArray(0 downto 0);
  signal place_1102_succs : BooleanArray(0 downto 0);
  signal place_1102_token : boolean;
  signal place_1103_preds : BooleanArray(0 downto 0);
  signal place_1103_succs : BooleanArray(0 downto 0);
  signal place_1103_token : boolean;
  signal place_1104_preds : BooleanArray(0 downto 0);
  signal place_1104_succs : BooleanArray(0 downto 0);
  signal place_1104_token : boolean;
  signal place_1105_preds : BooleanArray(0 downto 0);
  signal place_1105_succs : BooleanArray(0 downto 0);
  signal place_1105_token : boolean;
  signal place_1106_preds : BooleanArray(0 downto 0);
  signal place_1106_succs : BooleanArray(0 downto 0);
  signal place_1106_token : boolean;
  signal place_1107_preds : BooleanArray(0 downto 0);
  signal place_1107_succs : BooleanArray(0 downto 0);
  signal place_1107_token : boolean;
  signal place_1108_preds : BooleanArray(0 downto 0);
  signal place_1108_succs : BooleanArray(0 downto 0);
  signal place_1108_token : boolean;
  signal place_1109_preds : BooleanArray(0 downto 0);
  signal place_1109_succs : BooleanArray(0 downto 0);
  signal place_1109_token : boolean;
  signal place_1110_preds : BooleanArray(0 downto 0);
  signal place_1110_succs : BooleanArray(0 downto 0);
  signal place_1110_token : boolean;
  signal place_1111_preds : BooleanArray(0 downto 0);
  signal place_1111_succs : BooleanArray(0 downto 0);
  signal place_1111_token : boolean;
  signal place_1112_preds : BooleanArray(0 downto 0);
  signal place_1112_succs : BooleanArray(0 downto 0);
  signal place_1112_token : boolean;
  signal place_1113_preds : BooleanArray(0 downto 0);
  signal place_1113_succs : BooleanArray(0 downto 0);
  signal place_1113_token : boolean;
  signal place_1114_preds : BooleanArray(0 downto 0);
  signal place_1114_succs : BooleanArray(0 downto 0);
  signal place_1114_token : boolean;
  signal place_1115_preds : BooleanArray(0 downto 0);
  signal place_1115_succs : BooleanArray(0 downto 0);
  signal place_1115_token : boolean;
  signal place_1116_preds : BooleanArray(0 downto 0);
  signal place_1116_succs : BooleanArray(0 downto 0);
  signal place_1116_token : boolean;
  signal place_1117_preds : BooleanArray(0 downto 0);
  signal place_1117_succs : BooleanArray(0 downto 0);
  signal place_1117_token : boolean;
  signal place_1118_preds : BooleanArray(0 downto 0);
  signal place_1118_succs : BooleanArray(0 downto 0);
  signal place_1118_token : boolean;
  signal place_1119_preds : BooleanArray(0 downto 0);
  signal place_1119_succs : BooleanArray(0 downto 0);
  signal place_1119_token : boolean;
  signal place_1120_preds : BooleanArray(0 downto 0);
  signal place_1120_succs : BooleanArray(0 downto 0);
  signal place_1120_token : boolean;
  signal place_1121_preds : BooleanArray(0 downto 0);
  signal place_1121_succs : BooleanArray(0 downto 0);
  signal place_1121_token : boolean;
  signal place_1122_preds : BooleanArray(0 downto 0);
  signal place_1122_succs : BooleanArray(0 downto 0);
  signal place_1122_token : boolean;
  signal place_1123_preds : BooleanArray(0 downto 0);
  signal place_1123_succs : BooleanArray(0 downto 0);
  signal place_1123_token : boolean;
  signal place_1124_preds : BooleanArray(0 downto 0);
  signal place_1124_succs : BooleanArray(0 downto 0);
  signal place_1124_token : boolean;
  signal place_1125_preds : BooleanArray(0 downto 0);
  signal place_1125_succs : BooleanArray(0 downto 0);
  signal place_1125_token : boolean;
  signal place_1126_preds : BooleanArray(0 downto 0);
  signal place_1126_succs : BooleanArray(0 downto 0);
  signal place_1126_token : boolean;
  signal place_1127_preds : BooleanArray(0 downto 0);
  signal place_1127_succs : BooleanArray(0 downto 0);
  signal place_1127_token : boolean;
  signal place_1128_preds : BooleanArray(0 downto 0);
  signal place_1128_succs : BooleanArray(0 downto 0);
  signal place_1128_token : boolean;
  signal place_1129_preds : BooleanArray(0 downto 0);
  signal place_1129_succs : BooleanArray(0 downto 0);
  signal place_1129_token : boolean;
  signal place_1130_preds : BooleanArray(0 downto 0);
  signal place_1130_succs : BooleanArray(0 downto 0);
  signal place_1130_token : boolean;
  signal place_1131_preds : BooleanArray(0 downto 0);
  signal place_1131_succs : BooleanArray(0 downto 0);
  signal place_1131_token : boolean;
  signal place_1132_preds : BooleanArray(0 downto 0);
  signal place_1132_succs : BooleanArray(0 downto 0);
  signal place_1132_token : boolean;
  signal place_1133_preds : BooleanArray(0 downto 0);
  signal place_1133_succs : BooleanArray(0 downto 0);
  signal place_1133_token : boolean;
  signal place_1134_preds : BooleanArray(0 downto 0);
  signal place_1134_succs : BooleanArray(0 downto 0);
  signal place_1134_token : boolean;
  signal place_1135_preds : BooleanArray(0 downto 0);
  signal place_1135_succs : BooleanArray(0 downto 0);
  signal place_1135_token : boolean;
  signal place_1136_preds : BooleanArray(0 downto 0);
  signal place_1136_succs : BooleanArray(0 downto 0);
  signal place_1136_token : boolean;
  signal place_1137_preds : BooleanArray(0 downto 0);
  signal place_1137_succs : BooleanArray(0 downto 0);
  signal place_1137_token : boolean;
  signal place_1138_preds : BooleanArray(0 downto 0);
  signal place_1138_succs : BooleanArray(0 downto 0);
  signal place_1138_token : boolean;
  signal place_1139_preds : BooleanArray(0 downto 0);
  signal place_1139_succs : BooleanArray(0 downto 0);
  signal place_1139_token : boolean;
  signal place_1140_preds : BooleanArray(0 downto 0);
  signal place_1140_succs : BooleanArray(0 downto 0);
  signal place_1140_token : boolean;
  signal place_1141_preds : BooleanArray(0 downto 0);
  signal place_1141_succs : BooleanArray(0 downto 0);
  signal place_1141_token : boolean;
  signal place_1142_preds : BooleanArray(0 downto 0);
  signal place_1142_succs : BooleanArray(0 downto 0);
  signal place_1142_token : boolean;
  signal place_1143_preds : BooleanArray(0 downto 0);
  signal place_1143_succs : BooleanArray(0 downto 0);
  signal place_1143_token : boolean;
  signal place_1144_preds : BooleanArray(0 downto 0);
  signal place_1144_succs : BooleanArray(0 downto 0);
  signal place_1144_token : boolean;
  signal place_1145_preds : BooleanArray(0 downto 0);
  signal place_1145_succs : BooleanArray(0 downto 0);
  signal place_1145_token : boolean;
  signal place_1146_preds : BooleanArray(0 downto 0);
  signal place_1146_succs : BooleanArray(0 downto 0);
  signal place_1146_token : boolean;
  signal place_1147_preds : BooleanArray(0 downto 0);
  signal place_1147_succs : BooleanArray(0 downto 0);
  signal place_1147_token : boolean;
  signal place_1148_preds : BooleanArray(0 downto 0);
  signal place_1148_succs : BooleanArray(0 downto 0);
  signal place_1148_token : boolean;
  signal place_1149_preds : BooleanArray(0 downto 0);
  signal place_1149_succs : BooleanArray(0 downto 0);
  signal place_1149_token : boolean;
  signal place_1150_preds : BooleanArray(0 downto 0);
  signal place_1150_succs : BooleanArray(0 downto 0);
  signal place_1150_token : boolean;
  signal place_1151_preds : BooleanArray(0 downto 0);
  signal place_1151_succs : BooleanArray(0 downto 0);
  signal place_1151_token : boolean;
  signal place_1152_preds : BooleanArray(0 downto 0);
  signal place_1152_succs : BooleanArray(0 downto 0);
  signal place_1152_token : boolean;
  signal place_1153_preds : BooleanArray(0 downto 0);
  signal place_1153_succs : BooleanArray(0 downto 0);
  signal place_1153_token : boolean;
  signal place_1154_preds : BooleanArray(0 downto 0);
  signal place_1154_succs : BooleanArray(0 downto 0);
  signal place_1154_token : boolean;
  signal place_1155_preds : BooleanArray(0 downto 0);
  signal place_1155_succs : BooleanArray(0 downto 0);
  signal place_1155_token : boolean;
  signal place_1156_preds : BooleanArray(0 downto 0);
  signal place_1156_succs : BooleanArray(0 downto 0);
  signal place_1156_token : boolean;
  signal place_1157_preds : BooleanArray(0 downto 0);
  signal place_1157_succs : BooleanArray(0 downto 0);
  signal place_1157_token : boolean;
  signal place_1158_preds : BooleanArray(0 downto 0);
  signal place_1158_succs : BooleanArray(0 downto 0);
  signal place_1158_token : boolean;
  signal place_1159_preds : BooleanArray(0 downto 0);
  signal place_1159_succs : BooleanArray(0 downto 0);
  signal place_1159_token : boolean;
  signal place_1160_preds : BooleanArray(0 downto 0);
  signal place_1160_succs : BooleanArray(0 downto 0);
  signal place_1160_token : boolean;
  signal place_1161_preds : BooleanArray(0 downto 0);
  signal place_1161_succs : BooleanArray(0 downto 0);
  signal place_1161_token : boolean;
  signal place_1162_preds : BooleanArray(0 downto 0);
  signal place_1162_succs : BooleanArray(0 downto 0);
  signal place_1162_token : boolean;
  signal place_1163_preds : BooleanArray(0 downto 0);
  signal place_1163_succs : BooleanArray(0 downto 0);
  signal place_1163_token : boolean;
  signal place_1164_preds : BooleanArray(0 downto 0);
  signal place_1164_succs : BooleanArray(0 downto 0);
  signal place_1164_token : boolean;
  signal place_1165_preds : BooleanArray(0 downto 0);
  signal place_1165_succs : BooleanArray(0 downto 0);
  signal place_1165_token : boolean;
  signal place_1166_preds : BooleanArray(0 downto 0);
  signal place_1166_succs : BooleanArray(0 downto 0);
  signal place_1166_token : boolean;
  signal place_1167_preds : BooleanArray(0 downto 0);
  signal place_1167_succs : BooleanArray(0 downto 0);
  signal place_1167_token : boolean;
  signal place_1168_preds : BooleanArray(0 downto 0);
  signal place_1168_succs : BooleanArray(0 downto 0);
  signal place_1168_token : boolean;
  signal place_1169_preds : BooleanArray(0 downto 0);
  signal place_1169_succs : BooleanArray(0 downto 0);
  signal place_1169_token : boolean;
  signal place_1170_preds : BooleanArray(0 downto 0);
  signal place_1170_succs : BooleanArray(0 downto 0);
  signal place_1170_token : boolean;
  signal place_1171_preds : BooleanArray(0 downto 0);
  signal place_1171_succs : BooleanArray(0 downto 0);
  signal place_1171_token : boolean;
  signal place_1172_preds : BooleanArray(0 downto 0);
  signal place_1172_succs : BooleanArray(0 downto 0);
  signal place_1172_token : boolean;
  signal place_1173_preds : BooleanArray(0 downto 0);
  signal place_1173_succs : BooleanArray(0 downto 0);
  signal place_1173_token : boolean;
  signal place_1174_preds : BooleanArray(0 downto 0);
  signal place_1174_succs : BooleanArray(0 downto 0);
  signal place_1174_token : boolean;
  signal place_1175_preds : BooleanArray(0 downto 0);
  signal place_1175_succs : BooleanArray(0 downto 0);
  signal place_1175_token : boolean;
  signal place_1176_preds : BooleanArray(0 downto 0);
  signal place_1176_succs : BooleanArray(0 downto 0);
  signal place_1176_token : boolean;
  signal place_1177_preds : BooleanArray(0 downto 0);
  signal place_1177_succs : BooleanArray(0 downto 0);
  signal place_1177_token : boolean;
  signal place_1178_preds : BooleanArray(0 downto 0);
  signal place_1178_succs : BooleanArray(0 downto 0);
  signal place_1178_token : boolean;
  signal place_1179_preds : BooleanArray(0 downto 0);
  signal place_1179_succs : BooleanArray(0 downto 0);
  signal place_1179_token : boolean;
  signal place_1180_preds : BooleanArray(0 downto 0);
  signal place_1180_succs : BooleanArray(0 downto 0);
  signal place_1180_token : boolean;
  signal place_1181_preds : BooleanArray(0 downto 0);
  signal place_1181_succs : BooleanArray(0 downto 0);
  signal place_1181_token : boolean;
  signal place_1182_preds : BooleanArray(0 downto 0);
  signal place_1182_succs : BooleanArray(0 downto 0);
  signal place_1182_token : boolean;
  signal place_1183_preds : BooleanArray(0 downto 0);
  signal place_1183_succs : BooleanArray(0 downto 0);
  signal place_1183_token : boolean;
  signal place_1184_preds : BooleanArray(0 downto 0);
  signal place_1184_succs : BooleanArray(0 downto 0);
  signal place_1184_token : boolean;
  signal place_1185_preds : BooleanArray(0 downto 0);
  signal place_1185_succs : BooleanArray(0 downto 0);
  signal place_1185_token : boolean;
  signal place_1186_preds : BooleanArray(0 downto 0);
  signal place_1186_succs : BooleanArray(0 downto 0);
  signal place_1186_token : boolean;
  signal place_1187_preds : BooleanArray(0 downto 0);
  signal place_1187_succs : BooleanArray(0 downto 0);
  signal place_1187_token : boolean;
  signal place_1188_preds : BooleanArray(0 downto 0);
  signal place_1188_succs : BooleanArray(0 downto 0);
  signal place_1188_token : boolean;
  signal place_1189_preds : BooleanArray(0 downto 0);
  signal place_1189_succs : BooleanArray(0 downto 0);
  signal place_1189_token : boolean;
  signal place_1190_preds : BooleanArray(0 downto 0);
  signal place_1190_succs : BooleanArray(0 downto 0);
  signal place_1190_token : boolean;
  signal place_1191_preds : BooleanArray(0 downto 0);
  signal place_1191_succs : BooleanArray(0 downto 0);
  signal place_1191_token : boolean;
  signal place_1192_preds : BooleanArray(0 downto 0);
  signal place_1192_succs : BooleanArray(0 downto 0);
  signal place_1192_token : boolean;
  signal place_1193_preds : BooleanArray(0 downto 0);
  signal place_1193_succs : BooleanArray(0 downto 0);
  signal place_1193_token : boolean;
  signal place_1194_preds : BooleanArray(0 downto 0);
  signal place_1194_succs : BooleanArray(0 downto 0);
  signal place_1194_token : boolean;
  signal place_1195_preds : BooleanArray(0 downto 0);
  signal place_1195_succs : BooleanArray(0 downto 0);
  signal place_1195_token : boolean;
  signal place_1196_preds : BooleanArray(0 downto 0);
  signal place_1196_succs : BooleanArray(0 downto 0);
  signal place_1196_token : boolean;
  signal place_1197_preds : BooleanArray(0 downto 0);
  signal place_1197_succs : BooleanArray(0 downto 0);
  signal place_1197_token : boolean;
  signal place_1198_preds : BooleanArray(0 downto 0);
  signal place_1198_succs : BooleanArray(0 downto 0);
  signal place_1198_token : boolean;
  signal place_1199_preds : BooleanArray(0 downto 0);
  signal place_1199_succs : BooleanArray(0 downto 0);
  signal place_1199_token : boolean;
  signal place_1200_preds : BooleanArray(0 downto 0);
  signal place_1200_succs : BooleanArray(0 downto 0);
  signal place_1200_token : boolean;
  signal place_1201_preds : BooleanArray(0 downto 0);
  signal place_1201_succs : BooleanArray(0 downto 0);
  signal place_1201_token : boolean;
  signal place_1202_preds : BooleanArray(0 downto 0);
  signal place_1202_succs : BooleanArray(0 downto 0);
  signal place_1202_token : boolean;
  signal place_1203_preds : BooleanArray(0 downto 0);
  signal place_1203_succs : BooleanArray(0 downto 0);
  signal place_1203_token : boolean;
  signal place_1204_preds : BooleanArray(0 downto 0);
  signal place_1204_succs : BooleanArray(0 downto 0);
  signal place_1204_token : boolean;
  signal place_1205_preds : BooleanArray(0 downto 0);
  signal place_1205_succs : BooleanArray(0 downto 0);
  signal place_1205_token : boolean;
  signal place_1206_preds : BooleanArray(0 downto 0);
  signal place_1206_succs : BooleanArray(0 downto 0);
  signal place_1206_token : boolean;
  signal place_1207_preds : BooleanArray(0 downto 0);
  signal place_1207_succs : BooleanArray(0 downto 0);
  signal place_1207_token : boolean;
  signal place_1208_preds : BooleanArray(0 downto 0);
  signal place_1208_succs : BooleanArray(0 downto 0);
  signal place_1208_token : boolean;
  signal place_1209_preds : BooleanArray(0 downto 0);
  signal place_1209_succs : BooleanArray(0 downto 0);
  signal place_1209_token : boolean;
  signal place_1210_preds : BooleanArray(0 downto 0);
  signal place_1210_succs : BooleanArray(0 downto 0);
  signal place_1210_token : boolean;
  signal place_1211_preds : BooleanArray(0 downto 0);
  signal place_1211_succs : BooleanArray(0 downto 0);
  signal place_1211_token : boolean;
  signal place_1212_preds : BooleanArray(0 downto 0);
  signal place_1212_succs : BooleanArray(0 downto 0);
  signal place_1212_token : boolean;
  signal place_1213_preds : BooleanArray(0 downto 0);
  signal place_1213_succs : BooleanArray(0 downto 0);
  signal place_1213_token : boolean;
  signal place_1214_preds : BooleanArray(0 downto 0);
  signal place_1214_succs : BooleanArray(0 downto 0);
  signal place_1214_token : boolean;
  signal place_1215_preds : BooleanArray(0 downto 0);
  signal place_1215_succs : BooleanArray(0 downto 0);
  signal place_1215_token : boolean;
  signal place_1216_preds : BooleanArray(0 downto 0);
  signal place_1216_succs : BooleanArray(0 downto 0);
  signal place_1216_token : boolean;
  signal place_1217_preds : BooleanArray(0 downto 0);
  signal place_1217_succs : BooleanArray(0 downto 0);
  signal place_1217_token : boolean;
  signal place_1218_preds : BooleanArray(0 downto 0);
  signal place_1218_succs : BooleanArray(0 downto 0);
  signal place_1218_token : boolean;
  signal place_1219_preds : BooleanArray(0 downto 0);
  signal place_1219_succs : BooleanArray(0 downto 0);
  signal place_1219_token : boolean;
  signal place_1220_preds : BooleanArray(0 downto 0);
  signal place_1220_succs : BooleanArray(0 downto 0);
  signal place_1220_token : boolean;
  signal place_1221_preds : BooleanArray(0 downto 0);
  signal place_1221_succs : BooleanArray(0 downto 0);
  signal place_1221_token : boolean;
  signal place_1222_preds : BooleanArray(0 downto 0);
  signal place_1222_succs : BooleanArray(0 downto 0);
  signal place_1222_token : boolean;
  signal place_1223_preds : BooleanArray(0 downto 0);
  signal place_1223_succs : BooleanArray(0 downto 0);
  signal place_1223_token : boolean;
  signal place_1224_preds : BooleanArray(0 downto 0);
  signal place_1224_succs : BooleanArray(0 downto 0);
  signal place_1224_token : boolean;
  signal place_1225_preds : BooleanArray(0 downto 0);
  signal place_1225_succs : BooleanArray(0 downto 0);
  signal place_1225_token : boolean;
  signal place_1226_preds : BooleanArray(0 downto 0);
  signal place_1226_succs : BooleanArray(0 downto 0);
  signal place_1226_token : boolean;
  signal place_1227_preds : BooleanArray(0 downto 0);
  signal place_1227_succs : BooleanArray(0 downto 0);
  signal place_1227_token : boolean;
  signal place_1228_preds : BooleanArray(0 downto 0);
  signal place_1228_succs : BooleanArray(0 downto 0);
  signal place_1228_token : boolean;
  signal place_1229_preds : BooleanArray(0 downto 0);
  signal place_1229_succs : BooleanArray(0 downto 0);
  signal place_1229_token : boolean;
  signal place_1230_preds : BooleanArray(0 downto 0);
  signal place_1230_succs : BooleanArray(0 downto 0);
  signal place_1230_token : boolean;
  signal place_1231_preds : BooleanArray(0 downto 0);
  signal place_1231_succs : BooleanArray(0 downto 0);
  signal place_1231_token : boolean;
  signal place_1232_preds : BooleanArray(0 downto 0);
  signal place_1232_succs : BooleanArray(0 downto 0);
  signal place_1232_token : boolean;
  signal place_1233_preds : BooleanArray(0 downto 0);
  signal place_1233_succs : BooleanArray(0 downto 0);
  signal place_1233_token : boolean;
  signal place_1234_preds : BooleanArray(0 downto 0);
  signal place_1234_succs : BooleanArray(0 downto 0);
  signal place_1234_token : boolean;
  signal place_1235_preds : BooleanArray(0 downto 0);
  signal place_1235_succs : BooleanArray(0 downto 0);
  signal place_1235_token : boolean;
  signal place_1236_preds : BooleanArray(0 downto 0);
  signal place_1236_succs : BooleanArray(0 downto 0);
  signal place_1236_token : boolean;
  signal place_1237_preds : BooleanArray(0 downto 0);
  signal place_1237_succs : BooleanArray(0 downto 0);
  signal place_1237_token : boolean;
  signal place_1238_preds : BooleanArray(0 downto 0);
  signal place_1238_succs : BooleanArray(0 downto 0);
  signal place_1238_token : boolean;
  signal place_1239_preds : BooleanArray(0 downto 0);
  signal place_1239_succs : BooleanArray(0 downto 0);
  signal place_1239_token : boolean;
  signal place_1240_preds : BooleanArray(0 downto 0);
  signal place_1240_succs : BooleanArray(0 downto 0);
  signal place_1240_token : boolean;
  signal place_1241_preds : BooleanArray(0 downto 0);
  signal place_1241_succs : BooleanArray(0 downto 0);
  signal place_1241_token : boolean;
  signal place_1242_preds : BooleanArray(0 downto 0);
  signal place_1242_succs : BooleanArray(0 downto 0);
  signal place_1242_token : boolean;
  signal place_1243_preds : BooleanArray(0 downto 0);
  signal place_1243_succs : BooleanArray(0 downto 0);
  signal place_1243_token : boolean;
  signal place_1244_preds : BooleanArray(0 downto 0);
  signal place_1244_succs : BooleanArray(0 downto 0);
  signal place_1244_token : boolean;
  signal place_1245_preds : BooleanArray(0 downto 0);
  signal place_1245_succs : BooleanArray(0 downto 0);
  signal place_1245_token : boolean;
  signal place_1246_preds : BooleanArray(0 downto 0);
  signal place_1246_succs : BooleanArray(0 downto 0);
  signal place_1246_token : boolean;
  signal place_1247_preds : BooleanArray(0 downto 0);
  signal place_1247_succs : BooleanArray(0 downto 0);
  signal place_1247_token : boolean;
  signal place_1248_preds : BooleanArray(0 downto 0);
  signal place_1248_succs : BooleanArray(0 downto 0);
  signal place_1248_token : boolean;
  signal place_1249_preds : BooleanArray(0 downto 0);
  signal place_1249_succs : BooleanArray(0 downto 0);
  signal place_1249_token : boolean;
  signal place_1250_preds : BooleanArray(0 downto 0);
  signal place_1250_succs : BooleanArray(0 downto 0);
  signal place_1250_token : boolean;
  signal place_1251_preds : BooleanArray(0 downto 0);
  signal place_1251_succs : BooleanArray(0 downto 0);
  signal place_1251_token : boolean;
  signal place_1252_preds : BooleanArray(0 downto 0);
  signal place_1252_succs : BooleanArray(0 downto 0);
  signal place_1252_token : boolean;
  signal place_1253_preds : BooleanArray(0 downto 0);
  signal place_1253_succs : BooleanArray(0 downto 0);
  signal place_1253_token : boolean;
  signal place_1254_preds : BooleanArray(0 downto 0);
  signal place_1254_succs : BooleanArray(0 downto 0);
  signal place_1254_token : boolean;
  signal place_1255_preds : BooleanArray(0 downto 0);
  signal place_1255_succs : BooleanArray(0 downto 0);
  signal place_1255_token : boolean;
  signal place_1256_preds : BooleanArray(0 downto 0);
  signal place_1256_succs : BooleanArray(0 downto 0);
  signal place_1256_token : boolean;
  signal place_1257_preds : BooleanArray(0 downto 0);
  signal place_1257_succs : BooleanArray(0 downto 0);
  signal place_1257_token : boolean;
  signal place_1258_preds : BooleanArray(0 downto 0);
  signal place_1258_succs : BooleanArray(0 downto 0);
  signal place_1258_token : boolean;
  signal place_1259_preds : BooleanArray(0 downto 0);
  signal place_1259_succs : BooleanArray(0 downto 0);
  signal place_1259_token : boolean;
  signal place_1260_preds : BooleanArray(0 downto 0);
  signal place_1260_succs : BooleanArray(0 downto 0);
  signal place_1260_token : boolean;
  signal place_1261_preds : BooleanArray(0 downto 0);
  signal place_1261_succs : BooleanArray(0 downto 0);
  signal place_1261_token : boolean;
  signal place_1262_preds : BooleanArray(0 downto 0);
  signal place_1262_succs : BooleanArray(0 downto 0);
  signal place_1262_token : boolean;
  signal place_1263_preds : BooleanArray(0 downto 0);
  signal place_1263_succs : BooleanArray(0 downto 0);
  signal place_1263_token : boolean;
  signal place_1264_preds : BooleanArray(0 downto 0);
  signal place_1264_succs : BooleanArray(0 downto 0);
  signal place_1264_token : boolean;
  signal place_1265_preds : BooleanArray(0 downto 0);
  signal place_1265_succs : BooleanArray(0 downto 0);
  signal place_1265_token : boolean;
  signal place_1266_preds : BooleanArray(0 downto 0);
  signal place_1266_succs : BooleanArray(0 downto 0);
  signal place_1266_token : boolean;
  signal place_1267_preds : BooleanArray(0 downto 0);
  signal place_1267_succs : BooleanArray(0 downto 0);
  signal place_1267_token : boolean;
  signal place_1268_preds : BooleanArray(0 downto 0);
  signal place_1268_succs : BooleanArray(0 downto 0);
  signal place_1268_token : boolean;
  signal place_1269_preds : BooleanArray(0 downto 0);
  signal place_1269_succs : BooleanArray(0 downto 0);
  signal place_1269_token : boolean;
  signal place_1270_preds : BooleanArray(0 downto 0);
  signal place_1270_succs : BooleanArray(0 downto 0);
  signal place_1270_token : boolean;
  signal place_1271_preds : BooleanArray(0 downto 0);
  signal place_1271_succs : BooleanArray(0 downto 0);
  signal place_1271_token : boolean;
  signal place_1272_preds : BooleanArray(0 downto 0);
  signal place_1272_succs : BooleanArray(0 downto 0);
  signal place_1272_token : boolean;
  signal place_1273_preds : BooleanArray(0 downto 0);
  signal place_1273_succs : BooleanArray(0 downto 0);
  signal place_1273_token : boolean;
  signal place_1274_preds : BooleanArray(0 downto 0);
  signal place_1274_succs : BooleanArray(0 downto 0);
  signal place_1274_token : boolean;
  signal place_1275_preds : BooleanArray(0 downto 0);
  signal place_1275_succs : BooleanArray(0 downto 0);
  signal place_1275_token : boolean;
  signal place_1276_preds : BooleanArray(0 downto 0);
  signal place_1276_succs : BooleanArray(0 downto 0);
  signal place_1276_token : boolean;
  signal place_1277_preds : BooleanArray(0 downto 0);
  signal place_1277_succs : BooleanArray(0 downto 0);
  signal place_1277_token : boolean;
  signal place_1278_preds : BooleanArray(0 downto 0);
  signal place_1278_succs : BooleanArray(0 downto 0);
  signal place_1278_token : boolean;
  signal place_1279_preds : BooleanArray(0 downto 0);
  signal place_1279_succs : BooleanArray(0 downto 0);
  signal place_1279_token : boolean;
  signal place_1280_preds : BooleanArray(0 downto 0);
  signal place_1280_succs : BooleanArray(0 downto 0);
  signal place_1280_token : boolean;
  signal place_1281_preds : BooleanArray(0 downto 0);
  signal place_1281_succs : BooleanArray(0 downto 0);
  signal place_1281_token : boolean;
  signal place_1282_preds : BooleanArray(0 downto 0);
  signal place_1282_succs : BooleanArray(0 downto 0);
  signal place_1282_token : boolean;
  signal place_1283_preds : BooleanArray(0 downto 0);
  signal place_1283_succs : BooleanArray(0 downto 0);
  signal place_1283_token : boolean;
  signal place_1284_preds : BooleanArray(0 downto 0);
  signal place_1284_succs : BooleanArray(0 downto 0);
  signal place_1284_token : boolean;
  signal place_1285_preds : BooleanArray(0 downto 0);
  signal place_1285_succs : BooleanArray(0 downto 0);
  signal place_1285_token : boolean;
  signal place_1286_preds : BooleanArray(0 downto 0);
  signal place_1286_succs : BooleanArray(0 downto 0);
  signal place_1286_token : boolean;
  signal place_1287_preds : BooleanArray(0 downto 0);
  signal place_1287_succs : BooleanArray(0 downto 0);
  signal place_1287_token : boolean;
  signal place_1288_preds : BooleanArray(0 downto 0);
  signal place_1288_succs : BooleanArray(0 downto 0);
  signal place_1288_token : boolean;
  signal place_1289_preds : BooleanArray(0 downto 0);
  signal place_1289_succs : BooleanArray(0 downto 0);
  signal place_1289_token : boolean;
  signal place_1290_preds : BooleanArray(0 downto 0);
  signal place_1290_succs : BooleanArray(0 downto 0);
  signal place_1290_token : boolean;
  signal place_1291_preds : BooleanArray(0 downto 0);
  signal place_1291_succs : BooleanArray(0 downto 0);
  signal place_1291_token : boolean;
  signal place_1292_preds : BooleanArray(0 downto 0);
  signal place_1292_succs : BooleanArray(0 downto 0);
  signal place_1292_token : boolean;
  signal place_1293_preds : BooleanArray(0 downto 0);
  signal place_1293_succs : BooleanArray(0 downto 0);
  signal place_1293_token : boolean;
  signal place_1294_preds : BooleanArray(0 downto 0);
  signal place_1294_succs : BooleanArray(0 downto 0);
  signal place_1294_token : boolean;
  signal place_1295_preds : BooleanArray(0 downto 0);
  signal place_1295_succs : BooleanArray(0 downto 0);
  signal place_1295_token : boolean;
  signal place_1296_preds : BooleanArray(0 downto 0);
  signal place_1296_succs : BooleanArray(0 downto 0);
  signal place_1296_token : boolean;
  signal place_1297_preds : BooleanArray(0 downto 0);
  signal place_1297_succs : BooleanArray(0 downto 0);
  signal place_1297_token : boolean;
  signal place_1298_preds : BooleanArray(0 downto 0);
  signal place_1298_succs : BooleanArray(0 downto 0);
  signal place_1298_token : boolean;
  signal place_1299_preds : BooleanArray(0 downto 0);
  signal place_1299_succs : BooleanArray(0 downto 0);
  signal place_1299_token : boolean;
  signal place_1300_preds : BooleanArray(0 downto 0);
  signal place_1300_succs : BooleanArray(0 downto 0);
  signal place_1300_token : boolean;
  signal place_1301_preds : BooleanArray(0 downto 0);
  signal place_1301_succs : BooleanArray(0 downto 0);
  signal place_1301_token : boolean;
  signal place_1302_preds : BooleanArray(0 downto 0);
  signal place_1302_succs : BooleanArray(0 downto 0);
  signal place_1302_token : boolean;
  signal place_1303_preds : BooleanArray(0 downto 0);
  signal place_1303_succs : BooleanArray(0 downto 0);
  signal place_1303_token : boolean;
  signal place_1304_preds : BooleanArray(0 downto 0);
  signal place_1304_succs : BooleanArray(0 downto 0);
  signal place_1304_token : boolean;
  signal place_1305_preds : BooleanArray(0 downto 0);
  signal place_1305_succs : BooleanArray(0 downto 0);
  signal place_1305_token : boolean;
  signal place_1306_preds : BooleanArray(0 downto 0);
  signal place_1306_succs : BooleanArray(0 downto 0);
  signal place_1306_token : boolean;
  signal place_1307_preds : BooleanArray(0 downto 0);
  signal place_1307_succs : BooleanArray(0 downto 0);
  signal place_1307_token : boolean;
  signal place_1308_preds : BooleanArray(0 downto 0);
  signal place_1308_succs : BooleanArray(0 downto 0);
  signal place_1308_token : boolean;
  signal place_1309_preds : BooleanArray(0 downto 0);
  signal place_1309_succs : BooleanArray(0 downto 0);
  signal place_1309_token : boolean;
  signal place_1310_preds : BooleanArray(0 downto 0);
  signal place_1310_succs : BooleanArray(0 downto 0);
  signal place_1310_token : boolean;
  signal place_1311_preds : BooleanArray(0 downto 0);
  signal place_1311_succs : BooleanArray(0 downto 0);
  signal place_1311_token : boolean;
  signal place_1312_preds : BooleanArray(0 downto 0);
  signal place_1312_succs : BooleanArray(0 downto 0);
  signal place_1312_token : boolean;
  signal place_1313_preds : BooleanArray(0 downto 0);
  signal place_1313_succs : BooleanArray(0 downto 0);
  signal place_1313_token : boolean;
  signal place_1314_preds : BooleanArray(0 downto 0);
  signal place_1314_succs : BooleanArray(0 downto 0);
  signal place_1314_token : boolean;
  signal place_1315_preds : BooleanArray(0 downto 0);
  signal place_1315_succs : BooleanArray(0 downto 0);
  signal place_1315_token : boolean;
  signal place_1316_preds : BooleanArray(0 downto 0);
  signal place_1316_succs : BooleanArray(0 downto 0);
  signal place_1316_token : boolean;
  signal place_1317_preds : BooleanArray(0 downto 0);
  signal place_1317_succs : BooleanArray(0 downto 0);
  signal place_1317_token : boolean;
  signal place_1318_preds : BooleanArray(0 downto 0);
  signal place_1318_succs : BooleanArray(0 downto 0);
  signal place_1318_token : boolean;
  signal place_1319_preds : BooleanArray(0 downto 0);
  signal place_1319_succs : BooleanArray(0 downto 0);
  signal place_1319_token : boolean;
  signal place_1320_preds : BooleanArray(0 downto 0);
  signal place_1320_succs : BooleanArray(0 downto 0);
  signal place_1320_token : boolean;
  signal place_1321_preds : BooleanArray(0 downto 0);
  signal place_1321_succs : BooleanArray(0 downto 0);
  signal place_1321_token : boolean;
  signal place_1322_preds : BooleanArray(0 downto 0);
  signal place_1322_succs : BooleanArray(0 downto 0);
  signal place_1322_token : boolean;
  signal place_1323_preds : BooleanArray(0 downto 0);
  signal place_1323_succs : BooleanArray(0 downto 0);
  signal place_1323_token : boolean;
  signal place_1324_preds : BooleanArray(0 downto 0);
  signal place_1324_succs : BooleanArray(0 downto 0);
  signal place_1324_token : boolean;
  signal place_1325_preds : BooleanArray(0 downto 0);
  signal place_1325_succs : BooleanArray(0 downto 0);
  signal place_1325_token : boolean;
  signal place_1326_preds : BooleanArray(0 downto 0);
  signal place_1326_succs : BooleanArray(0 downto 0);
  signal place_1326_token : boolean;
  signal place_1327_preds : BooleanArray(0 downto 0);
  signal place_1327_succs : BooleanArray(0 downto 0);
  signal place_1327_token : boolean;
  signal place_1328_preds : BooleanArray(0 downto 0);
  signal place_1328_succs : BooleanArray(0 downto 0);
  signal place_1328_token : boolean;
  signal place_1329_preds : BooleanArray(0 downto 0);
  signal place_1329_succs : BooleanArray(0 downto 0);
  signal place_1329_token : boolean;
  signal place_1330_preds : BooleanArray(0 downto 0);
  signal place_1330_succs : BooleanArray(0 downto 0);
  signal place_1330_token : boolean;
  signal place_1331_preds : BooleanArray(0 downto 0);
  signal place_1331_succs : BooleanArray(0 downto 0);
  signal place_1331_token : boolean;
  signal place_1332_preds : BooleanArray(0 downto 0);
  signal place_1332_succs : BooleanArray(0 downto 0);
  signal place_1332_token : boolean;
  signal place_1333_preds : BooleanArray(0 downto 0);
  signal place_1333_succs : BooleanArray(0 downto 0);
  signal place_1333_token : boolean;
  signal place_1334_preds : BooleanArray(0 downto 0);
  signal place_1334_succs : BooleanArray(0 downto 0);
  signal place_1334_token : boolean;
  signal place_1335_preds : BooleanArray(0 downto 0);
  signal place_1335_succs : BooleanArray(0 downto 0);
  signal place_1335_token : boolean;
  signal place_1336_preds : BooleanArray(0 downto 0);
  signal place_1336_succs : BooleanArray(0 downto 0);
  signal place_1336_token : boolean;
  signal place_1337_preds : BooleanArray(0 downto 0);
  signal place_1337_succs : BooleanArray(0 downto 0);
  signal place_1337_token : boolean;
  signal place_1338_preds : BooleanArray(0 downto 0);
  signal place_1338_succs : BooleanArray(0 downto 0);
  signal place_1338_token : boolean;
  signal place_1339_preds : BooleanArray(0 downto 0);
  signal place_1339_succs : BooleanArray(0 downto 0);
  signal place_1339_token : boolean;
  signal place_1340_preds : BooleanArray(0 downto 0);
  signal place_1340_succs : BooleanArray(0 downto 0);
  signal place_1340_token : boolean;
  signal place_1341_preds : BooleanArray(0 downto 0);
  signal place_1341_succs : BooleanArray(0 downto 0);
  signal place_1341_token : boolean;
  signal place_1342_preds : BooleanArray(0 downto 0);
  signal place_1342_succs : BooleanArray(0 downto 0);
  signal place_1342_token : boolean;
  signal place_1343_preds : BooleanArray(0 downto 0);
  signal place_1343_succs : BooleanArray(0 downto 0);
  signal place_1343_token : boolean;
  signal place_1344_preds : BooleanArray(0 downto 0);
  signal place_1344_succs : BooleanArray(0 downto 0);
  signal place_1344_token : boolean;
  signal place_1345_preds : BooleanArray(0 downto 0);
  signal place_1345_succs : BooleanArray(0 downto 0);
  signal place_1345_token : boolean;
  signal place_1346_preds : BooleanArray(0 downto 0);
  signal place_1346_succs : BooleanArray(0 downto 0);
  signal place_1346_token : boolean;
  signal place_1347_preds : BooleanArray(0 downto 0);
  signal place_1347_succs : BooleanArray(0 downto 0);
  signal place_1347_token : boolean;
  signal place_1348_preds : BooleanArray(0 downto 0);
  signal place_1348_succs : BooleanArray(0 downto 0);
  signal place_1348_token : boolean;
  signal place_1349_preds : BooleanArray(0 downto 0);
  signal place_1349_succs : BooleanArray(0 downto 0);
  signal place_1349_token : boolean;
  signal place_1350_preds : BooleanArray(0 downto 0);
  signal place_1350_succs : BooleanArray(0 downto 0);
  signal place_1350_token : boolean;
  signal place_1351_preds : BooleanArray(0 downto 0);
  signal place_1351_succs : BooleanArray(0 downto 0);
  signal place_1351_token : boolean;
  signal place_1352_preds : BooleanArray(0 downto 0);
  signal place_1352_succs : BooleanArray(0 downto 0);
  signal place_1352_token : boolean;
  signal place_1353_preds : BooleanArray(0 downto 0);
  signal place_1353_succs : BooleanArray(0 downto 0);
  signal place_1353_token : boolean;
  signal place_1354_preds : BooleanArray(0 downto 0);
  signal place_1354_succs : BooleanArray(0 downto 0);
  signal place_1354_token : boolean;
  signal place_1355_preds : BooleanArray(0 downto 0);
  signal place_1355_succs : BooleanArray(0 downto 0);
  signal place_1355_token : boolean;
  signal place_1356_preds : BooleanArray(0 downto 0);
  signal place_1356_succs : BooleanArray(0 downto 0);
  signal place_1356_token : boolean;
  signal place_1357_preds : BooleanArray(0 downto 0);
  signal place_1357_succs : BooleanArray(0 downto 0);
  signal place_1357_token : boolean;
  signal place_1358_preds : BooleanArray(0 downto 0);
  signal place_1358_succs : BooleanArray(0 downto 0);
  signal place_1358_token : boolean;
  signal place_1359_preds : BooleanArray(0 downto 0);
  signal place_1359_succs : BooleanArray(0 downto 0);
  signal place_1359_token : boolean;
  signal place_1360_preds : BooleanArray(0 downto 0);
  signal place_1360_succs : BooleanArray(0 downto 0);
  signal place_1360_token : boolean;
  signal place_1361_preds : BooleanArray(0 downto 0);
  signal place_1361_succs : BooleanArray(0 downto 0);
  signal place_1361_token : boolean;
  signal place_1362_preds : BooleanArray(0 downto 0);
  signal place_1362_succs : BooleanArray(0 downto 0);
  signal place_1362_token : boolean;
  signal place_1363_preds : BooleanArray(0 downto 0);
  signal place_1363_succs : BooleanArray(0 downto 0);
  signal place_1363_token : boolean;
  signal place_1364_preds : BooleanArray(0 downto 0);
  signal place_1364_succs : BooleanArray(0 downto 0);
  signal place_1364_token : boolean;
  signal place_1365_preds : BooleanArray(0 downto 0);
  signal place_1365_succs : BooleanArray(0 downto 0);
  signal place_1365_token : boolean;
  signal place_1366_preds : BooleanArray(0 downto 0);
  signal place_1366_succs : BooleanArray(0 downto 0);
  signal place_1366_token : boolean;
  signal place_1367_preds : BooleanArray(0 downto 0);
  signal place_1367_succs : BooleanArray(0 downto 0);
  signal place_1367_token : boolean;
  signal place_1368_preds : BooleanArray(0 downto 0);
  signal place_1368_succs : BooleanArray(0 downto 0);
  signal place_1368_token : boolean;
  signal place_1369_preds : BooleanArray(0 downto 0);
  signal place_1369_succs : BooleanArray(0 downto 0);
  signal place_1369_token : boolean;
  signal place_1370_preds : BooleanArray(0 downto 0);
  signal place_1370_succs : BooleanArray(0 downto 0);
  signal place_1370_token : boolean;
  signal place_1371_preds : BooleanArray(0 downto 0);
  signal place_1371_succs : BooleanArray(0 downto 0);
  signal place_1371_token : boolean;
  signal place_1372_preds : BooleanArray(0 downto 0);
  signal place_1372_succs : BooleanArray(0 downto 0);
  signal place_1372_token : boolean;
  signal place_1373_preds : BooleanArray(0 downto 0);
  signal place_1373_succs : BooleanArray(0 downto 0);
  signal place_1373_token : boolean;
  signal place_1374_preds : BooleanArray(0 downto 0);
  signal place_1374_succs : BooleanArray(0 downto 0);
  signal place_1374_token : boolean;
  signal place_1375_preds : BooleanArray(0 downto 0);
  signal place_1375_succs : BooleanArray(0 downto 0);
  signal place_1375_token : boolean;
  signal place_1376_preds : BooleanArray(0 downto 0);
  signal place_1376_succs : BooleanArray(0 downto 0);
  signal place_1376_token : boolean;
  signal place_1377_preds : BooleanArray(0 downto 0);
  signal place_1377_succs : BooleanArray(0 downto 0);
  signal place_1377_token : boolean;
  signal place_1378_preds : BooleanArray(0 downto 0);
  signal place_1378_succs : BooleanArray(0 downto 0);
  signal place_1378_token : boolean;
  signal place_1379_preds : BooleanArray(0 downto 0);
  signal place_1379_succs : BooleanArray(0 downto 0);
  signal place_1379_token : boolean;
  signal place_1380_preds : BooleanArray(0 downto 0);
  signal place_1380_succs : BooleanArray(0 downto 0);
  signal place_1380_token : boolean;
  signal place_1381_preds : BooleanArray(0 downto 0);
  signal place_1381_succs : BooleanArray(0 downto 0);
  signal place_1381_token : boolean;
  signal place_1382_preds : BooleanArray(0 downto 0);
  signal place_1382_succs : BooleanArray(0 downto 0);
  signal place_1382_token : boolean;
  signal place_1383_preds : BooleanArray(0 downto 0);
  signal place_1383_succs : BooleanArray(0 downto 0);
  signal place_1383_token : boolean;
  signal place_1384_preds : BooleanArray(0 downto 0);
  signal place_1384_succs : BooleanArray(0 downto 0);
  signal place_1384_token : boolean;
  signal place_1385_preds : BooleanArray(0 downto 0);
  signal place_1385_succs : BooleanArray(0 downto 0);
  signal place_1385_token : boolean;

  signal transition_1_symbol_out : boolean;
  signal transition_1_preds : BooleanArray(0 downto 0);
  signal transition_2_symbol_out : boolean;
  signal transition_2_preds : BooleanArray(0 downto 0);
  signal transition_3_symbol_out : boolean;
  signal transition_3_preds : BooleanArray(1 downto 0);
  signal transition_4_symbol_out : boolean;
  signal transition_4_preds : BooleanArray(0 downto 0);
  signal transition_5_symbol_out : boolean;
  signal transition_5_preds : BooleanArray(1 downto 0);
  signal transition_7_symbol_out : boolean;
  signal transition_7_preds : BooleanArray(0 downto 0);
  signal transition_8_symbol_out : boolean;
  signal transition_8_preds : BooleanArray(0 downto 0);
  signal transition_9_symbol_out : boolean;
  signal transition_9_preds : BooleanArray(0 downto 0);
  signal transition_10_symbol_out : boolean;
  signal transition_10_preds : BooleanArray(1 downto 0);
  signal transition_11_symbol_out : boolean;
  signal transition_11_preds : BooleanArray(0 downto 0);
  signal transition_12_symbol_out : boolean;
  signal transition_12_preds : BooleanArray(1 downto 0);
  signal transition_14_symbol_out : boolean;
  signal transition_14_preds : BooleanArray(0 downto 0);
  signal transition_15_symbol_out : boolean;
  signal transition_15_preds : BooleanArray(0 downto 0);
  signal transition_16_symbol_out : boolean;
  signal transition_16_preds : BooleanArray(0 downto 0);
  signal transition_17_symbol_out : boolean;
  signal transition_17_preds : BooleanArray(0 downto 0);
  signal transition_19_symbol_out : boolean;
  signal transition_19_preds : BooleanArray(0 downto 0);
  signal transition_20_symbol_out : boolean;
  signal transition_20_preds : BooleanArray(0 downto 0);
  signal transition_21_symbol_out : boolean;
  signal transition_21_preds : BooleanArray(0 downto 0);
  signal transition_22_symbol_out : boolean;
  signal transition_22_preds : BooleanArray(0 downto 0);
  signal transition_23_symbol_out : boolean;
  signal transition_23_preds : BooleanArray(0 downto 0);
  signal transition_25_symbol_out : boolean;
  signal transition_25_preds : BooleanArray(0 downto 0);
  signal transition_26_symbol_out : boolean;
  signal transition_26_preds : BooleanArray(0 downto 0);
  signal transition_27_symbol_out : boolean;
  signal transition_27_preds : BooleanArray(0 downto 0);
  signal transition_29_symbol_out : boolean;
  signal transition_29_preds : BooleanArray(0 downto 0);
  signal transition_30_symbol_out : boolean;
  signal transition_30_preds : BooleanArray(0 downto 0);
  signal transition_31_symbol_out : boolean;
  signal transition_31_preds : BooleanArray(0 downto 0);
  signal transition_32_symbol_out : boolean;
  signal transition_32_preds : BooleanArray(0 downto 0);
  signal transition_33_symbol_out : boolean;
  signal transition_33_preds : BooleanArray(0 downto 0);
  signal transition_34_symbol_out : boolean;
  signal transition_34_preds : BooleanArray(0 downto 0);
  signal transition_35_symbol_out : boolean;
  signal transition_35_preds : BooleanArray(0 downto 0);
  signal transition_39_symbol_out : boolean;
  signal transition_39_preds : BooleanArray(0 downto 0);
  signal transition_40_symbol_out : boolean;
  signal transition_40_preds : BooleanArray(0 downto 0);
  signal transition_41_symbol_out : boolean;
  signal transition_41_preds : BooleanArray(0 downto 0);
  signal transition_42_symbol_out : boolean;
  signal transition_42_preds : BooleanArray(0 downto 0);
  signal transition_46_symbol_out : boolean;
  signal transition_46_preds : BooleanArray(0 downto 0);
  signal transition_47_symbol_out : boolean;
  signal transition_47_preds : BooleanArray(0 downto 0);
  signal transition_48_symbol_out : boolean;
  signal transition_48_preds : BooleanArray(0 downto 0);
  signal transition_49_symbol_out : boolean;
  signal transition_49_preds : BooleanArray(0 downto 0);
  signal transition_53_symbol_out : boolean;
  signal transition_53_preds : BooleanArray(1 downto 0);
  signal transition_54_symbol_out : boolean;
  signal transition_54_preds : BooleanArray(0 downto 0);
  signal transition_55_symbol_out : boolean;
  signal transition_55_preds : BooleanArray(0 downto 0);
  signal transition_56_symbol_out : boolean;
  signal transition_56_preds : BooleanArray(0 downto 0);
  signal transition_57_symbol_out : boolean;
  signal transition_57_preds : BooleanArray(0 downto 0);
  signal transition_61_symbol_out : boolean;
  signal transition_61_preds : BooleanArray(0 downto 0);
  signal transition_62_symbol_out : boolean;
  signal transition_62_preds : BooleanArray(0 downto 0);
  signal transition_63_symbol_out : boolean;
  signal transition_63_preds : BooleanArray(0 downto 0);
  signal transition_64_symbol_out : boolean;
  signal transition_64_preds : BooleanArray(0 downto 0);
  signal transition_68_symbol_out : boolean;
  signal transition_68_preds : BooleanArray(1 downto 0);
  signal transition_69_symbol_out : boolean;
  signal transition_69_preds : BooleanArray(0 downto 0);
  signal transition_70_symbol_out : boolean;
  signal transition_70_preds : BooleanArray(0 downto 0);
  signal transition_71_symbol_out : boolean;
  signal transition_71_preds : BooleanArray(0 downto 0);
  signal transition_72_symbol_out : boolean;
  signal transition_72_preds : BooleanArray(0 downto 0);
  signal transition_76_symbol_out : boolean;
  signal transition_76_preds : BooleanArray(0 downto 0);
  signal transition_77_symbol_out : boolean;
  signal transition_77_preds : BooleanArray(0 downto 0);
  signal transition_78_symbol_out : boolean;
  signal transition_78_preds : BooleanArray(0 downto 0);
  signal transition_79_symbol_out : boolean;
  signal transition_79_preds : BooleanArray(0 downto 0);
  signal transition_83_symbol_out : boolean;
  signal transition_83_preds : BooleanArray(0 downto 0);
  signal transition_84_symbol_out : boolean;
  signal transition_84_preds : BooleanArray(0 downto 0);
  signal transition_85_symbol_out : boolean;
  signal transition_85_preds : BooleanArray(0 downto 0);
  signal transition_86_symbol_out : boolean;
  signal transition_86_preds : BooleanArray(0 downto 0);
  signal transition_90_symbol_out : boolean;
  signal transition_90_preds : BooleanArray(0 downto 0);
  signal transition_91_symbol_out : boolean;
  signal transition_91_preds : BooleanArray(0 downto 0);
  signal transition_92_symbol_out : boolean;
  signal transition_92_preds : BooleanArray(0 downto 0);
  signal transition_93_symbol_out : boolean;
  signal transition_93_preds : BooleanArray(0 downto 0);
  signal transition_97_symbol_out : boolean;
  signal transition_97_preds : BooleanArray(1 downto 0);
  signal transition_98_symbol_out : boolean;
  signal transition_98_preds : BooleanArray(0 downto 0);
  signal transition_99_symbol_out : boolean;
  signal transition_99_preds : BooleanArray(0 downto 0);
  signal transition_100_symbol_out : boolean;
  signal transition_100_preds : BooleanArray(0 downto 0);
  signal transition_101_symbol_out : boolean;
  signal transition_101_preds : BooleanArray(0 downto 0);
  signal transition_105_symbol_out : boolean;
  signal transition_105_preds : BooleanArray(0 downto 0);
  signal transition_106_symbol_out : boolean;
  signal transition_106_preds : BooleanArray(0 downto 0);
  signal transition_107_symbol_out : boolean;
  signal transition_107_preds : BooleanArray(0 downto 0);
  signal transition_108_symbol_out : boolean;
  signal transition_108_preds : BooleanArray(0 downto 0);
  signal transition_112_symbol_out : boolean;
  signal transition_112_preds : BooleanArray(1 downto 0);
  signal transition_113_symbol_out : boolean;
  signal transition_113_preds : BooleanArray(0 downto 0);
  signal transition_114_symbol_out : boolean;
  signal transition_114_preds : BooleanArray(0 downto 0);
  signal transition_115_symbol_out : boolean;
  signal transition_115_preds : BooleanArray(0 downto 0);
  signal transition_116_symbol_out : boolean;
  signal transition_116_preds : BooleanArray(0 downto 0);
  signal transition_120_symbol_out : boolean;
  signal transition_120_preds : BooleanArray(0 downto 0);
  signal transition_121_symbol_out : boolean;
  signal transition_121_preds : BooleanArray(0 downto 0);
  signal transition_122_symbol_out : boolean;
  signal transition_122_preds : BooleanArray(0 downto 0);
  signal transition_123_symbol_out : boolean;
  signal transition_123_preds : BooleanArray(0 downto 0);
  signal transition_127_symbol_out : boolean;
  signal transition_127_preds : BooleanArray(0 downto 0);
  signal transition_128_symbol_out : boolean;
  signal transition_128_preds : BooleanArray(0 downto 0);
  signal transition_129_symbol_out : boolean;
  signal transition_129_preds : BooleanArray(0 downto 0);
  signal transition_130_symbol_out : boolean;
  signal transition_130_preds : BooleanArray(0 downto 0);
  signal transition_134_symbol_out : boolean;
  signal transition_134_preds : BooleanArray(0 downto 0);
  signal transition_135_symbol_out : boolean;
  signal transition_135_preds : BooleanArray(0 downto 0);
  signal transition_136_symbol_out : boolean;
  signal transition_136_preds : BooleanArray(0 downto 0);
  signal transition_137_symbol_out : boolean;
  signal transition_137_preds : BooleanArray(0 downto 0);
  signal transition_141_symbol_out : boolean;
  signal transition_141_preds : BooleanArray(1 downto 0);
  signal transition_142_symbol_out : boolean;
  signal transition_142_preds : BooleanArray(0 downto 0);
  signal transition_143_symbol_out : boolean;
  signal transition_143_preds : BooleanArray(0 downto 0);
  signal transition_144_symbol_out : boolean;
  signal transition_144_preds : BooleanArray(0 downto 0);
  signal transition_145_symbol_out : boolean;
  signal transition_145_preds : BooleanArray(0 downto 0);
  signal transition_149_symbol_out : boolean;
  signal transition_149_preds : BooleanArray(0 downto 0);
  signal transition_150_symbol_out : boolean;
  signal transition_150_preds : BooleanArray(0 downto 0);
  signal transition_151_symbol_out : boolean;
  signal transition_151_preds : BooleanArray(0 downto 0);
  signal transition_152_symbol_out : boolean;
  signal transition_152_preds : BooleanArray(0 downto 0);
  signal transition_156_symbol_out : boolean;
  signal transition_156_preds : BooleanArray(0 downto 0);
  signal transition_157_symbol_out : boolean;
  signal transition_157_preds : BooleanArray(0 downto 0);
  signal transition_158_symbol_out : boolean;
  signal transition_158_preds : BooleanArray(0 downto 0);
  signal transition_159_symbol_out : boolean;
  signal transition_159_preds : BooleanArray(0 downto 0);
  signal transition_163_symbol_out : boolean;
  signal transition_163_preds : BooleanArray(1 downto 0);
  signal transition_164_symbol_out : boolean;
  signal transition_164_preds : BooleanArray(0 downto 0);
  signal transition_166_symbol_out : boolean;
  signal transition_166_preds : BooleanArray(0 downto 0);
  signal transition_167_symbol_out : boolean;
  signal transition_167_preds : BooleanArray(0 downto 0);
  signal transition_168_symbol_out : boolean;
  signal transition_168_preds : BooleanArray(2 downto 0);
  signal transition_169_symbol_out : boolean;
  signal transition_169_preds : BooleanArray(0 downto 0);
  signal transition_170_symbol_out : boolean;
  signal transition_170_preds : BooleanArray(0 downto 0);
  signal transition_171_symbol_out : boolean;
  signal transition_171_preds : BooleanArray(0 downto 0);
  signal transition_172_symbol_out : boolean;
  signal transition_172_preds : BooleanArray(0 downto 0);
  signal transition_176_symbol_out : boolean;
  signal transition_176_preds : BooleanArray(0 downto 0);
  signal transition_177_symbol_out : boolean;
  signal transition_177_preds : BooleanArray(0 downto 0);
  signal transition_178_symbol_out : boolean;
  signal transition_178_preds : BooleanArray(0 downto 0);
  signal transition_179_symbol_out : boolean;
  signal transition_179_preds : BooleanArray(0 downto 0);
  signal transition_183_symbol_out : boolean;
  signal transition_183_preds : BooleanArray(0 downto 0);
  signal transition_184_symbol_out : boolean;
  signal transition_184_preds : BooleanArray(0 downto 0);
  signal transition_185_symbol_out : boolean;
  signal transition_185_preds : BooleanArray(0 downto 0);
  signal transition_186_symbol_out : boolean;
  signal transition_186_preds : BooleanArray(0 downto 0);
  signal transition_190_symbol_out : boolean;
  signal transition_190_preds : BooleanArray(1 downto 0);
  signal transition_191_symbol_out : boolean;
  signal transition_191_preds : BooleanArray(0 downto 0);
  signal transition_192_symbol_out : boolean;
  signal transition_192_preds : BooleanArray(0 downto 0);
  signal transition_193_symbol_out : boolean;
  signal transition_193_preds : BooleanArray(0 downto 0);
  signal transition_194_symbol_out : boolean;
  signal transition_194_preds : BooleanArray(0 downto 0);
  signal transition_198_symbol_out : boolean;
  signal transition_198_preds : BooleanArray(0 downto 0);
  signal transition_199_symbol_out : boolean;
  signal transition_199_preds : BooleanArray(0 downto 0);
  signal transition_200_symbol_out : boolean;
  signal transition_200_preds : BooleanArray(0 downto 0);
  signal transition_201_symbol_out : boolean;
  signal transition_201_preds : BooleanArray(0 downto 0);
  signal transition_205_symbol_out : boolean;
  signal transition_205_preds : BooleanArray(0 downto 0);
  signal transition_206_symbol_out : boolean;
  signal transition_206_preds : BooleanArray(0 downto 0);
  signal transition_207_symbol_out : boolean;
  signal transition_207_preds : BooleanArray(0 downto 0);
  signal transition_208_symbol_out : boolean;
  signal transition_208_preds : BooleanArray(0 downto 0);
  signal transition_212_symbol_out : boolean;
  signal transition_212_preds : BooleanArray(1 downto 0);
  signal transition_214_symbol_out : boolean;
  signal transition_214_preds : BooleanArray(0 downto 0);
  signal transition_215_symbol_out : boolean;
  signal transition_215_preds : BooleanArray(0 downto 0);
  signal transition_216_symbol_out : boolean;
  signal transition_216_preds : BooleanArray(2 downto 0);
  signal transition_217_symbol_out : boolean;
  signal transition_217_preds : BooleanArray(0 downto 0);
  signal transition_218_symbol_out : boolean;
  signal transition_218_preds : BooleanArray(0 downto 0);
  signal transition_219_symbol_out : boolean;
  signal transition_219_preds : BooleanArray(0 downto 0);
  signal transition_220_symbol_out : boolean;
  signal transition_220_preds : BooleanArray(0 downto 0);
  signal transition_224_symbol_out : boolean;
  signal transition_224_preds : BooleanArray(0 downto 0);
  signal transition_225_symbol_out : boolean;
  signal transition_225_preds : BooleanArray(0 downto 0);
  signal transition_226_symbol_out : boolean;
  signal transition_226_preds : BooleanArray(0 downto 0);
  signal transition_227_symbol_out : boolean;
  signal transition_227_preds : BooleanArray(0 downto 0);
  signal transition_231_symbol_out : boolean;
  signal transition_231_preds : BooleanArray(0 downto 0);
  signal transition_233_symbol_out : boolean;
  signal transition_233_preds : BooleanArray(0 downto 0);
  signal transition_234_symbol_out : boolean;
  signal transition_234_preds : BooleanArray(0 downto 0);
  signal transition_235_symbol_out : boolean;
  signal transition_235_preds : BooleanArray(0 downto 0);
  signal transition_237_symbol_out : boolean;
  signal transition_237_preds : BooleanArray(0 downto 0);
  signal transition_238_symbol_out : boolean;
  signal transition_238_preds : BooleanArray(0 downto 0);
  signal transition_239_symbol_out : boolean;
  signal transition_239_preds : BooleanArray(0 downto 0);
  signal transition_240_symbol_out : boolean;
  signal transition_240_preds : BooleanArray(0 downto 0);
  signal transition_241_symbol_out : boolean;
  signal transition_241_preds : BooleanArray(0 downto 0);
  signal transition_242_symbol_out : boolean;
  signal transition_242_preds : BooleanArray(0 downto 0);
  signal transition_243_symbol_out : boolean;
  signal transition_243_preds : BooleanArray(0 downto 0);
  signal transition_247_symbol_out : boolean;
  signal transition_247_preds : BooleanArray(0 downto 0);
  signal transition_248_symbol_out : boolean;
  signal transition_248_preds : BooleanArray(0 downto 0);
  signal transition_249_symbol_out : boolean;
  signal transition_249_preds : BooleanArray(0 downto 0);
  signal transition_250_symbol_out : boolean;
  signal transition_250_preds : BooleanArray(0 downto 0);
  signal transition_254_symbol_out : boolean;
  signal transition_254_preds : BooleanArray(0 downto 0);
  signal transition_255_symbol_out : boolean;
  signal transition_255_preds : BooleanArray(0 downto 0);
  signal transition_256_symbol_out : boolean;
  signal transition_256_preds : BooleanArray(0 downto 0);
  signal transition_257_symbol_out : boolean;
  signal transition_257_preds : BooleanArray(0 downto 0);
  signal transition_261_symbol_out : boolean;
  signal transition_261_preds : BooleanArray(1 downto 0);
  signal transition_262_symbol_out : boolean;
  signal transition_262_preds : BooleanArray(0 downto 0);
  signal transition_263_symbol_out : boolean;
  signal transition_263_preds : BooleanArray(0 downto 0);
  signal transition_264_symbol_out : boolean;
  signal transition_264_preds : BooleanArray(0 downto 0);
  signal transition_265_symbol_out : boolean;
  signal transition_265_preds : BooleanArray(0 downto 0);
  signal transition_269_symbol_out : boolean;
  signal transition_269_preds : BooleanArray(0 downto 0);
  signal transition_270_symbol_out : boolean;
  signal transition_270_preds : BooleanArray(0 downto 0);
  signal transition_271_symbol_out : boolean;
  signal transition_271_preds : BooleanArray(0 downto 0);
  signal transition_272_symbol_out : boolean;
  signal transition_272_preds : BooleanArray(0 downto 0);
  signal transition_276_symbol_out : boolean;
  signal transition_276_preds : BooleanArray(1 downto 0);
  signal transition_277_symbol_out : boolean;
  signal transition_277_preds : BooleanArray(0 downto 0);
  signal transition_278_symbol_out : boolean;
  signal transition_278_preds : BooleanArray(0 downto 0);
  signal transition_279_symbol_out : boolean;
  signal transition_279_preds : BooleanArray(0 downto 0);
  signal transition_280_symbol_out : boolean;
  signal transition_280_preds : BooleanArray(0 downto 0);
  signal transition_284_symbol_out : boolean;
  signal transition_284_preds : BooleanArray(0 downto 0);
  signal transition_285_symbol_out : boolean;
  signal transition_285_preds : BooleanArray(0 downto 0);
  signal transition_286_symbol_out : boolean;
  signal transition_286_preds : BooleanArray(0 downto 0);
  signal transition_287_symbol_out : boolean;
  signal transition_287_preds : BooleanArray(0 downto 0);
  signal transition_291_symbol_out : boolean;
  signal transition_291_preds : BooleanArray(0 downto 0);
  signal transition_292_symbol_out : boolean;
  signal transition_292_preds : BooleanArray(0 downto 0);
  signal transition_293_symbol_out : boolean;
  signal transition_293_preds : BooleanArray(0 downto 0);
  signal transition_294_symbol_out : boolean;
  signal transition_294_preds : BooleanArray(0 downto 0);
  signal transition_298_symbol_out : boolean;
  signal transition_298_preds : BooleanArray(0 downto 0);
  signal transition_299_symbol_out : boolean;
  signal transition_299_preds : BooleanArray(0 downto 0);
  signal transition_300_symbol_out : boolean;
  signal transition_300_preds : BooleanArray(0 downto 0);
  signal transition_301_symbol_out : boolean;
  signal transition_301_preds : BooleanArray(0 downto 0);
  signal transition_305_symbol_out : boolean;
  signal transition_305_preds : BooleanArray(1 downto 0);
  signal transition_306_symbol_out : boolean;
  signal transition_306_preds : BooleanArray(0 downto 0);
  signal transition_307_symbol_out : boolean;
  signal transition_307_preds : BooleanArray(0 downto 0);
  signal transition_308_symbol_out : boolean;
  signal transition_308_preds : BooleanArray(0 downto 0);
  signal transition_309_symbol_out : boolean;
  signal transition_309_preds : BooleanArray(0 downto 0);
  signal transition_313_symbol_out : boolean;
  signal transition_313_preds : BooleanArray(0 downto 0);
  signal transition_314_symbol_out : boolean;
  signal transition_314_preds : BooleanArray(0 downto 0);
  signal transition_315_symbol_out : boolean;
  signal transition_315_preds : BooleanArray(0 downto 0);
  signal transition_316_symbol_out : boolean;
  signal transition_316_preds : BooleanArray(0 downto 0);
  signal transition_320_symbol_out : boolean;
  signal transition_320_preds : BooleanArray(1 downto 0);
  signal transition_321_symbol_out : boolean;
  signal transition_321_preds : BooleanArray(0 downto 0);
  signal transition_322_symbol_out : boolean;
  signal transition_322_preds : BooleanArray(0 downto 0);
  signal transition_323_symbol_out : boolean;
  signal transition_323_preds : BooleanArray(0 downto 0);
  signal transition_324_symbol_out : boolean;
  signal transition_324_preds : BooleanArray(0 downto 0);
  signal transition_328_symbol_out : boolean;
  signal transition_328_preds : BooleanArray(0 downto 0);
  signal transition_329_symbol_out : boolean;
  signal transition_329_preds : BooleanArray(0 downto 0);
  signal transition_330_symbol_out : boolean;
  signal transition_330_preds : BooleanArray(0 downto 0);
  signal transition_331_symbol_out : boolean;
  signal transition_331_preds : BooleanArray(0 downto 0);
  signal transition_335_symbol_out : boolean;
  signal transition_335_preds : BooleanArray(0 downto 0);
  signal transition_336_symbol_out : boolean;
  signal transition_336_preds : BooleanArray(0 downto 0);
  signal transition_337_symbol_out : boolean;
  signal transition_337_preds : BooleanArray(0 downto 0);
  signal transition_338_symbol_out : boolean;
  signal transition_338_preds : BooleanArray(0 downto 0);
  signal transition_342_symbol_out : boolean;
  signal transition_342_preds : BooleanArray(0 downto 0);
  signal transition_343_symbol_out : boolean;
  signal transition_343_preds : BooleanArray(0 downto 0);
  signal transition_344_symbol_out : boolean;
  signal transition_344_preds : BooleanArray(0 downto 0);
  signal transition_345_symbol_out : boolean;
  signal transition_345_preds : BooleanArray(0 downto 0);
  signal transition_349_symbol_out : boolean;
  signal transition_349_preds : BooleanArray(1 downto 0);
  signal transition_350_symbol_out : boolean;
  signal transition_350_preds : BooleanArray(0 downto 0);
  signal transition_351_symbol_out : boolean;
  signal transition_351_preds : BooleanArray(0 downto 0);
  signal transition_352_symbol_out : boolean;
  signal transition_352_preds : BooleanArray(0 downto 0);
  signal transition_353_symbol_out : boolean;
  signal transition_353_preds : BooleanArray(0 downto 0);
  signal transition_357_symbol_out : boolean;
  signal transition_357_preds : BooleanArray(0 downto 0);
  signal transition_358_symbol_out : boolean;
  signal transition_358_preds : BooleanArray(0 downto 0);
  signal transition_359_symbol_out : boolean;
  signal transition_359_preds : BooleanArray(0 downto 0);
  signal transition_360_symbol_out : boolean;
  signal transition_360_preds : BooleanArray(0 downto 0);
  signal transition_364_symbol_out : boolean;
  signal transition_364_preds : BooleanArray(0 downto 0);
  signal transition_365_symbol_out : boolean;
  signal transition_365_preds : BooleanArray(0 downto 0);
  signal transition_366_symbol_out : boolean;
  signal transition_366_preds : BooleanArray(0 downto 0);
  signal transition_367_symbol_out : boolean;
  signal transition_367_preds : BooleanArray(0 downto 0);
  signal transition_371_symbol_out : boolean;
  signal transition_371_preds : BooleanArray(1 downto 0);
  signal transition_372_symbol_out : boolean;
  signal transition_372_preds : BooleanArray(0 downto 0);
  signal transition_373_symbol_out : boolean;
  signal transition_373_preds : BooleanArray(0 downto 0);
  signal transition_374_symbol_out : boolean;
  signal transition_374_preds : BooleanArray(0 downto 0);
  signal transition_375_symbol_out : boolean;
  signal transition_375_preds : BooleanArray(0 downto 0);
  signal transition_376_symbol_out : boolean;
  signal transition_376_preds : BooleanArray(0 downto 0);
  signal transition_381_symbol_out : boolean;
  signal transition_381_preds : BooleanArray(0 downto 0);
  signal transition_382_symbol_out : boolean;
  signal transition_382_preds : BooleanArray(0 downto 0);
  signal transition_383_symbol_out : boolean;
  signal transition_383_preds : BooleanArray(2 downto 0);
  signal transition_384_symbol_out : boolean;
  signal transition_384_preds : BooleanArray(0 downto 0);
  signal transition_385_symbol_out : boolean;
  signal transition_385_preds : BooleanArray(0 downto 0);
  signal transition_386_symbol_out : boolean;
  signal transition_386_preds : BooleanArray(0 downto 0);
  signal transition_387_symbol_out : boolean;
  signal transition_387_preds : BooleanArray(0 downto 0);
  signal transition_391_symbol_out : boolean;
  signal transition_391_preds : BooleanArray(0 downto 0);
  signal transition_392_symbol_out : boolean;
  signal transition_392_preds : BooleanArray(0 downto 0);
  signal transition_393_symbol_out : boolean;
  signal transition_393_preds : BooleanArray(0 downto 0);
  signal transition_394_symbol_out : boolean;
  signal transition_394_preds : BooleanArray(0 downto 0);
  signal transition_398_symbol_out : boolean;
  signal transition_398_preds : BooleanArray(0 downto 0);
  signal transition_399_symbol_out : boolean;
  signal transition_399_preds : BooleanArray(0 downto 0);
  signal transition_400_symbol_out : boolean;
  signal transition_400_preds : BooleanArray(0 downto 0);
  signal transition_401_symbol_out : boolean;
  signal transition_401_preds : BooleanArray(0 downto 0);
  signal transition_405_symbol_out : boolean;
  signal transition_405_preds : BooleanArray(1 downto 0);
  signal transition_406_symbol_out : boolean;
  signal transition_406_preds : BooleanArray(0 downto 0);
  signal transition_407_symbol_out : boolean;
  signal transition_407_preds : BooleanArray(0 downto 0);
  signal transition_408_symbol_out : boolean;
  signal transition_408_preds : BooleanArray(0 downto 0);
  signal transition_409_symbol_out : boolean;
  signal transition_409_preds : BooleanArray(0 downto 0);
  signal transition_413_symbol_out : boolean;
  signal transition_413_preds : BooleanArray(0 downto 0);
  signal transition_414_symbol_out : boolean;
  signal transition_414_preds : BooleanArray(0 downto 0);
  signal transition_415_symbol_out : boolean;
  signal transition_415_preds : BooleanArray(0 downto 0);
  signal transition_416_symbol_out : boolean;
  signal transition_416_preds : BooleanArray(0 downto 0);
  signal transition_420_symbol_out : boolean;
  signal transition_420_preds : BooleanArray(0 downto 0);
  signal transition_421_symbol_out : boolean;
  signal transition_421_preds : BooleanArray(0 downto 0);
  signal transition_422_symbol_out : boolean;
  signal transition_422_preds : BooleanArray(0 downto 0);
  signal transition_423_symbol_out : boolean;
  signal transition_423_preds : BooleanArray(0 downto 0);
  signal transition_427_symbol_out : boolean;
  signal transition_427_preds : BooleanArray(1 downto 0);
  signal transition_428_symbol_out : boolean;
  signal transition_428_preds : BooleanArray(0 downto 0);
  signal transition_429_symbol_out : boolean;
  signal transition_429_preds : BooleanArray(0 downto 0);
  signal transition_430_symbol_out : boolean;
  signal transition_430_preds : BooleanArray(0 downto 0);
  signal transition_431_symbol_out : boolean;
  signal transition_431_preds : BooleanArray(0 downto 0);
  signal transition_436_symbol_out : boolean;
  signal transition_436_preds : BooleanArray(0 downto 0);
  signal transition_437_symbol_out : boolean;
  signal transition_437_preds : BooleanArray(0 downto 0);
  signal transition_438_symbol_out : boolean;
  signal transition_438_preds : BooleanArray(2 downto 0);
  signal transition_439_symbol_out : boolean;
  signal transition_439_preds : BooleanArray(0 downto 0);
  signal transition_440_symbol_out : boolean;
  signal transition_440_preds : BooleanArray(0 downto 0);
  signal transition_441_symbol_out : boolean;
  signal transition_441_preds : BooleanArray(0 downto 0);
  signal transition_442_symbol_out : boolean;
  signal transition_442_preds : BooleanArray(0 downto 0);
  signal transition_446_symbol_out : boolean;
  signal transition_446_preds : BooleanArray(0 downto 0);
  signal transition_447_symbol_out : boolean;
  signal transition_447_preds : BooleanArray(0 downto 0);
  signal transition_448_symbol_out : boolean;
  signal transition_448_preds : BooleanArray(0 downto 0);
  signal transition_449_symbol_out : boolean;
  signal transition_449_preds : BooleanArray(0 downto 0);
  signal transition_453_symbol_out : boolean;
  signal transition_453_preds : BooleanArray(0 downto 0);
  signal transition_454_symbol_out : boolean;
  signal transition_454_preds : BooleanArray(0 downto 0);
  signal transition_455_symbol_out : boolean;
  signal transition_455_preds : BooleanArray(0 downto 0);
  signal transition_456_symbol_out : boolean;
  signal transition_456_preds : BooleanArray(0 downto 0);
  signal transition_460_symbol_out : boolean;
  signal transition_460_preds : BooleanArray(0 downto 0);
  signal transition_461_symbol_out : boolean;
  signal transition_461_preds : BooleanArray(0 downto 0);
  signal transition_462_symbol_out : boolean;
  signal transition_462_preds : BooleanArray(0 downto 0);
  signal transition_463_symbol_out : boolean;
  signal transition_463_preds : BooleanArray(0 downto 0);
  signal transition_467_symbol_out : boolean;
  signal transition_467_preds : BooleanArray(0 downto 0);
  signal transition_468_symbol_out : boolean;
  signal transition_468_preds : BooleanArray(0 downto 0);
  signal transition_469_symbol_out : boolean;
  signal transition_469_preds : BooleanArray(0 downto 0);
  signal transition_470_symbol_out : boolean;
  signal transition_470_preds : BooleanArray(0 downto 0);
  signal transition_474_symbol_out : boolean;
  signal transition_474_preds : BooleanArray(1 downto 0);
  signal transition_475_symbol_out : boolean;
  signal transition_475_preds : BooleanArray(0 downto 0);
  signal transition_476_symbol_out : boolean;
  signal transition_476_preds : BooleanArray(0 downto 0);
  signal transition_477_symbol_out : boolean;
  signal transition_477_preds : BooleanArray(0 downto 0);
  signal transition_478_symbol_out : boolean;
  signal transition_478_preds : BooleanArray(0 downto 0);
  signal transition_482_symbol_out : boolean;
  signal transition_482_preds : BooleanArray(0 downto 0);
  signal transition_483_symbol_out : boolean;
  signal transition_483_preds : BooleanArray(0 downto 0);
  signal transition_484_symbol_out : boolean;
  signal transition_484_preds : BooleanArray(0 downto 0);
  signal transition_485_symbol_out : boolean;
  signal transition_485_preds : BooleanArray(0 downto 0);
  signal transition_489_symbol_out : boolean;
  signal transition_489_preds : BooleanArray(1 downto 0);
  signal transition_490_symbol_out : boolean;
  signal transition_490_preds : BooleanArray(0 downto 0);
  signal transition_491_symbol_out : boolean;
  signal transition_491_preds : BooleanArray(0 downto 0);
  signal transition_492_symbol_out : boolean;
  signal transition_492_preds : BooleanArray(0 downto 0);
  signal transition_493_symbol_out : boolean;
  signal transition_493_preds : BooleanArray(0 downto 0);
  signal transition_498_symbol_out : boolean;
  signal transition_498_preds : BooleanArray(0 downto 0);
  signal transition_499_symbol_out : boolean;
  signal transition_499_preds : BooleanArray(0 downto 0);
  signal transition_500_symbol_out : boolean;
  signal transition_500_preds : BooleanArray(1 downto 0);
  signal transition_501_symbol_out : boolean;
  signal transition_501_preds : BooleanArray(0 downto 0);
  signal transition_502_symbol_out : boolean;
  signal transition_502_preds : BooleanArray(0 downto 0);
  signal transition_503_symbol_out : boolean;
  signal transition_503_preds : BooleanArray(0 downto 0);
  signal transition_504_symbol_out : boolean;
  signal transition_504_preds : BooleanArray(0 downto 0);
  signal transition_508_symbol_out : boolean;
  signal transition_508_preds : BooleanArray(0 downto 0);
  signal transition_509_symbol_out : boolean;
  signal transition_509_preds : BooleanArray(0 downto 0);
  signal transition_510_symbol_out : boolean;
  signal transition_510_preds : BooleanArray(0 downto 0);
  signal transition_511_symbol_out : boolean;
  signal transition_511_preds : BooleanArray(0 downto 0);
  signal transition_515_symbol_out : boolean;
  signal transition_515_preds : BooleanArray(0 downto 0);
  signal transition_516_symbol_out : boolean;
  signal transition_516_preds : BooleanArray(0 downto 0);
  signal transition_517_symbol_out : boolean;
  signal transition_517_preds : BooleanArray(0 downto 0);
  signal transition_518_symbol_out : boolean;
  signal transition_518_preds : BooleanArray(0 downto 0);
  signal transition_522_symbol_out : boolean;
  signal transition_522_preds : BooleanArray(1 downto 0);
  signal transition_523_symbol_out : boolean;
  signal transition_523_preds : BooleanArray(0 downto 0);
  signal transition_524_symbol_out : boolean;
  signal transition_524_preds : BooleanArray(0 downto 0);
  signal transition_525_symbol_out : boolean;
  signal transition_525_preds : BooleanArray(0 downto 0);
  signal transition_526_symbol_out : boolean;
  signal transition_526_preds : BooleanArray(0 downto 0);
  signal transition_530_symbol_out : boolean;
  signal transition_530_preds : BooleanArray(0 downto 0);
  signal transition_531_symbol_out : boolean;
  signal transition_531_preds : BooleanArray(0 downto 0);
  signal transition_532_symbol_out : boolean;
  signal transition_532_preds : BooleanArray(0 downto 0);
  signal transition_533_symbol_out : boolean;
  signal transition_533_preds : BooleanArray(0 downto 0);
  signal transition_537_symbol_out : boolean;
  signal transition_537_preds : BooleanArray(1 downto 0);
  signal transition_538_symbol_out : boolean;
  signal transition_538_preds : BooleanArray(0 downto 0);
  signal transition_539_symbol_out : boolean;
  signal transition_539_preds : BooleanArray(0 downto 0);
  signal transition_540_symbol_out : boolean;
  signal transition_540_preds : BooleanArray(0 downto 0);
  signal transition_541_symbol_out : boolean;
  signal transition_541_preds : BooleanArray(0 downto 0);
  signal transition_546_symbol_out : boolean;
  signal transition_546_preds : BooleanArray(0 downto 0);
  signal transition_547_symbol_out : boolean;
  signal transition_547_preds : BooleanArray(0 downto 0);
  signal transition_548_symbol_out : boolean;
  signal transition_548_preds : BooleanArray(1 downto 0);
  signal transition_549_symbol_out : boolean;
  signal transition_549_preds : BooleanArray(0 downto 0);
  signal transition_550_symbol_out : boolean;
  signal transition_550_preds : BooleanArray(0 downto 0);
  signal transition_551_symbol_out : boolean;
  signal transition_551_preds : BooleanArray(0 downto 0);
  signal transition_552_symbol_out : boolean;
  signal transition_552_preds : BooleanArray(0 downto 0);
  signal transition_556_symbol_out : boolean;
  signal transition_556_preds : BooleanArray(0 downto 0);
  signal transition_557_symbol_out : boolean;
  signal transition_557_preds : BooleanArray(0 downto 0);
  signal transition_558_symbol_out : boolean;
  signal transition_558_preds : BooleanArray(0 downto 0);
  signal transition_559_symbol_out : boolean;
  signal transition_559_preds : BooleanArray(0 downto 0);
  signal transition_563_symbol_out : boolean;
  signal transition_563_preds : BooleanArray(0 downto 0);
  signal transition_564_symbol_out : boolean;
  signal transition_564_preds : BooleanArray(0 downto 0);
  signal transition_565_symbol_out : boolean;
  signal transition_565_preds : BooleanArray(0 downto 0);
  signal transition_566_symbol_out : boolean;
  signal transition_566_preds : BooleanArray(0 downto 0);
  signal transition_570_symbol_out : boolean;
  signal transition_570_preds : BooleanArray(1 downto 0);
  signal transition_571_symbol_out : boolean;
  signal transition_571_preds : BooleanArray(0 downto 0);
  signal transition_572_symbol_out : boolean;
  signal transition_572_preds : BooleanArray(0 downto 0);
  signal transition_573_symbol_out : boolean;
  signal transition_573_preds : BooleanArray(0 downto 0);
  signal transition_574_symbol_out : boolean;
  signal transition_574_preds : BooleanArray(0 downto 0);
  signal transition_578_symbol_out : boolean;
  signal transition_578_preds : BooleanArray(0 downto 0);
  signal transition_579_symbol_out : boolean;
  signal transition_579_preds : BooleanArray(0 downto 0);
  signal transition_580_symbol_out : boolean;
  signal transition_580_preds : BooleanArray(0 downto 0);
  signal transition_581_symbol_out : boolean;
  signal transition_581_preds : BooleanArray(0 downto 0);
  signal transition_585_symbol_out : boolean;
  signal transition_585_preds : BooleanArray(1 downto 0);
  signal transition_586_symbol_out : boolean;
  signal transition_586_preds : BooleanArray(0 downto 0);
  signal transition_587_symbol_out : boolean;
  signal transition_587_preds : BooleanArray(0 downto 0);
  signal transition_588_symbol_out : boolean;
  signal transition_588_preds : BooleanArray(0 downto 0);
  signal transition_589_symbol_out : boolean;
  signal transition_589_preds : BooleanArray(0 downto 0);
  signal transition_594_symbol_out : boolean;
  signal transition_594_preds : BooleanArray(0 downto 0);
  signal transition_595_symbol_out : boolean;
  signal transition_595_preds : BooleanArray(0 downto 0);
  signal transition_596_symbol_out : boolean;
  signal transition_596_preds : BooleanArray(1 downto 0);
  signal transition_597_symbol_out : boolean;
  signal transition_597_preds : BooleanArray(0 downto 0);
  signal transition_598_symbol_out : boolean;
  signal transition_598_preds : BooleanArray(0 downto 0);
  signal transition_599_symbol_out : boolean;
  signal transition_599_preds : BooleanArray(0 downto 0);
  signal transition_600_symbol_out : boolean;
  signal transition_600_preds : BooleanArray(0 downto 0);
  signal transition_604_symbol_out : boolean;
  signal transition_604_preds : BooleanArray(0 downto 0);
  signal transition_605_symbol_out : boolean;
  signal transition_605_preds : BooleanArray(0 downto 0);
  signal transition_606_symbol_out : boolean;
  signal transition_606_preds : BooleanArray(0 downto 0);
  signal transition_607_symbol_out : boolean;
  signal transition_607_preds : BooleanArray(0 downto 0);
  signal transition_611_symbol_out : boolean;
  signal transition_611_preds : BooleanArray(0 downto 0);
  signal transition_612_symbol_out : boolean;
  signal transition_612_preds : BooleanArray(0 downto 0);
  signal transition_613_symbol_out : boolean;
  signal transition_613_preds : BooleanArray(0 downto 0);
  signal transition_614_symbol_out : boolean;
  signal transition_614_preds : BooleanArray(0 downto 0);
  signal transition_618_symbol_out : boolean;
  signal transition_618_preds : BooleanArray(1 downto 0);
  signal transition_619_symbol_out : boolean;
  signal transition_619_preds : BooleanArray(0 downto 0);
  signal transition_620_symbol_out : boolean;
  signal transition_620_preds : BooleanArray(0 downto 0);
  signal transition_621_symbol_out : boolean;
  signal transition_621_preds : BooleanArray(0 downto 0);
  signal transition_622_symbol_out : boolean;
  signal transition_622_preds : BooleanArray(0 downto 0);
  signal transition_626_symbol_out : boolean;
  signal transition_626_preds : BooleanArray(0 downto 0);
  signal transition_627_symbol_out : boolean;
  signal transition_627_preds : BooleanArray(0 downto 0);
  signal transition_628_symbol_out : boolean;
  signal transition_628_preds : BooleanArray(0 downto 0);
  signal transition_629_symbol_out : boolean;
  signal transition_629_preds : BooleanArray(0 downto 0);
  signal transition_633_symbol_out : boolean;
  signal transition_633_preds : BooleanArray(1 downto 0);
  signal transition_634_symbol_out : boolean;
  signal transition_634_preds : BooleanArray(0 downto 0);
  signal transition_635_symbol_out : boolean;
  signal transition_635_preds : BooleanArray(0 downto 0);
  signal transition_636_symbol_out : boolean;
  signal transition_636_preds : BooleanArray(0 downto 0);
  signal transition_637_symbol_out : boolean;
  signal transition_637_preds : BooleanArray(0 downto 0);
  signal transition_642_symbol_out : boolean;
  signal transition_642_preds : BooleanArray(0 downto 0);
  signal transition_643_symbol_out : boolean;
  signal transition_643_preds : BooleanArray(0 downto 0);
  signal transition_644_symbol_out : boolean;
  signal transition_644_preds : BooleanArray(1 downto 0);
  signal transition_645_symbol_out : boolean;
  signal transition_645_preds : BooleanArray(0 downto 0);
  signal transition_646_symbol_out : boolean;
  signal transition_646_preds : BooleanArray(0 downto 0);
  signal transition_647_symbol_out : boolean;
  signal transition_647_preds : BooleanArray(0 downto 0);
  signal transition_648_symbol_out : boolean;
  signal transition_648_preds : BooleanArray(0 downto 0);
  signal transition_652_symbol_out : boolean;
  signal transition_652_preds : BooleanArray(0 downto 0);
  signal transition_653_symbol_out : boolean;
  signal transition_653_preds : BooleanArray(0 downto 0);
  signal transition_654_symbol_out : boolean;
  signal transition_654_preds : BooleanArray(0 downto 0);
  signal transition_655_symbol_out : boolean;
  signal transition_655_preds : BooleanArray(0 downto 0);
  signal transition_659_symbol_out : boolean;
  signal transition_659_preds : BooleanArray(0 downto 0);
  signal transition_660_symbol_out : boolean;
  signal transition_660_preds : BooleanArray(0 downto 0);
  signal transition_661_symbol_out : boolean;
  signal transition_661_preds : BooleanArray(0 downto 0);
  signal transition_662_symbol_out : boolean;
  signal transition_662_preds : BooleanArray(0 downto 0);
  signal transition_666_symbol_out : boolean;
  signal transition_666_preds : BooleanArray(1 downto 0);
  signal transition_667_symbol_out : boolean;
  signal transition_667_preds : BooleanArray(0 downto 0);
  signal transition_668_symbol_out : boolean;
  signal transition_668_preds : BooleanArray(0 downto 0);
  signal transition_669_symbol_out : boolean;
  signal transition_669_preds : BooleanArray(0 downto 0);
  signal transition_670_symbol_out : boolean;
  signal transition_670_preds : BooleanArray(0 downto 0);
  signal transition_674_symbol_out : boolean;
  signal transition_674_preds : BooleanArray(0 downto 0);
  signal transition_675_symbol_out : boolean;
  signal transition_675_preds : BooleanArray(0 downto 0);
  signal transition_676_symbol_out : boolean;
  signal transition_676_preds : BooleanArray(0 downto 0);
  signal transition_677_symbol_out : boolean;
  signal transition_677_preds : BooleanArray(0 downto 0);
  signal transition_681_symbol_out : boolean;
  signal transition_681_preds : BooleanArray(1 downto 0);
  signal transition_682_symbol_out : boolean;
  signal transition_682_preds : BooleanArray(0 downto 0);
  signal transition_683_symbol_out : boolean;
  signal transition_683_preds : BooleanArray(0 downto 0);
  signal transition_684_symbol_out : boolean;
  signal transition_684_preds : BooleanArray(0 downto 0);
  signal transition_685_symbol_out : boolean;
  signal transition_685_preds : BooleanArray(0 downto 0);
  signal transition_690_symbol_out : boolean;
  signal transition_690_preds : BooleanArray(0 downto 0);
  signal transition_691_symbol_out : boolean;
  signal transition_691_preds : BooleanArray(0 downto 0);
  signal transition_692_symbol_out : boolean;
  signal transition_692_preds : BooleanArray(1 downto 0);
  signal transition_693_symbol_out : boolean;
  signal transition_693_preds : BooleanArray(0 downto 0);
  signal transition_694_symbol_out : boolean;
  signal transition_694_preds : BooleanArray(0 downto 0);
  signal transition_695_symbol_out : boolean;
  signal transition_695_preds : BooleanArray(0 downto 0);
  signal transition_696_symbol_out : boolean;
  signal transition_696_preds : BooleanArray(0 downto 0);
  signal transition_700_symbol_out : boolean;
  signal transition_700_preds : BooleanArray(0 downto 0);
  signal transition_701_symbol_out : boolean;
  signal transition_701_preds : BooleanArray(0 downto 0);
  signal transition_702_symbol_out : boolean;
  signal transition_702_preds : BooleanArray(0 downto 0);
  signal transition_703_symbol_out : boolean;
  signal transition_703_preds : BooleanArray(0 downto 0);
  signal transition_707_symbol_out : boolean;
  signal transition_707_preds : BooleanArray(0 downto 0);
  signal transition_708_symbol_out : boolean;
  signal transition_708_preds : BooleanArray(0 downto 0);
  signal transition_709_symbol_out : boolean;
  signal transition_709_preds : BooleanArray(0 downto 0);
  signal transition_710_symbol_out : boolean;
  signal transition_710_preds : BooleanArray(0 downto 0);
  signal transition_714_symbol_out : boolean;
  signal transition_714_preds : BooleanArray(1 downto 0);
  signal transition_715_symbol_out : boolean;
  signal transition_715_preds : BooleanArray(0 downto 0);
  signal transition_716_symbol_out : boolean;
  signal transition_716_preds : BooleanArray(0 downto 0);
  signal transition_717_symbol_out : boolean;
  signal transition_717_preds : BooleanArray(0 downto 0);
  signal transition_718_symbol_out : boolean;
  signal transition_718_preds : BooleanArray(0 downto 0);
  signal transition_722_symbol_out : boolean;
  signal transition_722_preds : BooleanArray(0 downto 0);
  signal transition_723_symbol_out : boolean;
  signal transition_723_preds : BooleanArray(0 downto 0);
  signal transition_724_symbol_out : boolean;
  signal transition_724_preds : BooleanArray(0 downto 0);
  signal transition_725_symbol_out : boolean;
  signal transition_725_preds : BooleanArray(0 downto 0);
  signal transition_729_symbol_out : boolean;
  signal transition_729_preds : BooleanArray(1 downto 0);
  signal transition_730_symbol_out : boolean;
  signal transition_730_preds : BooleanArray(0 downto 0);
  signal transition_731_symbol_out : boolean;
  signal transition_731_preds : BooleanArray(0 downto 0);
  signal transition_732_symbol_out : boolean;
  signal transition_732_preds : BooleanArray(0 downto 0);
  signal transition_733_symbol_out : boolean;
  signal transition_733_preds : BooleanArray(0 downto 0);
  signal transition_738_symbol_out : boolean;
  signal transition_738_preds : BooleanArray(0 downto 0);
  signal transition_739_symbol_out : boolean;
  signal transition_739_preds : BooleanArray(0 downto 0);
  signal transition_740_symbol_out : boolean;
  signal transition_740_preds : BooleanArray(1 downto 0);
  signal transition_741_symbol_out : boolean;
  signal transition_741_preds : BooleanArray(0 downto 0);
  signal transition_742_symbol_out : boolean;
  signal transition_742_preds : BooleanArray(0 downto 0);
  signal transition_743_symbol_out : boolean;
  signal transition_743_preds : BooleanArray(0 downto 0);
  signal transition_744_symbol_out : boolean;
  signal transition_744_preds : BooleanArray(0 downto 0);
  signal transition_748_symbol_out : boolean;
  signal transition_748_preds : BooleanArray(0 downto 0);
  signal transition_749_symbol_out : boolean;
  signal transition_749_preds : BooleanArray(0 downto 0);
  signal transition_750_symbol_out : boolean;
  signal transition_750_preds : BooleanArray(0 downto 0);
  signal transition_751_symbol_out : boolean;
  signal transition_751_preds : BooleanArray(0 downto 0);
  signal transition_755_symbol_out : boolean;
  signal transition_755_preds : BooleanArray(0 downto 0);
  signal transition_756_symbol_out : boolean;
  signal transition_756_preds : BooleanArray(0 downto 0);
  signal transition_757_symbol_out : boolean;
  signal transition_757_preds : BooleanArray(0 downto 0);
  signal transition_758_symbol_out : boolean;
  signal transition_758_preds : BooleanArray(0 downto 0);
  signal transition_762_symbol_out : boolean;
  signal transition_762_preds : BooleanArray(1 downto 0);
  signal transition_763_symbol_out : boolean;
  signal transition_763_preds : BooleanArray(0 downto 0);
  signal transition_764_symbol_out : boolean;
  signal transition_764_preds : BooleanArray(0 downto 0);
  signal transition_765_symbol_out : boolean;
  signal transition_765_preds : BooleanArray(0 downto 0);
  signal transition_766_symbol_out : boolean;
  signal transition_766_preds : BooleanArray(0 downto 0);
  signal transition_770_symbol_out : boolean;
  signal transition_770_preds : BooleanArray(0 downto 0);
  signal transition_771_symbol_out : boolean;
  signal transition_771_preds : BooleanArray(0 downto 0);
  signal transition_772_symbol_out : boolean;
  signal transition_772_preds : BooleanArray(0 downto 0);
  signal transition_773_symbol_out : boolean;
  signal transition_773_preds : BooleanArray(0 downto 0);
  signal transition_777_symbol_out : boolean;
  signal transition_777_preds : BooleanArray(1 downto 0);
  signal transition_778_symbol_out : boolean;
  signal transition_778_preds : BooleanArray(0 downto 0);
  signal transition_779_symbol_out : boolean;
  signal transition_779_preds : BooleanArray(0 downto 0);
  signal transition_780_symbol_out : boolean;
  signal transition_780_preds : BooleanArray(0 downto 0);
  signal transition_781_symbol_out : boolean;
  signal transition_781_preds : BooleanArray(0 downto 0);
  signal transition_786_symbol_out : boolean;
  signal transition_786_preds : BooleanArray(0 downto 0);
  signal transition_787_symbol_out : boolean;
  signal transition_787_preds : BooleanArray(0 downto 0);
  signal transition_788_symbol_out : boolean;
  signal transition_788_preds : BooleanArray(1 downto 0);
  signal transition_789_symbol_out : boolean;
  signal transition_789_preds : BooleanArray(0 downto 0);
  signal transition_790_symbol_out : boolean;
  signal transition_790_preds : BooleanArray(0 downto 0);
  signal transition_791_symbol_out : boolean;
  signal transition_791_preds : BooleanArray(0 downto 0);
  signal transition_792_symbol_out : boolean;
  signal transition_792_preds : BooleanArray(0 downto 0);
  signal transition_796_symbol_out : boolean;
  signal transition_796_preds : BooleanArray(0 downto 0);
  signal transition_797_symbol_out : boolean;
  signal transition_797_preds : BooleanArray(0 downto 0);
  signal transition_798_symbol_out : boolean;
  signal transition_798_preds : BooleanArray(0 downto 0);
  signal transition_799_symbol_out : boolean;
  signal transition_799_preds : BooleanArray(0 downto 0);
  signal transition_803_symbol_out : boolean;
  signal transition_803_preds : BooleanArray(0 downto 0);
  signal transition_804_symbol_out : boolean;
  signal transition_804_preds : BooleanArray(0 downto 0);
  signal transition_805_symbol_out : boolean;
  signal transition_805_preds : BooleanArray(0 downto 0);
  signal transition_806_symbol_out : boolean;
  signal transition_806_preds : BooleanArray(0 downto 0);
  signal transition_810_symbol_out : boolean;
  signal transition_810_preds : BooleanArray(1 downto 0);
  signal transition_811_symbol_out : boolean;
  signal transition_811_preds : BooleanArray(0 downto 0);
  signal transition_812_symbol_out : boolean;
  signal transition_812_preds : BooleanArray(0 downto 0);
  signal transition_813_symbol_out : boolean;
  signal transition_813_preds : BooleanArray(0 downto 0);
  signal transition_814_symbol_out : boolean;
  signal transition_814_preds : BooleanArray(0 downto 0);
  signal transition_818_symbol_out : boolean;
  signal transition_818_preds : BooleanArray(0 downto 0);
  signal transition_819_symbol_out : boolean;
  signal transition_819_preds : BooleanArray(0 downto 0);
  signal transition_820_symbol_out : boolean;
  signal transition_820_preds : BooleanArray(0 downto 0);
  signal transition_821_symbol_out : boolean;
  signal transition_821_preds : BooleanArray(0 downto 0);
  signal transition_825_symbol_out : boolean;
  signal transition_825_preds : BooleanArray(1 downto 0);
  signal transition_826_symbol_out : boolean;
  signal transition_826_preds : BooleanArray(0 downto 0);
  signal transition_827_symbol_out : boolean;
  signal transition_827_preds : BooleanArray(0 downto 0);
  signal transition_828_symbol_out : boolean;
  signal transition_828_preds : BooleanArray(0 downto 0);
  signal transition_829_symbol_out : boolean;
  signal transition_829_preds : BooleanArray(0 downto 0);
  signal transition_834_symbol_out : boolean;
  signal transition_834_preds : BooleanArray(0 downto 0);
  signal transition_835_symbol_out : boolean;
  signal transition_835_preds : BooleanArray(0 downto 0);
  signal transition_836_symbol_out : boolean;
  signal transition_836_preds : BooleanArray(1 downto 0);
  signal transition_837_symbol_out : boolean;
  signal transition_837_preds : BooleanArray(0 downto 0);
  signal transition_838_symbol_out : boolean;
  signal transition_838_preds : BooleanArray(0 downto 0);
  signal transition_839_symbol_out : boolean;
  signal transition_839_preds : BooleanArray(0 downto 0);
  signal transition_840_symbol_out : boolean;
  signal transition_840_preds : BooleanArray(0 downto 0);
  signal transition_844_symbol_out : boolean;
  signal transition_844_preds : BooleanArray(0 downto 0);
  signal transition_845_symbol_out : boolean;
  signal transition_845_preds : BooleanArray(0 downto 0);
  signal transition_846_symbol_out : boolean;
  signal transition_846_preds : BooleanArray(0 downto 0);
  signal transition_847_symbol_out : boolean;
  signal transition_847_preds : BooleanArray(0 downto 0);
  signal transition_851_symbol_out : boolean;
  signal transition_851_preds : BooleanArray(0 downto 0);
  signal transition_852_symbol_out : boolean;
  signal transition_852_preds : BooleanArray(0 downto 0);
  signal transition_853_symbol_out : boolean;
  signal transition_853_preds : BooleanArray(0 downto 0);
  signal transition_854_symbol_out : boolean;
  signal transition_854_preds : BooleanArray(0 downto 0);
  signal transition_858_symbol_out : boolean;
  signal transition_858_preds : BooleanArray(1 downto 0);
  signal transition_859_symbol_out : boolean;
  signal transition_859_preds : BooleanArray(0 downto 0);
  signal transition_860_symbol_out : boolean;
  signal transition_860_preds : BooleanArray(0 downto 0);
  signal transition_861_symbol_out : boolean;
  signal transition_861_preds : BooleanArray(0 downto 0);
  signal transition_862_symbol_out : boolean;
  signal transition_862_preds : BooleanArray(0 downto 0);
  signal transition_866_symbol_out : boolean;
  signal transition_866_preds : BooleanArray(0 downto 0);
  signal transition_867_symbol_out : boolean;
  signal transition_867_preds : BooleanArray(0 downto 0);
  signal transition_868_symbol_out : boolean;
  signal transition_868_preds : BooleanArray(0 downto 0);
  signal transition_869_symbol_out : boolean;
  signal transition_869_preds : BooleanArray(0 downto 0);
  signal transition_873_symbol_out : boolean;
  signal transition_873_preds : BooleanArray(1 downto 0);
  signal transition_874_symbol_out : boolean;
  signal transition_874_preds : BooleanArray(0 downto 0);
  signal transition_875_symbol_out : boolean;
  signal transition_875_preds : BooleanArray(0 downto 0);
  signal transition_876_symbol_out : boolean;
  signal transition_876_preds : BooleanArray(0 downto 0);
  signal transition_877_symbol_out : boolean;
  signal transition_877_preds : BooleanArray(0 downto 0);
  signal transition_882_symbol_out : boolean;
  signal transition_882_preds : BooleanArray(0 downto 0);
  signal transition_883_symbol_out : boolean;
  signal transition_883_preds : BooleanArray(0 downto 0);
  signal transition_884_symbol_out : boolean;
  signal transition_884_preds : BooleanArray(1 downto 0);
  signal transition_885_symbol_out : boolean;
  signal transition_885_preds : BooleanArray(0 downto 0);
  signal transition_886_symbol_out : boolean;
  signal transition_886_preds : BooleanArray(0 downto 0);
  signal transition_887_symbol_out : boolean;
  signal transition_887_preds : BooleanArray(0 downto 0);
  signal transition_888_symbol_out : boolean;
  signal transition_888_preds : BooleanArray(0 downto 0);
  signal transition_892_symbol_out : boolean;
  signal transition_892_preds : BooleanArray(0 downto 0);
  signal transition_893_symbol_out : boolean;
  signal transition_893_preds : BooleanArray(0 downto 0);
  signal transition_894_symbol_out : boolean;
  signal transition_894_preds : BooleanArray(0 downto 0);
  signal transition_895_symbol_out : boolean;
  signal transition_895_preds : BooleanArray(0 downto 0);
  signal transition_899_symbol_out : boolean;
  signal transition_899_preds : BooleanArray(0 downto 0);
  signal transition_900_symbol_out : boolean;
  signal transition_900_preds : BooleanArray(0 downto 0);
  signal transition_901_symbol_out : boolean;
  signal transition_901_preds : BooleanArray(0 downto 0);
  signal transition_902_symbol_out : boolean;
  signal transition_902_preds : BooleanArray(0 downto 0);
  signal transition_906_symbol_out : boolean;
  signal transition_906_preds : BooleanArray(1 downto 0);
  signal transition_907_symbol_out : boolean;
  signal transition_907_preds : BooleanArray(0 downto 0);
  signal transition_908_symbol_out : boolean;
  signal transition_908_preds : BooleanArray(0 downto 0);
  signal transition_909_symbol_out : boolean;
  signal transition_909_preds : BooleanArray(0 downto 0);
  signal transition_910_symbol_out : boolean;
  signal transition_910_preds : BooleanArray(0 downto 0);
  signal transition_914_symbol_out : boolean;
  signal transition_914_preds : BooleanArray(0 downto 0);
  signal transition_915_symbol_out : boolean;
  signal transition_915_preds : BooleanArray(0 downto 0);
  signal transition_916_symbol_out : boolean;
  signal transition_916_preds : BooleanArray(0 downto 0);
  signal transition_917_symbol_out : boolean;
  signal transition_917_preds : BooleanArray(0 downto 0);
  signal transition_921_symbol_out : boolean;
  signal transition_921_preds : BooleanArray(1 downto 0);
  signal transition_922_symbol_out : boolean;
  signal transition_922_preds : BooleanArray(0 downto 0);
  signal transition_923_symbol_out : boolean;
  signal transition_923_preds : BooleanArray(0 downto 0);
  signal transition_924_symbol_out : boolean;
  signal transition_924_preds : BooleanArray(0 downto 0);
  signal transition_925_symbol_out : boolean;
  signal transition_925_preds : BooleanArray(0 downto 0);
  signal transition_930_symbol_out : boolean;
  signal transition_930_preds : BooleanArray(0 downto 0);
  signal transition_931_symbol_out : boolean;
  signal transition_931_preds : BooleanArray(0 downto 0);
  signal transition_932_symbol_out : boolean;
  signal transition_932_preds : BooleanArray(1 downto 0);
  signal transition_933_symbol_out : boolean;
  signal transition_933_preds : BooleanArray(0 downto 0);
  signal transition_934_symbol_out : boolean;
  signal transition_934_preds : BooleanArray(0 downto 0);
  signal transition_935_symbol_out : boolean;
  signal transition_935_preds : BooleanArray(0 downto 0);
  signal transition_936_symbol_out : boolean;
  signal transition_936_preds : BooleanArray(0 downto 0);
  signal transition_940_symbol_out : boolean;
  signal transition_940_preds : BooleanArray(0 downto 0);
  signal transition_941_symbol_out : boolean;
  signal transition_941_preds : BooleanArray(0 downto 0);
  signal transition_942_symbol_out : boolean;
  signal transition_942_preds : BooleanArray(0 downto 0);
  signal transition_943_symbol_out : boolean;
  signal transition_943_preds : BooleanArray(0 downto 0);
  signal transition_947_symbol_out : boolean;
  signal transition_947_preds : BooleanArray(0 downto 0);
  signal transition_948_symbol_out : boolean;
  signal transition_948_preds : BooleanArray(0 downto 0);
  signal transition_949_symbol_out : boolean;
  signal transition_949_preds : BooleanArray(0 downto 0);
  signal transition_950_symbol_out : boolean;
  signal transition_950_preds : BooleanArray(0 downto 0);
  signal transition_954_symbol_out : boolean;
  signal transition_954_preds : BooleanArray(1 downto 0);
  signal transition_955_symbol_out : boolean;
  signal transition_955_preds : BooleanArray(0 downto 0);
  signal transition_956_symbol_out : boolean;
  signal transition_956_preds : BooleanArray(0 downto 0);
  signal transition_957_symbol_out : boolean;
  signal transition_957_preds : BooleanArray(0 downto 0);
  signal transition_958_symbol_out : boolean;
  signal transition_958_preds : BooleanArray(0 downto 0);
  signal transition_962_symbol_out : boolean;
  signal transition_962_preds : BooleanArray(0 downto 0);
  signal transition_963_symbol_out : boolean;
  signal transition_963_preds : BooleanArray(0 downto 0);
  signal transition_964_symbol_out : boolean;
  signal transition_964_preds : BooleanArray(0 downto 0);
  signal transition_965_symbol_out : boolean;
  signal transition_965_preds : BooleanArray(0 downto 0);
  signal transition_969_symbol_out : boolean;
  signal transition_969_preds : BooleanArray(1 downto 0);
  signal transition_970_symbol_out : boolean;
  signal transition_970_preds : BooleanArray(0 downto 0);
  signal transition_971_symbol_out : boolean;
  signal transition_971_preds : BooleanArray(0 downto 0);
  signal transition_972_symbol_out : boolean;
  signal transition_972_preds : BooleanArray(0 downto 0);
  signal transition_973_symbol_out : boolean;
  signal transition_973_preds : BooleanArray(0 downto 0);
  signal transition_978_symbol_out : boolean;
  signal transition_978_preds : BooleanArray(0 downto 0);
  signal transition_979_symbol_out : boolean;
  signal transition_979_preds : BooleanArray(0 downto 0);
  signal transition_980_symbol_out : boolean;
  signal transition_980_preds : BooleanArray(1 downto 0);
  signal transition_981_symbol_out : boolean;
  signal transition_981_preds : BooleanArray(0 downto 0);
  signal transition_982_symbol_out : boolean;
  signal transition_982_preds : BooleanArray(0 downto 0);
  signal transition_983_symbol_out : boolean;
  signal transition_983_preds : BooleanArray(0 downto 0);
  signal transition_984_symbol_out : boolean;
  signal transition_984_preds : BooleanArray(0 downto 0);
  signal transition_988_symbol_out : boolean;
  signal transition_988_preds : BooleanArray(0 downto 0);
  signal transition_989_symbol_out : boolean;
  signal transition_989_preds : BooleanArray(0 downto 0);
  signal transition_990_symbol_out : boolean;
  signal transition_990_preds : BooleanArray(0 downto 0);
  signal transition_991_symbol_out : boolean;
  signal transition_991_preds : BooleanArray(0 downto 0);
  signal transition_995_symbol_out : boolean;
  signal transition_995_preds : BooleanArray(0 downto 0);
  signal transition_996_symbol_out : boolean;
  signal transition_996_preds : BooleanArray(0 downto 0);
  signal transition_997_symbol_out : boolean;
  signal transition_997_preds : BooleanArray(0 downto 0);
  signal transition_998_symbol_out : boolean;
  signal transition_998_preds : BooleanArray(0 downto 0);
  signal transition_1002_symbol_out : boolean;
  signal transition_1002_preds : BooleanArray(1 downto 0);
  signal transition_1003_symbol_out : boolean;
  signal transition_1003_preds : BooleanArray(0 downto 0);
  signal transition_1004_symbol_out : boolean;
  signal transition_1004_preds : BooleanArray(0 downto 0);
  signal transition_1005_symbol_out : boolean;
  signal transition_1005_preds : BooleanArray(0 downto 0);
  signal transition_1006_symbol_out : boolean;
  signal transition_1006_preds : BooleanArray(0 downto 0);
  signal transition_1010_symbol_out : boolean;
  signal transition_1010_preds : BooleanArray(0 downto 0);
  signal transition_1011_symbol_out : boolean;
  signal transition_1011_preds : BooleanArray(0 downto 0);
  signal transition_1012_symbol_out : boolean;
  signal transition_1012_preds : BooleanArray(0 downto 0);
  signal transition_1013_symbol_out : boolean;
  signal transition_1013_preds : BooleanArray(0 downto 0);
  signal transition_1017_symbol_out : boolean;
  signal transition_1017_preds : BooleanArray(1 downto 0);
  signal transition_1018_symbol_out : boolean;
  signal transition_1018_preds : BooleanArray(0 downto 0);
  signal transition_1019_symbol_out : boolean;
  signal transition_1019_preds : BooleanArray(0 downto 0);
  signal transition_1020_symbol_out : boolean;
  signal transition_1020_preds : BooleanArray(0 downto 0);
  signal transition_1021_symbol_out : boolean;
  signal transition_1021_preds : BooleanArray(0 downto 0);
  signal transition_1026_symbol_out : boolean;
  signal transition_1026_preds : BooleanArray(0 downto 0);
  signal transition_1027_symbol_out : boolean;
  signal transition_1027_preds : BooleanArray(0 downto 0);
  signal transition_1028_symbol_out : boolean;
  signal transition_1028_preds : BooleanArray(1 downto 0);
  signal transition_1030_symbol_out : boolean;
  signal transition_1030_preds : BooleanArray(0 downto 0);
  signal transition_1031_symbol_out : boolean;
  signal transition_1031_preds : BooleanArray(0 downto 0);
  signal transition_1033_symbol_out : boolean;
  signal transition_1033_preds : BooleanArray(0 downto 0);
  signal transition_1034_symbol_out : boolean;
  signal transition_1034_preds : BooleanArray(0 downto 0);
  signal transition_1035_symbol_out : boolean;
  signal transition_1035_preds : BooleanArray(0 downto 0);
  signal transition_1037_symbol_out : boolean;
  signal transition_1037_preds : BooleanArray(0 downto 0);
  signal transition_1038_symbol_out : boolean;
  signal transition_1038_preds : BooleanArray(0 downto 0);
  signal transition_1040_symbol_out : boolean;
  signal transition_1040_preds : BooleanArray(0 downto 0);
  signal transition_1041_symbol_out : boolean;
  signal transition_1041_preds : BooleanArray(0 downto 0);
  signal transition_1042_symbol_out : boolean;
  signal transition_1042_preds : BooleanArray(0 downto 0);
  signal transition_1043_symbol_out : boolean;
  signal transition_1043_preds : BooleanArray(0 downto 0);
  signal transition_1044_symbol_out : boolean;
  signal transition_1044_preds : BooleanArray(0 downto 0);
  signal transition_1045_symbol_out : boolean;
  signal transition_1045_preds : BooleanArray(0 downto 0);
  signal transition_1046_symbol_out : boolean;
  signal transition_1046_preds : BooleanArray(0 downto 0);
  signal transition_1051_symbol_out : boolean;
  signal transition_1051_preds : BooleanArray(0 downto 0);
  signal transition_1052_symbol_out : boolean;
  signal transition_1052_preds : BooleanArray(0 downto 0);
  signal transition_1054_symbol_out : boolean;
  signal transition_1054_preds : BooleanArray(0 downto 0);
  signal transition_1055_symbol_out : boolean;
  signal transition_1055_preds : BooleanArray(0 downto 0);
  signal transition_1056_symbol_out : boolean;
  signal transition_1056_preds : BooleanArray(0 downto 0);
  signal transition_1057_symbol_out : boolean;
  signal transition_1057_preds : BooleanArray(0 downto 0);
  signal transition_1058_symbol_out : boolean;
  signal transition_1058_preds : BooleanArray(0 downto 0);
  signal transition_1059_symbol_out : boolean;
  signal transition_1059_preds : BooleanArray(0 downto 0);
  signal transition_1063_symbol_out : boolean;
  signal transition_1063_preds : BooleanArray(0 downto 0);
  signal transition_1064_symbol_out : boolean;
  signal transition_1064_preds : BooleanArray(0 downto 0);
  signal transition_1065_symbol_out : boolean;
  signal transition_1065_preds : BooleanArray(0 downto 0);
  signal transition_1066_symbol_out : boolean;
  signal transition_1066_preds : BooleanArray(0 downto 0);
  signal transition_1070_symbol_out : boolean;
  signal transition_1070_preds : BooleanArray(1 downto 0);
  signal transition_1071_symbol_out : boolean;
  signal transition_1071_preds : BooleanArray(0 downto 0);
  signal transition_1072_symbol_out : boolean;
  signal transition_1072_preds : BooleanArray(0 downto 0);
  signal transition_1073_symbol_out : boolean;
  signal transition_1073_preds : BooleanArray(0 downto 0);
  signal transition_1074_symbol_out : boolean;
  signal transition_1074_preds : BooleanArray(0 downto 0);
  signal transition_1078_symbol_out : boolean;
  signal transition_1078_preds : BooleanArray(1 downto 0);
  signal transition_1080_symbol_out : boolean;
  signal transition_1080_preds : BooleanArray(0 downto 0);
  signal transition_1081_symbol_out : boolean;
  signal transition_1081_preds : BooleanArray(0 downto 0);

begin
  place_0_preds(0) <= transition_2_symbol_out;
  place_0_succs(0) <= transition_1_symbol_out;
  place_0 : place
    generic map(marking => true)
    port map(
      preds => place_0_preds,
      succs => place_0_succs,
      token => place_0_token,
      clk   => clk,
      reset => reset);

  place_6_preds(0) <= transition_9_symbol_out;
  place_6_succs(0) <= transition_7_symbol_out;
  place_6_succs(1) <= transition_8_symbol_out;
  place_6 : place
    generic map(marking => false)
    port map(
      preds => place_6_preds,
      succs => place_6_succs,
      token => place_6_token,
      clk   => clk,
      reset => reset);

  place_13_preds(0) <= transition_16_symbol_out;
  place_13_succs(0) <= transition_14_symbol_out;
  place_13_succs(1) <= transition_15_symbol_out;
  place_13 : place
    generic map(marking => false)
    port map(
      preds => place_13_preds,
      succs => place_13_succs,
      token => place_13_token,
      clk   => clk,
      reset => reset);

  place_18_preds(0) <= transition_20_symbol_out;
  place_18_succs(0) <= transition_19_symbol_out;
  place_18 : place
    generic map(marking => false)
    port map(
      preds => place_18_preds,
      succs => place_18_succs,
      token => place_18_token,
      clk   => clk,
      reset => reset);

  place_24_preds(0) <= transition_26_symbol_out;
  place_24_preds(1) <= transition_27_symbol_out;
  place_24_succs(0) <= transition_25_symbol_out;
  place_24 : place
    generic map(marking => false)
    port map(
      preds => place_24_preds,
      succs => place_24_succs,
      token => place_24_token,
      clk   => clk,
      reset => reset);

  place_28_preds(0) <= transition_30_symbol_out;
  place_28_preds(1) <= transition_31_symbol_out;
  place_28_succs(0) <= transition_29_symbol_out;
  place_28 : place
    generic map(marking => false)
    port map(
      preds => place_28_preds,
      succs => place_28_succs,
      token => place_28_token,
      clk   => clk,
      reset => reset);

  place_36_preds(0) <= transition_32_symbol_out;
  place_36_succs(0) <= transition_33_symbol_out;
  place_36 : place
    generic map(marking => false)
    port map(
      preds => place_36_preds,
      succs => place_36_succs,
      token => place_36_token,
      clk   => clk,
      reset => reset);

  place_37_preds(0) <= transition_33_symbol_out;
  place_37_succs(0) <= transition_34_symbol_out;
  place_37 : place
    generic map(marking => false)
    port map(
      preds => place_37_preds,
      succs => place_37_succs,
      token => place_37_token,
      clk   => clk,
      reset => reset);

  place_38_preds(0) <= transition_34_symbol_out;
  place_38_succs(0) <= transition_35_symbol_out;
  place_38 : place
    generic map(marking => false)
    port map(
      preds => place_38_preds,
      succs => place_38_succs,
      token => place_38_token,
      clk   => clk,
      reset => reset);

  place_43_preds(0) <= transition_39_symbol_out;
  place_43_succs(0) <= transition_40_symbol_out;
  place_43 : place
    generic map(marking => false)
    port map(
      preds => place_43_preds,
      succs => place_43_succs,
      token => place_43_token,
      clk   => clk,
      reset => reset);

  place_44_preds(0) <= transition_40_symbol_out;
  place_44_succs(0) <= transition_41_symbol_out;
  place_44 : place
    generic map(marking => false)
    port map(
      preds => place_44_preds,
      succs => place_44_succs,
      token => place_44_token,
      clk   => clk,
      reset => reset);

  place_45_preds(0) <= transition_41_symbol_out;
  place_45_succs(0) <= transition_42_symbol_out;
  place_45 : place
    generic map(marking => false)
    port map(
      preds => place_45_preds,
      succs => place_45_succs,
      token => place_45_token,
      clk   => clk,
      reset => reset);

  place_50_preds(0) <= transition_46_symbol_out;
  place_50_succs(0) <= transition_47_symbol_out;
  place_50 : place
    generic map(marking => false)
    port map(
      preds => place_50_preds,
      succs => place_50_succs,
      token => place_50_token,
      clk   => clk,
      reset => reset);

  place_51_preds(0) <= transition_47_symbol_out;
  place_51_succs(0) <= transition_48_symbol_out;
  place_51 : place
    generic map(marking => false)
    port map(
      preds => place_51_preds,
      succs => place_51_succs,
      token => place_51_token,
      clk   => clk,
      reset => reset);

  place_52_preds(0) <= transition_48_symbol_out;
  place_52_succs(0) <= transition_49_symbol_out;
  place_52 : place
    generic map(marking => false)
    port map(
      preds => place_52_preds,
      succs => place_52_succs,
      token => place_52_token,
      clk   => clk,
      reset => reset);

  place_58_preds(0) <= transition_54_symbol_out;
  place_58_succs(0) <= transition_55_symbol_out;
  place_58 : place
    generic map(marking => false)
    port map(
      preds => place_58_preds,
      succs => place_58_succs,
      token => place_58_token,
      clk   => clk,
      reset => reset);

  place_59_preds(0) <= transition_55_symbol_out;
  place_59_succs(0) <= transition_56_symbol_out;
  place_59 : place
    generic map(marking => false)
    port map(
      preds => place_59_preds,
      succs => place_59_succs,
      token => place_59_token,
      clk   => clk,
      reset => reset);

  place_60_preds(0) <= transition_56_symbol_out;
  place_60_succs(0) <= transition_57_symbol_out;
  place_60 : place
    generic map(marking => false)
    port map(
      preds => place_60_preds,
      succs => place_60_succs,
      token => place_60_token,
      clk   => clk,
      reset => reset);

  place_65_preds(0) <= transition_61_symbol_out;
  place_65_succs(0) <= transition_62_symbol_out;
  place_65 : place
    generic map(marking => false)
    port map(
      preds => place_65_preds,
      succs => place_65_succs,
      token => place_65_token,
      clk   => clk,
      reset => reset);

  place_66_preds(0) <= transition_62_symbol_out;
  place_66_succs(0) <= transition_63_symbol_out;
  place_66 : place
    generic map(marking => false)
    port map(
      preds => place_66_preds,
      succs => place_66_succs,
      token => place_66_token,
      clk   => clk,
      reset => reset);

  place_67_preds(0) <= transition_63_symbol_out;
  place_67_succs(0) <= transition_64_symbol_out;
  place_67 : place
    generic map(marking => false)
    port map(
      preds => place_67_preds,
      succs => place_67_succs,
      token => place_67_token,
      clk   => clk,
      reset => reset);

  place_73_preds(0) <= transition_69_symbol_out;
  place_73_succs(0) <= transition_70_symbol_out;
  place_73 : place
    generic map(marking => false)
    port map(
      preds => place_73_preds,
      succs => place_73_succs,
      token => place_73_token,
      clk   => clk,
      reset => reset);

  place_74_preds(0) <= transition_70_symbol_out;
  place_74_succs(0) <= transition_71_symbol_out;
  place_74 : place
    generic map(marking => false)
    port map(
      preds => place_74_preds,
      succs => place_74_succs,
      token => place_74_token,
      clk   => clk,
      reset => reset);

  place_75_preds(0) <= transition_71_symbol_out;
  place_75_succs(0) <= transition_72_symbol_out;
  place_75 : place
    generic map(marking => false)
    port map(
      preds => place_75_preds,
      succs => place_75_succs,
      token => place_75_token,
      clk   => clk,
      reset => reset);

  place_80_preds(0) <= transition_76_symbol_out;
  place_80_succs(0) <= transition_77_symbol_out;
  place_80 : place
    generic map(marking => false)
    port map(
      preds => place_80_preds,
      succs => place_80_succs,
      token => place_80_token,
      clk   => clk,
      reset => reset);

  place_81_preds(0) <= transition_77_symbol_out;
  place_81_succs(0) <= transition_78_symbol_out;
  place_81 : place
    generic map(marking => false)
    port map(
      preds => place_81_preds,
      succs => place_81_succs,
      token => place_81_token,
      clk   => clk,
      reset => reset);

  place_82_preds(0) <= transition_78_symbol_out;
  place_82_succs(0) <= transition_79_symbol_out;
  place_82 : place
    generic map(marking => false)
    port map(
      preds => place_82_preds,
      succs => place_82_succs,
      token => place_82_token,
      clk   => clk,
      reset => reset);

  place_87_preds(0) <= transition_83_symbol_out;
  place_87_succs(0) <= transition_84_symbol_out;
  place_87 : place
    generic map(marking => false)
    port map(
      preds => place_87_preds,
      succs => place_87_succs,
      token => place_87_token,
      clk   => clk,
      reset => reset);

  place_88_preds(0) <= transition_84_symbol_out;
  place_88_succs(0) <= transition_85_symbol_out;
  place_88 : place
    generic map(marking => false)
    port map(
      preds => place_88_preds,
      succs => place_88_succs,
      token => place_88_token,
      clk   => clk,
      reset => reset);

  place_89_preds(0) <= transition_85_symbol_out;
  place_89_succs(0) <= transition_86_symbol_out;
  place_89 : place
    generic map(marking => false)
    port map(
      preds => place_89_preds,
      succs => place_89_succs,
      token => place_89_token,
      clk   => clk,
      reset => reset);

  place_94_preds(0) <= transition_90_symbol_out;
  place_94_succs(0) <= transition_91_symbol_out;
  place_94 : place
    generic map(marking => false)
    port map(
      preds => place_94_preds,
      succs => place_94_succs,
      token => place_94_token,
      clk   => clk,
      reset => reset);

  place_95_preds(0) <= transition_91_symbol_out;
  place_95_succs(0) <= transition_92_symbol_out;
  place_95 : place
    generic map(marking => false)
    port map(
      preds => place_95_preds,
      succs => place_95_succs,
      token => place_95_token,
      clk   => clk,
      reset => reset);

  place_96_preds(0) <= transition_92_symbol_out;
  place_96_succs(0) <= transition_93_symbol_out;
  place_96 : place
    generic map(marking => false)
    port map(
      preds => place_96_preds,
      succs => place_96_succs,
      token => place_96_token,
      clk   => clk,
      reset => reset);

  place_102_preds(0) <= transition_98_symbol_out;
  place_102_succs(0) <= transition_99_symbol_out;
  place_102 : place
    generic map(marking => false)
    port map(
      preds => place_102_preds,
      succs => place_102_succs,
      token => place_102_token,
      clk   => clk,
      reset => reset);

  place_103_preds(0) <= transition_99_symbol_out;
  place_103_succs(0) <= transition_100_symbol_out;
  place_103 : place
    generic map(marking => false)
    port map(
      preds => place_103_preds,
      succs => place_103_succs,
      token => place_103_token,
      clk   => clk,
      reset => reset);

  place_104_preds(0) <= transition_100_symbol_out;
  place_104_succs(0) <= transition_101_symbol_out;
  place_104 : place
    generic map(marking => false)
    port map(
      preds => place_104_preds,
      succs => place_104_succs,
      token => place_104_token,
      clk   => clk,
      reset => reset);

  place_109_preds(0) <= transition_105_symbol_out;
  place_109_succs(0) <= transition_106_symbol_out;
  place_109 : place
    generic map(marking => false)
    port map(
      preds => place_109_preds,
      succs => place_109_succs,
      token => place_109_token,
      clk   => clk,
      reset => reset);

  place_110_preds(0) <= transition_106_symbol_out;
  place_110_succs(0) <= transition_107_symbol_out;
  place_110 : place
    generic map(marking => false)
    port map(
      preds => place_110_preds,
      succs => place_110_succs,
      token => place_110_token,
      clk   => clk,
      reset => reset);

  place_111_preds(0) <= transition_107_symbol_out;
  place_111_succs(0) <= transition_108_symbol_out;
  place_111 : place
    generic map(marking => false)
    port map(
      preds => place_111_preds,
      succs => place_111_succs,
      token => place_111_token,
      clk   => clk,
      reset => reset);

  place_117_preds(0) <= transition_113_symbol_out;
  place_117_succs(0) <= transition_114_symbol_out;
  place_117 : place
    generic map(marking => false)
    port map(
      preds => place_117_preds,
      succs => place_117_succs,
      token => place_117_token,
      clk   => clk,
      reset => reset);

  place_118_preds(0) <= transition_114_symbol_out;
  place_118_succs(0) <= transition_115_symbol_out;
  place_118 : place
    generic map(marking => false)
    port map(
      preds => place_118_preds,
      succs => place_118_succs,
      token => place_118_token,
      clk   => clk,
      reset => reset);

  place_119_preds(0) <= transition_115_symbol_out;
  place_119_succs(0) <= transition_116_symbol_out;
  place_119 : place
    generic map(marking => false)
    port map(
      preds => place_119_preds,
      succs => place_119_succs,
      token => place_119_token,
      clk   => clk,
      reset => reset);

  place_124_preds(0) <= transition_120_symbol_out;
  place_124_succs(0) <= transition_121_symbol_out;
  place_124 : place
    generic map(marking => false)
    port map(
      preds => place_124_preds,
      succs => place_124_succs,
      token => place_124_token,
      clk   => clk,
      reset => reset);

  place_125_preds(0) <= transition_121_symbol_out;
  place_125_succs(0) <= transition_122_symbol_out;
  place_125 : place
    generic map(marking => false)
    port map(
      preds => place_125_preds,
      succs => place_125_succs,
      token => place_125_token,
      clk   => clk,
      reset => reset);

  place_126_preds(0) <= transition_122_symbol_out;
  place_126_succs(0) <= transition_123_symbol_out;
  place_126 : place
    generic map(marking => false)
    port map(
      preds => place_126_preds,
      succs => place_126_succs,
      token => place_126_token,
      clk   => clk,
      reset => reset);

  place_131_preds(0) <= transition_127_symbol_out;
  place_131_succs(0) <= transition_128_symbol_out;
  place_131 : place
    generic map(marking => false)
    port map(
      preds => place_131_preds,
      succs => place_131_succs,
      token => place_131_token,
      clk   => clk,
      reset => reset);

  place_132_preds(0) <= transition_128_symbol_out;
  place_132_succs(0) <= transition_129_symbol_out;
  place_132 : place
    generic map(marking => false)
    port map(
      preds => place_132_preds,
      succs => place_132_succs,
      token => place_132_token,
      clk   => clk,
      reset => reset);

  place_133_preds(0) <= transition_129_symbol_out;
  place_133_succs(0) <= transition_130_symbol_out;
  place_133 : place
    generic map(marking => false)
    port map(
      preds => place_133_preds,
      succs => place_133_succs,
      token => place_133_token,
      clk   => clk,
      reset => reset);

  place_138_preds(0) <= transition_134_symbol_out;
  place_138_succs(0) <= transition_135_symbol_out;
  place_138 : place
    generic map(marking => false)
    port map(
      preds => place_138_preds,
      succs => place_138_succs,
      token => place_138_token,
      clk   => clk,
      reset => reset);

  place_139_preds(0) <= transition_135_symbol_out;
  place_139_succs(0) <= transition_136_symbol_out;
  place_139 : place
    generic map(marking => false)
    port map(
      preds => place_139_preds,
      succs => place_139_succs,
      token => place_139_token,
      clk   => clk,
      reset => reset);

  place_140_preds(0) <= transition_136_symbol_out;
  place_140_succs(0) <= transition_137_symbol_out;
  place_140 : place
    generic map(marking => false)
    port map(
      preds => place_140_preds,
      succs => place_140_succs,
      token => place_140_token,
      clk   => clk,
      reset => reset);

  place_146_preds(0) <= transition_142_symbol_out;
  place_146_succs(0) <= transition_143_symbol_out;
  place_146 : place
    generic map(marking => false)
    port map(
      preds => place_146_preds,
      succs => place_146_succs,
      token => place_146_token,
      clk   => clk,
      reset => reset);

  place_147_preds(0) <= transition_143_symbol_out;
  place_147_succs(0) <= transition_144_symbol_out;
  place_147 : place
    generic map(marking => false)
    port map(
      preds => place_147_preds,
      succs => place_147_succs,
      token => place_147_token,
      clk   => clk,
      reset => reset);

  place_148_preds(0) <= transition_144_symbol_out;
  place_148_succs(0) <= transition_145_symbol_out;
  place_148 : place
    generic map(marking => false)
    port map(
      preds => place_148_preds,
      succs => place_148_succs,
      token => place_148_token,
      clk   => clk,
      reset => reset);

  place_153_preds(0) <= transition_149_symbol_out;
  place_153_succs(0) <= transition_150_symbol_out;
  place_153 : place
    generic map(marking => false)
    port map(
      preds => place_153_preds,
      succs => place_153_succs,
      token => place_153_token,
      clk   => clk,
      reset => reset);

  place_154_preds(0) <= transition_150_symbol_out;
  place_154_succs(0) <= transition_151_symbol_out;
  place_154 : place
    generic map(marking => false)
    port map(
      preds => place_154_preds,
      succs => place_154_succs,
      token => place_154_token,
      clk   => clk,
      reset => reset);

  place_155_preds(0) <= transition_151_symbol_out;
  place_155_succs(0) <= transition_152_symbol_out;
  place_155 : place
    generic map(marking => false)
    port map(
      preds => place_155_preds,
      succs => place_155_succs,
      token => place_155_token,
      clk   => clk,
      reset => reset);

  place_160_preds(0) <= transition_156_symbol_out;
  place_160_succs(0) <= transition_157_symbol_out;
  place_160 : place
    generic map(marking => false)
    port map(
      preds => place_160_preds,
      succs => place_160_succs,
      token => place_160_token,
      clk   => clk,
      reset => reset);

  place_161_preds(0) <= transition_157_symbol_out;
  place_161_succs(0) <= transition_158_symbol_out;
  place_161 : place
    generic map(marking => false)
    port map(
      preds => place_161_preds,
      succs => place_161_succs,
      token => place_161_token,
      clk   => clk,
      reset => reset);

  place_162_preds(0) <= transition_158_symbol_out;
  place_162_succs(0) <= transition_159_symbol_out;
  place_162 : place
    generic map(marking => false)
    port map(
      preds => place_162_preds,
      succs => place_162_succs,
      token => place_162_token,
      clk   => clk,
      reset => reset);

  place_165_preds(0) <= transition_167_symbol_out;
  place_165_succs(0) <= transition_166_symbol_out;
  place_165 : place
    generic map(marking => false)
    port map(
      preds => place_165_preds,
      succs => place_165_succs,
      token => place_165_token,
      clk   => clk,
      reset => reset);

  place_173_preds(0) <= transition_169_symbol_out;
  place_173_succs(0) <= transition_170_symbol_out;
  place_173 : place
    generic map(marking => false)
    port map(
      preds => place_173_preds,
      succs => place_173_succs,
      token => place_173_token,
      clk   => clk,
      reset => reset);

  place_174_preds(0) <= transition_170_symbol_out;
  place_174_succs(0) <= transition_171_symbol_out;
  place_174 : place
    generic map(marking => false)
    port map(
      preds => place_174_preds,
      succs => place_174_succs,
      token => place_174_token,
      clk   => clk,
      reset => reset);

  place_175_preds(0) <= transition_171_symbol_out;
  place_175_succs(0) <= transition_172_symbol_out;
  place_175 : place
    generic map(marking => false)
    port map(
      preds => place_175_preds,
      succs => place_175_succs,
      token => place_175_token,
      clk   => clk,
      reset => reset);

  place_180_preds(0) <= transition_176_symbol_out;
  place_180_succs(0) <= transition_177_symbol_out;
  place_180 : place
    generic map(marking => false)
    port map(
      preds => place_180_preds,
      succs => place_180_succs,
      token => place_180_token,
      clk   => clk,
      reset => reset);

  place_181_preds(0) <= transition_177_symbol_out;
  place_181_succs(0) <= transition_178_symbol_out;
  place_181 : place
    generic map(marking => false)
    port map(
      preds => place_181_preds,
      succs => place_181_succs,
      token => place_181_token,
      clk   => clk,
      reset => reset);

  place_182_preds(0) <= transition_178_symbol_out;
  place_182_succs(0) <= transition_179_symbol_out;
  place_182 : place
    generic map(marking => false)
    port map(
      preds => place_182_preds,
      succs => place_182_succs,
      token => place_182_token,
      clk   => clk,
      reset => reset);

  place_187_preds(0) <= transition_183_symbol_out;
  place_187_succs(0) <= transition_184_symbol_out;
  place_187 : place
    generic map(marking => false)
    port map(
      preds => place_187_preds,
      succs => place_187_succs,
      token => place_187_token,
      clk   => clk,
      reset => reset);

  place_188_preds(0) <= transition_184_symbol_out;
  place_188_succs(0) <= transition_185_symbol_out;
  place_188 : place
    generic map(marking => false)
    port map(
      preds => place_188_preds,
      succs => place_188_succs,
      token => place_188_token,
      clk   => clk,
      reset => reset);

  place_189_preds(0) <= transition_185_symbol_out;
  place_189_succs(0) <= transition_186_symbol_out;
  place_189 : place
    generic map(marking => false)
    port map(
      preds => place_189_preds,
      succs => place_189_succs,
      token => place_189_token,
      clk   => clk,
      reset => reset);

  place_195_preds(0) <= transition_191_symbol_out;
  place_195_succs(0) <= transition_192_symbol_out;
  place_195 : place
    generic map(marking => false)
    port map(
      preds => place_195_preds,
      succs => place_195_succs,
      token => place_195_token,
      clk   => clk,
      reset => reset);

  place_196_preds(0) <= transition_192_symbol_out;
  place_196_succs(0) <= transition_193_symbol_out;
  place_196 : place
    generic map(marking => false)
    port map(
      preds => place_196_preds,
      succs => place_196_succs,
      token => place_196_token,
      clk   => clk,
      reset => reset);

  place_197_preds(0) <= transition_193_symbol_out;
  place_197_succs(0) <= transition_194_symbol_out;
  place_197 : place
    generic map(marking => false)
    port map(
      preds => place_197_preds,
      succs => place_197_succs,
      token => place_197_token,
      clk   => clk,
      reset => reset);

  place_202_preds(0) <= transition_198_symbol_out;
  place_202_succs(0) <= transition_199_symbol_out;
  place_202 : place
    generic map(marking => false)
    port map(
      preds => place_202_preds,
      succs => place_202_succs,
      token => place_202_token,
      clk   => clk,
      reset => reset);

  place_203_preds(0) <= transition_199_symbol_out;
  place_203_succs(0) <= transition_200_symbol_out;
  place_203 : place
    generic map(marking => false)
    port map(
      preds => place_203_preds,
      succs => place_203_succs,
      token => place_203_token,
      clk   => clk,
      reset => reset);

  place_204_preds(0) <= transition_200_symbol_out;
  place_204_succs(0) <= transition_201_symbol_out;
  place_204 : place
    generic map(marking => false)
    port map(
      preds => place_204_preds,
      succs => place_204_succs,
      token => place_204_token,
      clk   => clk,
      reset => reset);

  place_209_preds(0) <= transition_205_symbol_out;
  place_209_succs(0) <= transition_206_symbol_out;
  place_209 : place
    generic map(marking => false)
    port map(
      preds => place_209_preds,
      succs => place_209_succs,
      token => place_209_token,
      clk   => clk,
      reset => reset);

  place_210_preds(0) <= transition_206_symbol_out;
  place_210_succs(0) <= transition_207_symbol_out;
  place_210 : place
    generic map(marking => false)
    port map(
      preds => place_210_preds,
      succs => place_210_succs,
      token => place_210_token,
      clk   => clk,
      reset => reset);

  place_211_preds(0) <= transition_207_symbol_out;
  place_211_succs(0) <= transition_208_symbol_out;
  place_211 : place
    generic map(marking => false)
    port map(
      preds => place_211_preds,
      succs => place_211_succs,
      token => place_211_token,
      clk   => clk,
      reset => reset);

  place_213_preds(0) <= transition_215_symbol_out;
  place_213_succs(0) <= transition_214_symbol_out;
  place_213 : place
    generic map(marking => false)
    port map(
      preds => place_213_preds,
      succs => place_213_succs,
      token => place_213_token,
      clk   => clk,
      reset => reset);

  place_221_preds(0) <= transition_217_symbol_out;
  place_221_succs(0) <= transition_218_symbol_out;
  place_221 : place
    generic map(marking => false)
    port map(
      preds => place_221_preds,
      succs => place_221_succs,
      token => place_221_token,
      clk   => clk,
      reset => reset);

  place_222_preds(0) <= transition_218_symbol_out;
  place_222_succs(0) <= transition_219_symbol_out;
  place_222 : place
    generic map(marking => false)
    port map(
      preds => place_222_preds,
      succs => place_222_succs,
      token => place_222_token,
      clk   => clk,
      reset => reset);

  place_223_preds(0) <= transition_219_symbol_out;
  place_223_succs(0) <= transition_220_symbol_out;
  place_223 : place
    generic map(marking => false)
    port map(
      preds => place_223_preds,
      succs => place_223_succs,
      token => place_223_token,
      clk   => clk,
      reset => reset);

  place_228_preds(0) <= transition_224_symbol_out;
  place_228_succs(0) <= transition_225_symbol_out;
  place_228 : place
    generic map(marking => false)
    port map(
      preds => place_228_preds,
      succs => place_228_succs,
      token => place_228_token,
      clk   => clk,
      reset => reset);

  place_229_preds(0) <= transition_225_symbol_out;
  place_229_succs(0) <= transition_226_symbol_out;
  place_229 : place
    generic map(marking => false)
    port map(
      preds => place_229_preds,
      succs => place_229_succs,
      token => place_229_token,
      clk   => clk,
      reset => reset);

  place_230_preds(0) <= transition_226_symbol_out;
  place_230_succs(0) <= transition_227_symbol_out;
  place_230 : place
    generic map(marking => false)
    port map(
      preds => place_230_preds,
      succs => place_230_succs,
      token => place_230_token,
      clk   => clk,
      reset => reset);

  place_232_preds(0) <= transition_234_symbol_out;
  place_232_preds(1) <= transition_235_symbol_out;
  place_232_succs(0) <= transition_233_symbol_out;
  place_232 : place
    generic map(marking => false)
    port map(
      preds => place_232_preds,
      succs => place_232_succs,
      token => place_232_token,
      clk   => clk,
      reset => reset);

  place_236_preds(0) <= transition_238_symbol_out;
  place_236_preds(1) <= transition_239_symbol_out;
  place_236_succs(0) <= transition_237_symbol_out;
  place_236 : place
    generic map(marking => false)
    port map(
      preds => place_236_preds,
      succs => place_236_succs,
      token => place_236_token,
      clk   => clk,
      reset => reset);

  place_244_preds(0) <= transition_240_symbol_out;
  place_244_succs(0) <= transition_241_symbol_out;
  place_244 : place
    generic map(marking => false)
    port map(
      preds => place_244_preds,
      succs => place_244_succs,
      token => place_244_token,
      clk   => clk,
      reset => reset);

  place_245_preds(0) <= transition_241_symbol_out;
  place_245_succs(0) <= transition_242_symbol_out;
  place_245 : place
    generic map(marking => false)
    port map(
      preds => place_245_preds,
      succs => place_245_succs,
      token => place_245_token,
      clk   => clk,
      reset => reset);

  place_246_preds(0) <= transition_242_symbol_out;
  place_246_succs(0) <= transition_243_symbol_out;
  place_246 : place
    generic map(marking => false)
    port map(
      preds => place_246_preds,
      succs => place_246_succs,
      token => place_246_token,
      clk   => clk,
      reset => reset);

  place_251_preds(0) <= transition_247_symbol_out;
  place_251_succs(0) <= transition_248_symbol_out;
  place_251 : place
    generic map(marking => false)
    port map(
      preds => place_251_preds,
      succs => place_251_succs,
      token => place_251_token,
      clk   => clk,
      reset => reset);

  place_252_preds(0) <= transition_248_symbol_out;
  place_252_succs(0) <= transition_249_symbol_out;
  place_252 : place
    generic map(marking => false)
    port map(
      preds => place_252_preds,
      succs => place_252_succs,
      token => place_252_token,
      clk   => clk,
      reset => reset);

  place_253_preds(0) <= transition_249_symbol_out;
  place_253_succs(0) <= transition_250_symbol_out;
  place_253 : place
    generic map(marking => false)
    port map(
      preds => place_253_preds,
      succs => place_253_succs,
      token => place_253_token,
      clk   => clk,
      reset => reset);

  place_258_preds(0) <= transition_254_symbol_out;
  place_258_succs(0) <= transition_255_symbol_out;
  place_258 : place
    generic map(marking => false)
    port map(
      preds => place_258_preds,
      succs => place_258_succs,
      token => place_258_token,
      clk   => clk,
      reset => reset);

  place_259_preds(0) <= transition_255_symbol_out;
  place_259_succs(0) <= transition_256_symbol_out;
  place_259 : place
    generic map(marking => false)
    port map(
      preds => place_259_preds,
      succs => place_259_succs,
      token => place_259_token,
      clk   => clk,
      reset => reset);

  place_260_preds(0) <= transition_256_symbol_out;
  place_260_succs(0) <= transition_257_symbol_out;
  place_260 : place
    generic map(marking => false)
    port map(
      preds => place_260_preds,
      succs => place_260_succs,
      token => place_260_token,
      clk   => clk,
      reset => reset);

  place_266_preds(0) <= transition_262_symbol_out;
  place_266_succs(0) <= transition_263_symbol_out;
  place_266 : place
    generic map(marking => false)
    port map(
      preds => place_266_preds,
      succs => place_266_succs,
      token => place_266_token,
      clk   => clk,
      reset => reset);

  place_267_preds(0) <= transition_263_symbol_out;
  place_267_succs(0) <= transition_264_symbol_out;
  place_267 : place
    generic map(marking => false)
    port map(
      preds => place_267_preds,
      succs => place_267_succs,
      token => place_267_token,
      clk   => clk,
      reset => reset);

  place_268_preds(0) <= transition_264_symbol_out;
  place_268_succs(0) <= transition_265_symbol_out;
  place_268 : place
    generic map(marking => false)
    port map(
      preds => place_268_preds,
      succs => place_268_succs,
      token => place_268_token,
      clk   => clk,
      reset => reset);

  place_273_preds(0) <= transition_269_symbol_out;
  place_273_succs(0) <= transition_270_symbol_out;
  place_273 : place
    generic map(marking => false)
    port map(
      preds => place_273_preds,
      succs => place_273_succs,
      token => place_273_token,
      clk   => clk,
      reset => reset);

  place_274_preds(0) <= transition_270_symbol_out;
  place_274_succs(0) <= transition_271_symbol_out;
  place_274 : place
    generic map(marking => false)
    port map(
      preds => place_274_preds,
      succs => place_274_succs,
      token => place_274_token,
      clk   => clk,
      reset => reset);

  place_275_preds(0) <= transition_271_symbol_out;
  place_275_succs(0) <= transition_272_symbol_out;
  place_275 : place
    generic map(marking => false)
    port map(
      preds => place_275_preds,
      succs => place_275_succs,
      token => place_275_token,
      clk   => clk,
      reset => reset);

  place_281_preds(0) <= transition_277_symbol_out;
  place_281_succs(0) <= transition_278_symbol_out;
  place_281 : place
    generic map(marking => false)
    port map(
      preds => place_281_preds,
      succs => place_281_succs,
      token => place_281_token,
      clk   => clk,
      reset => reset);

  place_282_preds(0) <= transition_278_symbol_out;
  place_282_succs(0) <= transition_279_symbol_out;
  place_282 : place
    generic map(marking => false)
    port map(
      preds => place_282_preds,
      succs => place_282_succs,
      token => place_282_token,
      clk   => clk,
      reset => reset);

  place_283_preds(0) <= transition_279_symbol_out;
  place_283_succs(0) <= transition_280_symbol_out;
  place_283 : place
    generic map(marking => false)
    port map(
      preds => place_283_preds,
      succs => place_283_succs,
      token => place_283_token,
      clk   => clk,
      reset => reset);

  place_288_preds(0) <= transition_284_symbol_out;
  place_288_succs(0) <= transition_285_symbol_out;
  place_288 : place
    generic map(marking => false)
    port map(
      preds => place_288_preds,
      succs => place_288_succs,
      token => place_288_token,
      clk   => clk,
      reset => reset);

  place_289_preds(0) <= transition_285_symbol_out;
  place_289_succs(0) <= transition_286_symbol_out;
  place_289 : place
    generic map(marking => false)
    port map(
      preds => place_289_preds,
      succs => place_289_succs,
      token => place_289_token,
      clk   => clk,
      reset => reset);

  place_290_preds(0) <= transition_286_symbol_out;
  place_290_succs(0) <= transition_287_symbol_out;
  place_290 : place
    generic map(marking => false)
    port map(
      preds => place_290_preds,
      succs => place_290_succs,
      token => place_290_token,
      clk   => clk,
      reset => reset);

  place_295_preds(0) <= transition_291_symbol_out;
  place_295_succs(0) <= transition_292_symbol_out;
  place_295 : place
    generic map(marking => false)
    port map(
      preds => place_295_preds,
      succs => place_295_succs,
      token => place_295_token,
      clk   => clk,
      reset => reset);

  place_296_preds(0) <= transition_292_symbol_out;
  place_296_succs(0) <= transition_293_symbol_out;
  place_296 : place
    generic map(marking => false)
    port map(
      preds => place_296_preds,
      succs => place_296_succs,
      token => place_296_token,
      clk   => clk,
      reset => reset);

  place_297_preds(0) <= transition_293_symbol_out;
  place_297_succs(0) <= transition_294_symbol_out;
  place_297 : place
    generic map(marking => false)
    port map(
      preds => place_297_preds,
      succs => place_297_succs,
      token => place_297_token,
      clk   => clk,
      reset => reset);

  place_302_preds(0) <= transition_298_symbol_out;
  place_302_succs(0) <= transition_299_symbol_out;
  place_302 : place
    generic map(marking => false)
    port map(
      preds => place_302_preds,
      succs => place_302_succs,
      token => place_302_token,
      clk   => clk,
      reset => reset);

  place_303_preds(0) <= transition_299_symbol_out;
  place_303_succs(0) <= transition_300_symbol_out;
  place_303 : place
    generic map(marking => false)
    port map(
      preds => place_303_preds,
      succs => place_303_succs,
      token => place_303_token,
      clk   => clk,
      reset => reset);

  place_304_preds(0) <= transition_300_symbol_out;
  place_304_succs(0) <= transition_301_symbol_out;
  place_304 : place
    generic map(marking => false)
    port map(
      preds => place_304_preds,
      succs => place_304_succs,
      token => place_304_token,
      clk   => clk,
      reset => reset);

  place_310_preds(0) <= transition_306_symbol_out;
  place_310_succs(0) <= transition_307_symbol_out;
  place_310 : place
    generic map(marking => false)
    port map(
      preds => place_310_preds,
      succs => place_310_succs,
      token => place_310_token,
      clk   => clk,
      reset => reset);

  place_311_preds(0) <= transition_307_symbol_out;
  place_311_succs(0) <= transition_308_symbol_out;
  place_311 : place
    generic map(marking => false)
    port map(
      preds => place_311_preds,
      succs => place_311_succs,
      token => place_311_token,
      clk   => clk,
      reset => reset);

  place_312_preds(0) <= transition_308_symbol_out;
  place_312_succs(0) <= transition_309_symbol_out;
  place_312 : place
    generic map(marking => false)
    port map(
      preds => place_312_preds,
      succs => place_312_succs,
      token => place_312_token,
      clk   => clk,
      reset => reset);

  place_317_preds(0) <= transition_313_symbol_out;
  place_317_succs(0) <= transition_314_symbol_out;
  place_317 : place
    generic map(marking => false)
    port map(
      preds => place_317_preds,
      succs => place_317_succs,
      token => place_317_token,
      clk   => clk,
      reset => reset);

  place_318_preds(0) <= transition_314_symbol_out;
  place_318_succs(0) <= transition_315_symbol_out;
  place_318 : place
    generic map(marking => false)
    port map(
      preds => place_318_preds,
      succs => place_318_succs,
      token => place_318_token,
      clk   => clk,
      reset => reset);

  place_319_preds(0) <= transition_315_symbol_out;
  place_319_succs(0) <= transition_316_symbol_out;
  place_319 : place
    generic map(marking => false)
    port map(
      preds => place_319_preds,
      succs => place_319_succs,
      token => place_319_token,
      clk   => clk,
      reset => reset);

  place_325_preds(0) <= transition_321_symbol_out;
  place_325_succs(0) <= transition_322_symbol_out;
  place_325 : place
    generic map(marking => false)
    port map(
      preds => place_325_preds,
      succs => place_325_succs,
      token => place_325_token,
      clk   => clk,
      reset => reset);

  place_326_preds(0) <= transition_322_symbol_out;
  place_326_succs(0) <= transition_323_symbol_out;
  place_326 : place
    generic map(marking => false)
    port map(
      preds => place_326_preds,
      succs => place_326_succs,
      token => place_326_token,
      clk   => clk,
      reset => reset);

  place_327_preds(0) <= transition_323_symbol_out;
  place_327_succs(0) <= transition_324_symbol_out;
  place_327 : place
    generic map(marking => false)
    port map(
      preds => place_327_preds,
      succs => place_327_succs,
      token => place_327_token,
      clk   => clk,
      reset => reset);

  place_332_preds(0) <= transition_328_symbol_out;
  place_332_succs(0) <= transition_329_symbol_out;
  place_332 : place
    generic map(marking => false)
    port map(
      preds => place_332_preds,
      succs => place_332_succs,
      token => place_332_token,
      clk   => clk,
      reset => reset);

  place_333_preds(0) <= transition_329_symbol_out;
  place_333_succs(0) <= transition_330_symbol_out;
  place_333 : place
    generic map(marking => false)
    port map(
      preds => place_333_preds,
      succs => place_333_succs,
      token => place_333_token,
      clk   => clk,
      reset => reset);

  place_334_preds(0) <= transition_330_symbol_out;
  place_334_succs(0) <= transition_331_symbol_out;
  place_334 : place
    generic map(marking => false)
    port map(
      preds => place_334_preds,
      succs => place_334_succs,
      token => place_334_token,
      clk   => clk,
      reset => reset);

  place_339_preds(0) <= transition_335_symbol_out;
  place_339_succs(0) <= transition_336_symbol_out;
  place_339 : place
    generic map(marking => false)
    port map(
      preds => place_339_preds,
      succs => place_339_succs,
      token => place_339_token,
      clk   => clk,
      reset => reset);

  place_340_preds(0) <= transition_336_symbol_out;
  place_340_succs(0) <= transition_337_symbol_out;
  place_340 : place
    generic map(marking => false)
    port map(
      preds => place_340_preds,
      succs => place_340_succs,
      token => place_340_token,
      clk   => clk,
      reset => reset);

  place_341_preds(0) <= transition_337_symbol_out;
  place_341_succs(0) <= transition_338_symbol_out;
  place_341 : place
    generic map(marking => false)
    port map(
      preds => place_341_preds,
      succs => place_341_succs,
      token => place_341_token,
      clk   => clk,
      reset => reset);

  place_346_preds(0) <= transition_342_symbol_out;
  place_346_succs(0) <= transition_343_symbol_out;
  place_346 : place
    generic map(marking => false)
    port map(
      preds => place_346_preds,
      succs => place_346_succs,
      token => place_346_token,
      clk   => clk,
      reset => reset);

  place_347_preds(0) <= transition_343_symbol_out;
  place_347_succs(0) <= transition_344_symbol_out;
  place_347 : place
    generic map(marking => false)
    port map(
      preds => place_347_preds,
      succs => place_347_succs,
      token => place_347_token,
      clk   => clk,
      reset => reset);

  place_348_preds(0) <= transition_344_symbol_out;
  place_348_succs(0) <= transition_345_symbol_out;
  place_348 : place
    generic map(marking => false)
    port map(
      preds => place_348_preds,
      succs => place_348_succs,
      token => place_348_token,
      clk   => clk,
      reset => reset);

  place_354_preds(0) <= transition_350_symbol_out;
  place_354_succs(0) <= transition_351_symbol_out;
  place_354 : place
    generic map(marking => false)
    port map(
      preds => place_354_preds,
      succs => place_354_succs,
      token => place_354_token,
      clk   => clk,
      reset => reset);

  place_355_preds(0) <= transition_351_symbol_out;
  place_355_succs(0) <= transition_352_symbol_out;
  place_355 : place
    generic map(marking => false)
    port map(
      preds => place_355_preds,
      succs => place_355_succs,
      token => place_355_token,
      clk   => clk,
      reset => reset);

  place_356_preds(0) <= transition_352_symbol_out;
  place_356_succs(0) <= transition_353_symbol_out;
  place_356 : place
    generic map(marking => false)
    port map(
      preds => place_356_preds,
      succs => place_356_succs,
      token => place_356_token,
      clk   => clk,
      reset => reset);

  place_361_preds(0) <= transition_357_symbol_out;
  place_361_succs(0) <= transition_358_symbol_out;
  place_361 : place
    generic map(marking => false)
    port map(
      preds => place_361_preds,
      succs => place_361_succs,
      token => place_361_token,
      clk   => clk,
      reset => reset);

  place_362_preds(0) <= transition_358_symbol_out;
  place_362_succs(0) <= transition_359_symbol_out;
  place_362 : place
    generic map(marking => false)
    port map(
      preds => place_362_preds,
      succs => place_362_succs,
      token => place_362_token,
      clk   => clk,
      reset => reset);

  place_363_preds(0) <= transition_359_symbol_out;
  place_363_succs(0) <= transition_360_symbol_out;
  place_363 : place
    generic map(marking => false)
    port map(
      preds => place_363_preds,
      succs => place_363_succs,
      token => place_363_token,
      clk   => clk,
      reset => reset);

  place_368_preds(0) <= transition_364_symbol_out;
  place_368_succs(0) <= transition_365_symbol_out;
  place_368 : place
    generic map(marking => false)
    port map(
      preds => place_368_preds,
      succs => place_368_succs,
      token => place_368_token,
      clk   => clk,
      reset => reset);

  place_369_preds(0) <= transition_365_symbol_out;
  place_369_succs(0) <= transition_366_symbol_out;
  place_369 : place
    generic map(marking => false)
    port map(
      preds => place_369_preds,
      succs => place_369_succs,
      token => place_369_token,
      clk   => clk,
      reset => reset);

  place_370_preds(0) <= transition_366_symbol_out;
  place_370_succs(0) <= transition_367_symbol_out;
  place_370 : place
    generic map(marking => false)
    port map(
      preds => place_370_preds,
      succs => place_370_succs,
      token => place_370_token,
      clk   => clk,
      reset => reset);

  place_377_preds(0) <= transition_373_symbol_out;
  place_377_succs(0) <= transition_374_symbol_out;
  place_377 : place
    generic map(marking => false)
    port map(
      preds => place_377_preds,
      succs => place_377_succs,
      token => place_377_token,
      clk   => clk,
      reset => reset);

  place_378_preds(0) <= transition_374_symbol_out;
  place_378_succs(0) <= transition_375_symbol_out;
  place_378 : place
    generic map(marking => false)
    port map(
      preds => place_378_preds,
      succs => place_378_succs,
      token => place_378_token,
      clk   => clk,
      reset => reset);

  place_379_preds(0) <= transition_375_symbol_out;
  place_379_succs(0) <= transition_376_symbol_out;
  place_379 : place
    generic map(marking => false)
    port map(
      preds => place_379_preds,
      succs => place_379_succs,
      token => place_379_token,
      clk   => clk,
      reset => reset);

  place_380_preds(0) <= transition_382_symbol_out;
  place_380_succs(0) <= transition_381_symbol_out;
  place_380 : place
    generic map(marking => false)
    port map(
      preds => place_380_preds,
      succs => place_380_succs,
      token => place_380_token,
      clk   => clk,
      reset => reset);

  place_388_preds(0) <= transition_384_symbol_out;
  place_388_succs(0) <= transition_385_symbol_out;
  place_388 : place
    generic map(marking => false)
    port map(
      preds => place_388_preds,
      succs => place_388_succs,
      token => place_388_token,
      clk   => clk,
      reset => reset);

  place_389_preds(0) <= transition_385_symbol_out;
  place_389_succs(0) <= transition_386_symbol_out;
  place_389 : place
    generic map(marking => false)
    port map(
      preds => place_389_preds,
      succs => place_389_succs,
      token => place_389_token,
      clk   => clk,
      reset => reset);

  place_390_preds(0) <= transition_386_symbol_out;
  place_390_succs(0) <= transition_387_symbol_out;
  place_390 : place
    generic map(marking => false)
    port map(
      preds => place_390_preds,
      succs => place_390_succs,
      token => place_390_token,
      clk   => clk,
      reset => reset);

  place_395_preds(0) <= transition_391_symbol_out;
  place_395_succs(0) <= transition_392_symbol_out;
  place_395 : place
    generic map(marking => false)
    port map(
      preds => place_395_preds,
      succs => place_395_succs,
      token => place_395_token,
      clk   => clk,
      reset => reset);

  place_396_preds(0) <= transition_392_symbol_out;
  place_396_succs(0) <= transition_393_symbol_out;
  place_396 : place
    generic map(marking => false)
    port map(
      preds => place_396_preds,
      succs => place_396_succs,
      token => place_396_token,
      clk   => clk,
      reset => reset);

  place_397_preds(0) <= transition_393_symbol_out;
  place_397_succs(0) <= transition_394_symbol_out;
  place_397 : place
    generic map(marking => false)
    port map(
      preds => place_397_preds,
      succs => place_397_succs,
      token => place_397_token,
      clk   => clk,
      reset => reset);

  place_402_preds(0) <= transition_398_symbol_out;
  place_402_succs(0) <= transition_399_symbol_out;
  place_402 : place
    generic map(marking => false)
    port map(
      preds => place_402_preds,
      succs => place_402_succs,
      token => place_402_token,
      clk   => clk,
      reset => reset);

  place_403_preds(0) <= transition_399_symbol_out;
  place_403_succs(0) <= transition_400_symbol_out;
  place_403 : place
    generic map(marking => false)
    port map(
      preds => place_403_preds,
      succs => place_403_succs,
      token => place_403_token,
      clk   => clk,
      reset => reset);

  place_404_preds(0) <= transition_400_symbol_out;
  place_404_succs(0) <= transition_401_symbol_out;
  place_404 : place
    generic map(marking => false)
    port map(
      preds => place_404_preds,
      succs => place_404_succs,
      token => place_404_token,
      clk   => clk,
      reset => reset);

  place_410_preds(0) <= transition_406_symbol_out;
  place_410_succs(0) <= transition_407_symbol_out;
  place_410 : place
    generic map(marking => false)
    port map(
      preds => place_410_preds,
      succs => place_410_succs,
      token => place_410_token,
      clk   => clk,
      reset => reset);

  place_411_preds(0) <= transition_407_symbol_out;
  place_411_succs(0) <= transition_408_symbol_out;
  place_411 : place
    generic map(marking => false)
    port map(
      preds => place_411_preds,
      succs => place_411_succs,
      token => place_411_token,
      clk   => clk,
      reset => reset);

  place_412_preds(0) <= transition_408_symbol_out;
  place_412_succs(0) <= transition_409_symbol_out;
  place_412 : place
    generic map(marking => false)
    port map(
      preds => place_412_preds,
      succs => place_412_succs,
      token => place_412_token,
      clk   => clk,
      reset => reset);

  place_417_preds(0) <= transition_413_symbol_out;
  place_417_succs(0) <= transition_414_symbol_out;
  place_417 : place
    generic map(marking => false)
    port map(
      preds => place_417_preds,
      succs => place_417_succs,
      token => place_417_token,
      clk   => clk,
      reset => reset);

  place_418_preds(0) <= transition_414_symbol_out;
  place_418_succs(0) <= transition_415_symbol_out;
  place_418 : place
    generic map(marking => false)
    port map(
      preds => place_418_preds,
      succs => place_418_succs,
      token => place_418_token,
      clk   => clk,
      reset => reset);

  place_419_preds(0) <= transition_415_symbol_out;
  place_419_succs(0) <= transition_416_symbol_out;
  place_419 : place
    generic map(marking => false)
    port map(
      preds => place_419_preds,
      succs => place_419_succs,
      token => place_419_token,
      clk   => clk,
      reset => reset);

  place_424_preds(0) <= transition_420_symbol_out;
  place_424_succs(0) <= transition_421_symbol_out;
  place_424 : place
    generic map(marking => false)
    port map(
      preds => place_424_preds,
      succs => place_424_succs,
      token => place_424_token,
      clk   => clk,
      reset => reset);

  place_425_preds(0) <= transition_421_symbol_out;
  place_425_succs(0) <= transition_422_symbol_out;
  place_425 : place
    generic map(marking => false)
    port map(
      preds => place_425_preds,
      succs => place_425_succs,
      token => place_425_token,
      clk   => clk,
      reset => reset);

  place_426_preds(0) <= transition_422_symbol_out;
  place_426_succs(0) <= transition_423_symbol_out;
  place_426 : place
    generic map(marking => false)
    port map(
      preds => place_426_preds,
      succs => place_426_succs,
      token => place_426_token,
      clk   => clk,
      reset => reset);

  place_432_preds(0) <= transition_428_symbol_out;
  place_432_succs(0) <= transition_429_symbol_out;
  place_432 : place
    generic map(marking => false)
    port map(
      preds => place_432_preds,
      succs => place_432_succs,
      token => place_432_token,
      clk   => clk,
      reset => reset);

  place_433_preds(0) <= transition_429_symbol_out;
  place_433_succs(0) <= transition_430_symbol_out;
  place_433 : place
    generic map(marking => false)
    port map(
      preds => place_433_preds,
      succs => place_433_succs,
      token => place_433_token,
      clk   => clk,
      reset => reset);

  place_434_preds(0) <= transition_430_symbol_out;
  place_434_succs(0) <= transition_431_symbol_out;
  place_434 : place
    generic map(marking => false)
    port map(
      preds => place_434_preds,
      succs => place_434_succs,
      token => place_434_token,
      clk   => clk,
      reset => reset);

  place_435_preds(0) <= transition_437_symbol_out;
  place_435_succs(0) <= transition_436_symbol_out;
  place_435 : place
    generic map(marking => false)
    port map(
      preds => place_435_preds,
      succs => place_435_succs,
      token => place_435_token,
      clk   => clk,
      reset => reset);

  place_443_preds(0) <= transition_439_symbol_out;
  place_443_succs(0) <= transition_440_symbol_out;
  place_443 : place
    generic map(marking => false)
    port map(
      preds => place_443_preds,
      succs => place_443_succs,
      token => place_443_token,
      clk   => clk,
      reset => reset);

  place_444_preds(0) <= transition_440_symbol_out;
  place_444_succs(0) <= transition_441_symbol_out;
  place_444 : place
    generic map(marking => false)
    port map(
      preds => place_444_preds,
      succs => place_444_succs,
      token => place_444_token,
      clk   => clk,
      reset => reset);

  place_445_preds(0) <= transition_441_symbol_out;
  place_445_succs(0) <= transition_442_symbol_out;
  place_445 : place
    generic map(marking => false)
    port map(
      preds => place_445_preds,
      succs => place_445_succs,
      token => place_445_token,
      clk   => clk,
      reset => reset);

  place_450_preds(0) <= transition_446_symbol_out;
  place_450_succs(0) <= transition_447_symbol_out;
  place_450 : place
    generic map(marking => false)
    port map(
      preds => place_450_preds,
      succs => place_450_succs,
      token => place_450_token,
      clk   => clk,
      reset => reset);

  place_451_preds(0) <= transition_447_symbol_out;
  place_451_succs(0) <= transition_448_symbol_out;
  place_451 : place
    generic map(marking => false)
    port map(
      preds => place_451_preds,
      succs => place_451_succs,
      token => place_451_token,
      clk   => clk,
      reset => reset);

  place_452_preds(0) <= transition_448_symbol_out;
  place_452_succs(0) <= transition_449_symbol_out;
  place_452 : place
    generic map(marking => false)
    port map(
      preds => place_452_preds,
      succs => place_452_succs,
      token => place_452_token,
      clk   => clk,
      reset => reset);

  place_457_preds(0) <= transition_453_symbol_out;
  place_457_succs(0) <= transition_454_symbol_out;
  place_457 : place
    generic map(marking => false)
    port map(
      preds => place_457_preds,
      succs => place_457_succs,
      token => place_457_token,
      clk   => clk,
      reset => reset);

  place_458_preds(0) <= transition_454_symbol_out;
  place_458_succs(0) <= transition_455_symbol_out;
  place_458 : place
    generic map(marking => false)
    port map(
      preds => place_458_preds,
      succs => place_458_succs,
      token => place_458_token,
      clk   => clk,
      reset => reset);

  place_459_preds(0) <= transition_455_symbol_out;
  place_459_succs(0) <= transition_456_symbol_out;
  place_459 : place
    generic map(marking => false)
    port map(
      preds => place_459_preds,
      succs => place_459_succs,
      token => place_459_token,
      clk   => clk,
      reset => reset);

  place_464_preds(0) <= transition_460_symbol_out;
  place_464_succs(0) <= transition_461_symbol_out;
  place_464 : place
    generic map(marking => false)
    port map(
      preds => place_464_preds,
      succs => place_464_succs,
      token => place_464_token,
      clk   => clk,
      reset => reset);

  place_465_preds(0) <= transition_461_symbol_out;
  place_465_succs(0) <= transition_462_symbol_out;
  place_465 : place
    generic map(marking => false)
    port map(
      preds => place_465_preds,
      succs => place_465_succs,
      token => place_465_token,
      clk   => clk,
      reset => reset);

  place_466_preds(0) <= transition_462_symbol_out;
  place_466_succs(0) <= transition_463_symbol_out;
  place_466 : place
    generic map(marking => false)
    port map(
      preds => place_466_preds,
      succs => place_466_succs,
      token => place_466_token,
      clk   => clk,
      reset => reset);

  place_471_preds(0) <= transition_467_symbol_out;
  place_471_succs(0) <= transition_468_symbol_out;
  place_471 : place
    generic map(marking => false)
    port map(
      preds => place_471_preds,
      succs => place_471_succs,
      token => place_471_token,
      clk   => clk,
      reset => reset);

  place_472_preds(0) <= transition_468_symbol_out;
  place_472_succs(0) <= transition_469_symbol_out;
  place_472 : place
    generic map(marking => false)
    port map(
      preds => place_472_preds,
      succs => place_472_succs,
      token => place_472_token,
      clk   => clk,
      reset => reset);

  place_473_preds(0) <= transition_469_symbol_out;
  place_473_succs(0) <= transition_470_symbol_out;
  place_473 : place
    generic map(marking => false)
    port map(
      preds => place_473_preds,
      succs => place_473_succs,
      token => place_473_token,
      clk   => clk,
      reset => reset);

  place_479_preds(0) <= transition_475_symbol_out;
  place_479_succs(0) <= transition_476_symbol_out;
  place_479 : place
    generic map(marking => false)
    port map(
      preds => place_479_preds,
      succs => place_479_succs,
      token => place_479_token,
      clk   => clk,
      reset => reset);

  place_480_preds(0) <= transition_476_symbol_out;
  place_480_succs(0) <= transition_477_symbol_out;
  place_480 : place
    generic map(marking => false)
    port map(
      preds => place_480_preds,
      succs => place_480_succs,
      token => place_480_token,
      clk   => clk,
      reset => reset);

  place_481_preds(0) <= transition_477_symbol_out;
  place_481_succs(0) <= transition_478_symbol_out;
  place_481 : place
    generic map(marking => false)
    port map(
      preds => place_481_preds,
      succs => place_481_succs,
      token => place_481_token,
      clk   => clk,
      reset => reset);

  place_486_preds(0) <= transition_482_symbol_out;
  place_486_succs(0) <= transition_483_symbol_out;
  place_486 : place
    generic map(marking => false)
    port map(
      preds => place_486_preds,
      succs => place_486_succs,
      token => place_486_token,
      clk   => clk,
      reset => reset);

  place_487_preds(0) <= transition_483_symbol_out;
  place_487_succs(0) <= transition_484_symbol_out;
  place_487 : place
    generic map(marking => false)
    port map(
      preds => place_487_preds,
      succs => place_487_succs,
      token => place_487_token,
      clk   => clk,
      reset => reset);

  place_488_preds(0) <= transition_484_symbol_out;
  place_488_succs(0) <= transition_485_symbol_out;
  place_488 : place
    generic map(marking => false)
    port map(
      preds => place_488_preds,
      succs => place_488_succs,
      token => place_488_token,
      clk   => clk,
      reset => reset);

  place_494_preds(0) <= transition_490_symbol_out;
  place_494_succs(0) <= transition_491_symbol_out;
  place_494 : place
    generic map(marking => false)
    port map(
      preds => place_494_preds,
      succs => place_494_succs,
      token => place_494_token,
      clk   => clk,
      reset => reset);

  place_495_preds(0) <= transition_491_symbol_out;
  place_495_succs(0) <= transition_492_symbol_out;
  place_495 : place
    generic map(marking => false)
    port map(
      preds => place_495_preds,
      succs => place_495_succs,
      token => place_495_token,
      clk   => clk,
      reset => reset);

  place_496_preds(0) <= transition_492_symbol_out;
  place_496_succs(0) <= transition_493_symbol_out;
  place_496 : place
    generic map(marking => false)
    port map(
      preds => place_496_preds,
      succs => place_496_succs,
      token => place_496_token,
      clk   => clk,
      reset => reset);

  place_497_preds(0) <= transition_499_symbol_out;
  place_497_succs(0) <= transition_498_symbol_out;
  place_497 : place
    generic map(marking => false)
    port map(
      preds => place_497_preds,
      succs => place_497_succs,
      token => place_497_token,
      clk   => clk,
      reset => reset);

  place_505_preds(0) <= transition_501_symbol_out;
  place_505_succs(0) <= transition_502_symbol_out;
  place_505 : place
    generic map(marking => false)
    port map(
      preds => place_505_preds,
      succs => place_505_succs,
      token => place_505_token,
      clk   => clk,
      reset => reset);

  place_506_preds(0) <= transition_502_symbol_out;
  place_506_succs(0) <= transition_503_symbol_out;
  place_506 : place
    generic map(marking => false)
    port map(
      preds => place_506_preds,
      succs => place_506_succs,
      token => place_506_token,
      clk   => clk,
      reset => reset);

  place_507_preds(0) <= transition_503_symbol_out;
  place_507_succs(0) <= transition_504_symbol_out;
  place_507 : place
    generic map(marking => false)
    port map(
      preds => place_507_preds,
      succs => place_507_succs,
      token => place_507_token,
      clk   => clk,
      reset => reset);

  place_512_preds(0) <= transition_508_symbol_out;
  place_512_succs(0) <= transition_509_symbol_out;
  place_512 : place
    generic map(marking => false)
    port map(
      preds => place_512_preds,
      succs => place_512_succs,
      token => place_512_token,
      clk   => clk,
      reset => reset);

  place_513_preds(0) <= transition_509_symbol_out;
  place_513_succs(0) <= transition_510_symbol_out;
  place_513 : place
    generic map(marking => false)
    port map(
      preds => place_513_preds,
      succs => place_513_succs,
      token => place_513_token,
      clk   => clk,
      reset => reset);

  place_514_preds(0) <= transition_510_symbol_out;
  place_514_succs(0) <= transition_511_symbol_out;
  place_514 : place
    generic map(marking => false)
    port map(
      preds => place_514_preds,
      succs => place_514_succs,
      token => place_514_token,
      clk   => clk,
      reset => reset);

  place_519_preds(0) <= transition_515_symbol_out;
  place_519_succs(0) <= transition_516_symbol_out;
  place_519 : place
    generic map(marking => false)
    port map(
      preds => place_519_preds,
      succs => place_519_succs,
      token => place_519_token,
      clk   => clk,
      reset => reset);

  place_520_preds(0) <= transition_516_symbol_out;
  place_520_succs(0) <= transition_517_symbol_out;
  place_520 : place
    generic map(marking => false)
    port map(
      preds => place_520_preds,
      succs => place_520_succs,
      token => place_520_token,
      clk   => clk,
      reset => reset);

  place_521_preds(0) <= transition_517_symbol_out;
  place_521_succs(0) <= transition_518_symbol_out;
  place_521 : place
    generic map(marking => false)
    port map(
      preds => place_521_preds,
      succs => place_521_succs,
      token => place_521_token,
      clk   => clk,
      reset => reset);

  place_527_preds(0) <= transition_523_symbol_out;
  place_527_succs(0) <= transition_524_symbol_out;
  place_527 : place
    generic map(marking => false)
    port map(
      preds => place_527_preds,
      succs => place_527_succs,
      token => place_527_token,
      clk   => clk,
      reset => reset);

  place_528_preds(0) <= transition_524_symbol_out;
  place_528_succs(0) <= transition_525_symbol_out;
  place_528 : place
    generic map(marking => false)
    port map(
      preds => place_528_preds,
      succs => place_528_succs,
      token => place_528_token,
      clk   => clk,
      reset => reset);

  place_529_preds(0) <= transition_525_symbol_out;
  place_529_succs(0) <= transition_526_symbol_out;
  place_529 : place
    generic map(marking => false)
    port map(
      preds => place_529_preds,
      succs => place_529_succs,
      token => place_529_token,
      clk   => clk,
      reset => reset);

  place_534_preds(0) <= transition_530_symbol_out;
  place_534_succs(0) <= transition_531_symbol_out;
  place_534 : place
    generic map(marking => false)
    port map(
      preds => place_534_preds,
      succs => place_534_succs,
      token => place_534_token,
      clk   => clk,
      reset => reset);

  place_535_preds(0) <= transition_531_symbol_out;
  place_535_succs(0) <= transition_532_symbol_out;
  place_535 : place
    generic map(marking => false)
    port map(
      preds => place_535_preds,
      succs => place_535_succs,
      token => place_535_token,
      clk   => clk,
      reset => reset);

  place_536_preds(0) <= transition_532_symbol_out;
  place_536_succs(0) <= transition_533_symbol_out;
  place_536 : place
    generic map(marking => false)
    port map(
      preds => place_536_preds,
      succs => place_536_succs,
      token => place_536_token,
      clk   => clk,
      reset => reset);

  place_542_preds(0) <= transition_538_symbol_out;
  place_542_succs(0) <= transition_539_symbol_out;
  place_542 : place
    generic map(marking => false)
    port map(
      preds => place_542_preds,
      succs => place_542_succs,
      token => place_542_token,
      clk   => clk,
      reset => reset);

  place_543_preds(0) <= transition_539_symbol_out;
  place_543_succs(0) <= transition_540_symbol_out;
  place_543 : place
    generic map(marking => false)
    port map(
      preds => place_543_preds,
      succs => place_543_succs,
      token => place_543_token,
      clk   => clk,
      reset => reset);

  place_544_preds(0) <= transition_540_symbol_out;
  place_544_succs(0) <= transition_541_symbol_out;
  place_544 : place
    generic map(marking => false)
    port map(
      preds => place_544_preds,
      succs => place_544_succs,
      token => place_544_token,
      clk   => clk,
      reset => reset);

  place_545_preds(0) <= transition_547_symbol_out;
  place_545_succs(0) <= transition_546_symbol_out;
  place_545 : place
    generic map(marking => false)
    port map(
      preds => place_545_preds,
      succs => place_545_succs,
      token => place_545_token,
      clk   => clk,
      reset => reset);

  place_553_preds(0) <= transition_549_symbol_out;
  place_553_succs(0) <= transition_550_symbol_out;
  place_553 : place
    generic map(marking => false)
    port map(
      preds => place_553_preds,
      succs => place_553_succs,
      token => place_553_token,
      clk   => clk,
      reset => reset);

  place_554_preds(0) <= transition_550_symbol_out;
  place_554_succs(0) <= transition_551_symbol_out;
  place_554 : place
    generic map(marking => false)
    port map(
      preds => place_554_preds,
      succs => place_554_succs,
      token => place_554_token,
      clk   => clk,
      reset => reset);

  place_555_preds(0) <= transition_551_symbol_out;
  place_555_succs(0) <= transition_552_symbol_out;
  place_555 : place
    generic map(marking => false)
    port map(
      preds => place_555_preds,
      succs => place_555_succs,
      token => place_555_token,
      clk   => clk,
      reset => reset);

  place_560_preds(0) <= transition_556_symbol_out;
  place_560_succs(0) <= transition_557_symbol_out;
  place_560 : place
    generic map(marking => false)
    port map(
      preds => place_560_preds,
      succs => place_560_succs,
      token => place_560_token,
      clk   => clk,
      reset => reset);

  place_561_preds(0) <= transition_557_symbol_out;
  place_561_succs(0) <= transition_558_symbol_out;
  place_561 : place
    generic map(marking => false)
    port map(
      preds => place_561_preds,
      succs => place_561_succs,
      token => place_561_token,
      clk   => clk,
      reset => reset);

  place_562_preds(0) <= transition_558_symbol_out;
  place_562_succs(0) <= transition_559_symbol_out;
  place_562 : place
    generic map(marking => false)
    port map(
      preds => place_562_preds,
      succs => place_562_succs,
      token => place_562_token,
      clk   => clk,
      reset => reset);

  place_567_preds(0) <= transition_563_symbol_out;
  place_567_succs(0) <= transition_564_symbol_out;
  place_567 : place
    generic map(marking => false)
    port map(
      preds => place_567_preds,
      succs => place_567_succs,
      token => place_567_token,
      clk   => clk,
      reset => reset);

  place_568_preds(0) <= transition_564_symbol_out;
  place_568_succs(0) <= transition_565_symbol_out;
  place_568 : place
    generic map(marking => false)
    port map(
      preds => place_568_preds,
      succs => place_568_succs,
      token => place_568_token,
      clk   => clk,
      reset => reset);

  place_569_preds(0) <= transition_565_symbol_out;
  place_569_succs(0) <= transition_566_symbol_out;
  place_569 : place
    generic map(marking => false)
    port map(
      preds => place_569_preds,
      succs => place_569_succs,
      token => place_569_token,
      clk   => clk,
      reset => reset);

  place_575_preds(0) <= transition_571_symbol_out;
  place_575_succs(0) <= transition_572_symbol_out;
  place_575 : place
    generic map(marking => false)
    port map(
      preds => place_575_preds,
      succs => place_575_succs,
      token => place_575_token,
      clk   => clk,
      reset => reset);

  place_576_preds(0) <= transition_572_symbol_out;
  place_576_succs(0) <= transition_573_symbol_out;
  place_576 : place
    generic map(marking => false)
    port map(
      preds => place_576_preds,
      succs => place_576_succs,
      token => place_576_token,
      clk   => clk,
      reset => reset);

  place_577_preds(0) <= transition_573_symbol_out;
  place_577_succs(0) <= transition_574_symbol_out;
  place_577 : place
    generic map(marking => false)
    port map(
      preds => place_577_preds,
      succs => place_577_succs,
      token => place_577_token,
      clk   => clk,
      reset => reset);

  place_582_preds(0) <= transition_578_symbol_out;
  place_582_succs(0) <= transition_579_symbol_out;
  place_582 : place
    generic map(marking => false)
    port map(
      preds => place_582_preds,
      succs => place_582_succs,
      token => place_582_token,
      clk   => clk,
      reset => reset);

  place_583_preds(0) <= transition_579_symbol_out;
  place_583_succs(0) <= transition_580_symbol_out;
  place_583 : place
    generic map(marking => false)
    port map(
      preds => place_583_preds,
      succs => place_583_succs,
      token => place_583_token,
      clk   => clk,
      reset => reset);

  place_584_preds(0) <= transition_580_symbol_out;
  place_584_succs(0) <= transition_581_symbol_out;
  place_584 : place
    generic map(marking => false)
    port map(
      preds => place_584_preds,
      succs => place_584_succs,
      token => place_584_token,
      clk   => clk,
      reset => reset);

  place_590_preds(0) <= transition_586_symbol_out;
  place_590_succs(0) <= transition_587_symbol_out;
  place_590 : place
    generic map(marking => false)
    port map(
      preds => place_590_preds,
      succs => place_590_succs,
      token => place_590_token,
      clk   => clk,
      reset => reset);

  place_591_preds(0) <= transition_587_symbol_out;
  place_591_succs(0) <= transition_588_symbol_out;
  place_591 : place
    generic map(marking => false)
    port map(
      preds => place_591_preds,
      succs => place_591_succs,
      token => place_591_token,
      clk   => clk,
      reset => reset);

  place_592_preds(0) <= transition_588_symbol_out;
  place_592_succs(0) <= transition_589_symbol_out;
  place_592 : place
    generic map(marking => false)
    port map(
      preds => place_592_preds,
      succs => place_592_succs,
      token => place_592_token,
      clk   => clk,
      reset => reset);

  place_593_preds(0) <= transition_595_symbol_out;
  place_593_succs(0) <= transition_594_symbol_out;
  place_593 : place
    generic map(marking => false)
    port map(
      preds => place_593_preds,
      succs => place_593_succs,
      token => place_593_token,
      clk   => clk,
      reset => reset);

  place_601_preds(0) <= transition_597_symbol_out;
  place_601_succs(0) <= transition_598_symbol_out;
  place_601 : place
    generic map(marking => false)
    port map(
      preds => place_601_preds,
      succs => place_601_succs,
      token => place_601_token,
      clk   => clk,
      reset => reset);

  place_602_preds(0) <= transition_598_symbol_out;
  place_602_succs(0) <= transition_599_symbol_out;
  place_602 : place
    generic map(marking => false)
    port map(
      preds => place_602_preds,
      succs => place_602_succs,
      token => place_602_token,
      clk   => clk,
      reset => reset);

  place_603_preds(0) <= transition_599_symbol_out;
  place_603_succs(0) <= transition_600_symbol_out;
  place_603 : place
    generic map(marking => false)
    port map(
      preds => place_603_preds,
      succs => place_603_succs,
      token => place_603_token,
      clk   => clk,
      reset => reset);

  place_608_preds(0) <= transition_604_symbol_out;
  place_608_succs(0) <= transition_605_symbol_out;
  place_608 : place
    generic map(marking => false)
    port map(
      preds => place_608_preds,
      succs => place_608_succs,
      token => place_608_token,
      clk   => clk,
      reset => reset);

  place_609_preds(0) <= transition_605_symbol_out;
  place_609_succs(0) <= transition_606_symbol_out;
  place_609 : place
    generic map(marking => false)
    port map(
      preds => place_609_preds,
      succs => place_609_succs,
      token => place_609_token,
      clk   => clk,
      reset => reset);

  place_610_preds(0) <= transition_606_symbol_out;
  place_610_succs(0) <= transition_607_symbol_out;
  place_610 : place
    generic map(marking => false)
    port map(
      preds => place_610_preds,
      succs => place_610_succs,
      token => place_610_token,
      clk   => clk,
      reset => reset);

  place_615_preds(0) <= transition_611_symbol_out;
  place_615_succs(0) <= transition_612_symbol_out;
  place_615 : place
    generic map(marking => false)
    port map(
      preds => place_615_preds,
      succs => place_615_succs,
      token => place_615_token,
      clk   => clk,
      reset => reset);

  place_616_preds(0) <= transition_612_symbol_out;
  place_616_succs(0) <= transition_613_symbol_out;
  place_616 : place
    generic map(marking => false)
    port map(
      preds => place_616_preds,
      succs => place_616_succs,
      token => place_616_token,
      clk   => clk,
      reset => reset);

  place_617_preds(0) <= transition_613_symbol_out;
  place_617_succs(0) <= transition_614_symbol_out;
  place_617 : place
    generic map(marking => false)
    port map(
      preds => place_617_preds,
      succs => place_617_succs,
      token => place_617_token,
      clk   => clk,
      reset => reset);

  place_623_preds(0) <= transition_619_symbol_out;
  place_623_succs(0) <= transition_620_symbol_out;
  place_623 : place
    generic map(marking => false)
    port map(
      preds => place_623_preds,
      succs => place_623_succs,
      token => place_623_token,
      clk   => clk,
      reset => reset);

  place_624_preds(0) <= transition_620_symbol_out;
  place_624_succs(0) <= transition_621_symbol_out;
  place_624 : place
    generic map(marking => false)
    port map(
      preds => place_624_preds,
      succs => place_624_succs,
      token => place_624_token,
      clk   => clk,
      reset => reset);

  place_625_preds(0) <= transition_621_symbol_out;
  place_625_succs(0) <= transition_622_symbol_out;
  place_625 : place
    generic map(marking => false)
    port map(
      preds => place_625_preds,
      succs => place_625_succs,
      token => place_625_token,
      clk   => clk,
      reset => reset);

  place_630_preds(0) <= transition_626_symbol_out;
  place_630_succs(0) <= transition_627_symbol_out;
  place_630 : place
    generic map(marking => false)
    port map(
      preds => place_630_preds,
      succs => place_630_succs,
      token => place_630_token,
      clk   => clk,
      reset => reset);

  place_631_preds(0) <= transition_627_symbol_out;
  place_631_succs(0) <= transition_628_symbol_out;
  place_631 : place
    generic map(marking => false)
    port map(
      preds => place_631_preds,
      succs => place_631_succs,
      token => place_631_token,
      clk   => clk,
      reset => reset);

  place_632_preds(0) <= transition_628_symbol_out;
  place_632_succs(0) <= transition_629_symbol_out;
  place_632 : place
    generic map(marking => false)
    port map(
      preds => place_632_preds,
      succs => place_632_succs,
      token => place_632_token,
      clk   => clk,
      reset => reset);

  place_638_preds(0) <= transition_634_symbol_out;
  place_638_succs(0) <= transition_635_symbol_out;
  place_638 : place
    generic map(marking => false)
    port map(
      preds => place_638_preds,
      succs => place_638_succs,
      token => place_638_token,
      clk   => clk,
      reset => reset);

  place_639_preds(0) <= transition_635_symbol_out;
  place_639_succs(0) <= transition_636_symbol_out;
  place_639 : place
    generic map(marking => false)
    port map(
      preds => place_639_preds,
      succs => place_639_succs,
      token => place_639_token,
      clk   => clk,
      reset => reset);

  place_640_preds(0) <= transition_636_symbol_out;
  place_640_succs(0) <= transition_637_symbol_out;
  place_640 : place
    generic map(marking => false)
    port map(
      preds => place_640_preds,
      succs => place_640_succs,
      token => place_640_token,
      clk   => clk,
      reset => reset);

  place_641_preds(0) <= transition_643_symbol_out;
  place_641_succs(0) <= transition_642_symbol_out;
  place_641 : place
    generic map(marking => false)
    port map(
      preds => place_641_preds,
      succs => place_641_succs,
      token => place_641_token,
      clk   => clk,
      reset => reset);

  place_649_preds(0) <= transition_645_symbol_out;
  place_649_succs(0) <= transition_646_symbol_out;
  place_649 : place
    generic map(marking => false)
    port map(
      preds => place_649_preds,
      succs => place_649_succs,
      token => place_649_token,
      clk   => clk,
      reset => reset);

  place_650_preds(0) <= transition_646_symbol_out;
  place_650_succs(0) <= transition_647_symbol_out;
  place_650 : place
    generic map(marking => false)
    port map(
      preds => place_650_preds,
      succs => place_650_succs,
      token => place_650_token,
      clk   => clk,
      reset => reset);

  place_651_preds(0) <= transition_647_symbol_out;
  place_651_succs(0) <= transition_648_symbol_out;
  place_651 : place
    generic map(marking => false)
    port map(
      preds => place_651_preds,
      succs => place_651_succs,
      token => place_651_token,
      clk   => clk,
      reset => reset);

  place_656_preds(0) <= transition_652_symbol_out;
  place_656_succs(0) <= transition_653_symbol_out;
  place_656 : place
    generic map(marking => false)
    port map(
      preds => place_656_preds,
      succs => place_656_succs,
      token => place_656_token,
      clk   => clk,
      reset => reset);

  place_657_preds(0) <= transition_653_symbol_out;
  place_657_succs(0) <= transition_654_symbol_out;
  place_657 : place
    generic map(marking => false)
    port map(
      preds => place_657_preds,
      succs => place_657_succs,
      token => place_657_token,
      clk   => clk,
      reset => reset);

  place_658_preds(0) <= transition_654_symbol_out;
  place_658_succs(0) <= transition_655_symbol_out;
  place_658 : place
    generic map(marking => false)
    port map(
      preds => place_658_preds,
      succs => place_658_succs,
      token => place_658_token,
      clk   => clk,
      reset => reset);

  place_663_preds(0) <= transition_659_symbol_out;
  place_663_succs(0) <= transition_660_symbol_out;
  place_663 : place
    generic map(marking => false)
    port map(
      preds => place_663_preds,
      succs => place_663_succs,
      token => place_663_token,
      clk   => clk,
      reset => reset);

  place_664_preds(0) <= transition_660_symbol_out;
  place_664_succs(0) <= transition_661_symbol_out;
  place_664 : place
    generic map(marking => false)
    port map(
      preds => place_664_preds,
      succs => place_664_succs,
      token => place_664_token,
      clk   => clk,
      reset => reset);

  place_665_preds(0) <= transition_661_symbol_out;
  place_665_succs(0) <= transition_662_symbol_out;
  place_665 : place
    generic map(marking => false)
    port map(
      preds => place_665_preds,
      succs => place_665_succs,
      token => place_665_token,
      clk   => clk,
      reset => reset);

  place_671_preds(0) <= transition_667_symbol_out;
  place_671_succs(0) <= transition_668_symbol_out;
  place_671 : place
    generic map(marking => false)
    port map(
      preds => place_671_preds,
      succs => place_671_succs,
      token => place_671_token,
      clk   => clk,
      reset => reset);

  place_672_preds(0) <= transition_668_symbol_out;
  place_672_succs(0) <= transition_669_symbol_out;
  place_672 : place
    generic map(marking => false)
    port map(
      preds => place_672_preds,
      succs => place_672_succs,
      token => place_672_token,
      clk   => clk,
      reset => reset);

  place_673_preds(0) <= transition_669_symbol_out;
  place_673_succs(0) <= transition_670_symbol_out;
  place_673 : place
    generic map(marking => false)
    port map(
      preds => place_673_preds,
      succs => place_673_succs,
      token => place_673_token,
      clk   => clk,
      reset => reset);

  place_678_preds(0) <= transition_674_symbol_out;
  place_678_succs(0) <= transition_675_symbol_out;
  place_678 : place
    generic map(marking => false)
    port map(
      preds => place_678_preds,
      succs => place_678_succs,
      token => place_678_token,
      clk   => clk,
      reset => reset);

  place_679_preds(0) <= transition_675_symbol_out;
  place_679_succs(0) <= transition_676_symbol_out;
  place_679 : place
    generic map(marking => false)
    port map(
      preds => place_679_preds,
      succs => place_679_succs,
      token => place_679_token,
      clk   => clk,
      reset => reset);

  place_680_preds(0) <= transition_676_symbol_out;
  place_680_succs(0) <= transition_677_symbol_out;
  place_680 : place
    generic map(marking => false)
    port map(
      preds => place_680_preds,
      succs => place_680_succs,
      token => place_680_token,
      clk   => clk,
      reset => reset);

  place_686_preds(0) <= transition_682_symbol_out;
  place_686_succs(0) <= transition_683_symbol_out;
  place_686 : place
    generic map(marking => false)
    port map(
      preds => place_686_preds,
      succs => place_686_succs,
      token => place_686_token,
      clk   => clk,
      reset => reset);

  place_687_preds(0) <= transition_683_symbol_out;
  place_687_succs(0) <= transition_684_symbol_out;
  place_687 : place
    generic map(marking => false)
    port map(
      preds => place_687_preds,
      succs => place_687_succs,
      token => place_687_token,
      clk   => clk,
      reset => reset);

  place_688_preds(0) <= transition_684_symbol_out;
  place_688_succs(0) <= transition_685_symbol_out;
  place_688 : place
    generic map(marking => false)
    port map(
      preds => place_688_preds,
      succs => place_688_succs,
      token => place_688_token,
      clk   => clk,
      reset => reset);

  place_689_preds(0) <= transition_691_symbol_out;
  place_689_succs(0) <= transition_690_symbol_out;
  place_689 : place
    generic map(marking => false)
    port map(
      preds => place_689_preds,
      succs => place_689_succs,
      token => place_689_token,
      clk   => clk,
      reset => reset);

  place_697_preds(0) <= transition_693_symbol_out;
  place_697_succs(0) <= transition_694_symbol_out;
  place_697 : place
    generic map(marking => false)
    port map(
      preds => place_697_preds,
      succs => place_697_succs,
      token => place_697_token,
      clk   => clk,
      reset => reset);

  place_698_preds(0) <= transition_694_symbol_out;
  place_698_succs(0) <= transition_695_symbol_out;
  place_698 : place
    generic map(marking => false)
    port map(
      preds => place_698_preds,
      succs => place_698_succs,
      token => place_698_token,
      clk   => clk,
      reset => reset);

  place_699_preds(0) <= transition_695_symbol_out;
  place_699_succs(0) <= transition_696_symbol_out;
  place_699 : place
    generic map(marking => false)
    port map(
      preds => place_699_preds,
      succs => place_699_succs,
      token => place_699_token,
      clk   => clk,
      reset => reset);

  place_704_preds(0) <= transition_700_symbol_out;
  place_704_succs(0) <= transition_701_symbol_out;
  place_704 : place
    generic map(marking => false)
    port map(
      preds => place_704_preds,
      succs => place_704_succs,
      token => place_704_token,
      clk   => clk,
      reset => reset);

  place_705_preds(0) <= transition_701_symbol_out;
  place_705_succs(0) <= transition_702_symbol_out;
  place_705 : place
    generic map(marking => false)
    port map(
      preds => place_705_preds,
      succs => place_705_succs,
      token => place_705_token,
      clk   => clk,
      reset => reset);

  place_706_preds(0) <= transition_702_symbol_out;
  place_706_succs(0) <= transition_703_symbol_out;
  place_706 : place
    generic map(marking => false)
    port map(
      preds => place_706_preds,
      succs => place_706_succs,
      token => place_706_token,
      clk   => clk,
      reset => reset);

  place_711_preds(0) <= transition_707_symbol_out;
  place_711_succs(0) <= transition_708_symbol_out;
  place_711 : place
    generic map(marking => false)
    port map(
      preds => place_711_preds,
      succs => place_711_succs,
      token => place_711_token,
      clk   => clk,
      reset => reset);

  place_712_preds(0) <= transition_708_symbol_out;
  place_712_succs(0) <= transition_709_symbol_out;
  place_712 : place
    generic map(marking => false)
    port map(
      preds => place_712_preds,
      succs => place_712_succs,
      token => place_712_token,
      clk   => clk,
      reset => reset);

  place_713_preds(0) <= transition_709_symbol_out;
  place_713_succs(0) <= transition_710_symbol_out;
  place_713 : place
    generic map(marking => false)
    port map(
      preds => place_713_preds,
      succs => place_713_succs,
      token => place_713_token,
      clk   => clk,
      reset => reset);

  place_719_preds(0) <= transition_715_symbol_out;
  place_719_succs(0) <= transition_716_symbol_out;
  place_719 : place
    generic map(marking => false)
    port map(
      preds => place_719_preds,
      succs => place_719_succs,
      token => place_719_token,
      clk   => clk,
      reset => reset);

  place_720_preds(0) <= transition_716_symbol_out;
  place_720_succs(0) <= transition_717_symbol_out;
  place_720 : place
    generic map(marking => false)
    port map(
      preds => place_720_preds,
      succs => place_720_succs,
      token => place_720_token,
      clk   => clk,
      reset => reset);

  place_721_preds(0) <= transition_717_symbol_out;
  place_721_succs(0) <= transition_718_symbol_out;
  place_721 : place
    generic map(marking => false)
    port map(
      preds => place_721_preds,
      succs => place_721_succs,
      token => place_721_token,
      clk   => clk,
      reset => reset);

  place_726_preds(0) <= transition_722_symbol_out;
  place_726_succs(0) <= transition_723_symbol_out;
  place_726 : place
    generic map(marking => false)
    port map(
      preds => place_726_preds,
      succs => place_726_succs,
      token => place_726_token,
      clk   => clk,
      reset => reset);

  place_727_preds(0) <= transition_723_symbol_out;
  place_727_succs(0) <= transition_724_symbol_out;
  place_727 : place
    generic map(marking => false)
    port map(
      preds => place_727_preds,
      succs => place_727_succs,
      token => place_727_token,
      clk   => clk,
      reset => reset);

  place_728_preds(0) <= transition_724_symbol_out;
  place_728_succs(0) <= transition_725_symbol_out;
  place_728 : place
    generic map(marking => false)
    port map(
      preds => place_728_preds,
      succs => place_728_succs,
      token => place_728_token,
      clk   => clk,
      reset => reset);

  place_734_preds(0) <= transition_730_symbol_out;
  place_734_succs(0) <= transition_731_symbol_out;
  place_734 : place
    generic map(marking => false)
    port map(
      preds => place_734_preds,
      succs => place_734_succs,
      token => place_734_token,
      clk   => clk,
      reset => reset);

  place_735_preds(0) <= transition_731_symbol_out;
  place_735_succs(0) <= transition_732_symbol_out;
  place_735 : place
    generic map(marking => false)
    port map(
      preds => place_735_preds,
      succs => place_735_succs,
      token => place_735_token,
      clk   => clk,
      reset => reset);

  place_736_preds(0) <= transition_732_symbol_out;
  place_736_succs(0) <= transition_733_symbol_out;
  place_736 : place
    generic map(marking => false)
    port map(
      preds => place_736_preds,
      succs => place_736_succs,
      token => place_736_token,
      clk   => clk,
      reset => reset);

  place_737_preds(0) <= transition_739_symbol_out;
  place_737_succs(0) <= transition_738_symbol_out;
  place_737 : place
    generic map(marking => false)
    port map(
      preds => place_737_preds,
      succs => place_737_succs,
      token => place_737_token,
      clk   => clk,
      reset => reset);

  place_745_preds(0) <= transition_741_symbol_out;
  place_745_succs(0) <= transition_742_symbol_out;
  place_745 : place
    generic map(marking => false)
    port map(
      preds => place_745_preds,
      succs => place_745_succs,
      token => place_745_token,
      clk   => clk,
      reset => reset);

  place_746_preds(0) <= transition_742_symbol_out;
  place_746_succs(0) <= transition_743_symbol_out;
  place_746 : place
    generic map(marking => false)
    port map(
      preds => place_746_preds,
      succs => place_746_succs,
      token => place_746_token,
      clk   => clk,
      reset => reset);

  place_747_preds(0) <= transition_743_symbol_out;
  place_747_succs(0) <= transition_744_symbol_out;
  place_747 : place
    generic map(marking => false)
    port map(
      preds => place_747_preds,
      succs => place_747_succs,
      token => place_747_token,
      clk   => clk,
      reset => reset);

  place_752_preds(0) <= transition_748_symbol_out;
  place_752_succs(0) <= transition_749_symbol_out;
  place_752 : place
    generic map(marking => false)
    port map(
      preds => place_752_preds,
      succs => place_752_succs,
      token => place_752_token,
      clk   => clk,
      reset => reset);

  place_753_preds(0) <= transition_749_symbol_out;
  place_753_succs(0) <= transition_750_symbol_out;
  place_753 : place
    generic map(marking => false)
    port map(
      preds => place_753_preds,
      succs => place_753_succs,
      token => place_753_token,
      clk   => clk,
      reset => reset);

  place_754_preds(0) <= transition_750_symbol_out;
  place_754_succs(0) <= transition_751_symbol_out;
  place_754 : place
    generic map(marking => false)
    port map(
      preds => place_754_preds,
      succs => place_754_succs,
      token => place_754_token,
      clk   => clk,
      reset => reset);

  place_759_preds(0) <= transition_755_symbol_out;
  place_759_succs(0) <= transition_756_symbol_out;
  place_759 : place
    generic map(marking => false)
    port map(
      preds => place_759_preds,
      succs => place_759_succs,
      token => place_759_token,
      clk   => clk,
      reset => reset);

  place_760_preds(0) <= transition_756_symbol_out;
  place_760_succs(0) <= transition_757_symbol_out;
  place_760 : place
    generic map(marking => false)
    port map(
      preds => place_760_preds,
      succs => place_760_succs,
      token => place_760_token,
      clk   => clk,
      reset => reset);

  place_761_preds(0) <= transition_757_symbol_out;
  place_761_succs(0) <= transition_758_symbol_out;
  place_761 : place
    generic map(marking => false)
    port map(
      preds => place_761_preds,
      succs => place_761_succs,
      token => place_761_token,
      clk   => clk,
      reset => reset);

  place_767_preds(0) <= transition_763_symbol_out;
  place_767_succs(0) <= transition_764_symbol_out;
  place_767 : place
    generic map(marking => false)
    port map(
      preds => place_767_preds,
      succs => place_767_succs,
      token => place_767_token,
      clk   => clk,
      reset => reset);

  place_768_preds(0) <= transition_764_symbol_out;
  place_768_succs(0) <= transition_765_symbol_out;
  place_768 : place
    generic map(marking => false)
    port map(
      preds => place_768_preds,
      succs => place_768_succs,
      token => place_768_token,
      clk   => clk,
      reset => reset);

  place_769_preds(0) <= transition_765_symbol_out;
  place_769_succs(0) <= transition_766_symbol_out;
  place_769 : place
    generic map(marking => false)
    port map(
      preds => place_769_preds,
      succs => place_769_succs,
      token => place_769_token,
      clk   => clk,
      reset => reset);

  place_774_preds(0) <= transition_770_symbol_out;
  place_774_succs(0) <= transition_771_symbol_out;
  place_774 : place
    generic map(marking => false)
    port map(
      preds => place_774_preds,
      succs => place_774_succs,
      token => place_774_token,
      clk   => clk,
      reset => reset);

  place_775_preds(0) <= transition_771_symbol_out;
  place_775_succs(0) <= transition_772_symbol_out;
  place_775 : place
    generic map(marking => false)
    port map(
      preds => place_775_preds,
      succs => place_775_succs,
      token => place_775_token,
      clk   => clk,
      reset => reset);

  place_776_preds(0) <= transition_772_symbol_out;
  place_776_succs(0) <= transition_773_symbol_out;
  place_776 : place
    generic map(marking => false)
    port map(
      preds => place_776_preds,
      succs => place_776_succs,
      token => place_776_token,
      clk   => clk,
      reset => reset);

  place_782_preds(0) <= transition_778_symbol_out;
  place_782_succs(0) <= transition_779_symbol_out;
  place_782 : place
    generic map(marking => false)
    port map(
      preds => place_782_preds,
      succs => place_782_succs,
      token => place_782_token,
      clk   => clk,
      reset => reset);

  place_783_preds(0) <= transition_779_symbol_out;
  place_783_succs(0) <= transition_780_symbol_out;
  place_783 : place
    generic map(marking => false)
    port map(
      preds => place_783_preds,
      succs => place_783_succs,
      token => place_783_token,
      clk   => clk,
      reset => reset);

  place_784_preds(0) <= transition_780_symbol_out;
  place_784_succs(0) <= transition_781_symbol_out;
  place_784 : place
    generic map(marking => false)
    port map(
      preds => place_784_preds,
      succs => place_784_succs,
      token => place_784_token,
      clk   => clk,
      reset => reset);

  place_785_preds(0) <= transition_787_symbol_out;
  place_785_succs(0) <= transition_786_symbol_out;
  place_785 : place
    generic map(marking => false)
    port map(
      preds => place_785_preds,
      succs => place_785_succs,
      token => place_785_token,
      clk   => clk,
      reset => reset);

  place_793_preds(0) <= transition_789_symbol_out;
  place_793_succs(0) <= transition_790_symbol_out;
  place_793 : place
    generic map(marking => false)
    port map(
      preds => place_793_preds,
      succs => place_793_succs,
      token => place_793_token,
      clk   => clk,
      reset => reset);

  place_794_preds(0) <= transition_790_symbol_out;
  place_794_succs(0) <= transition_791_symbol_out;
  place_794 : place
    generic map(marking => false)
    port map(
      preds => place_794_preds,
      succs => place_794_succs,
      token => place_794_token,
      clk   => clk,
      reset => reset);

  place_795_preds(0) <= transition_791_symbol_out;
  place_795_succs(0) <= transition_792_symbol_out;
  place_795 : place
    generic map(marking => false)
    port map(
      preds => place_795_preds,
      succs => place_795_succs,
      token => place_795_token,
      clk   => clk,
      reset => reset);

  place_800_preds(0) <= transition_796_symbol_out;
  place_800_succs(0) <= transition_797_symbol_out;
  place_800 : place
    generic map(marking => false)
    port map(
      preds => place_800_preds,
      succs => place_800_succs,
      token => place_800_token,
      clk   => clk,
      reset => reset);

  place_801_preds(0) <= transition_797_symbol_out;
  place_801_succs(0) <= transition_798_symbol_out;
  place_801 : place
    generic map(marking => false)
    port map(
      preds => place_801_preds,
      succs => place_801_succs,
      token => place_801_token,
      clk   => clk,
      reset => reset);

  place_802_preds(0) <= transition_798_symbol_out;
  place_802_succs(0) <= transition_799_symbol_out;
  place_802 : place
    generic map(marking => false)
    port map(
      preds => place_802_preds,
      succs => place_802_succs,
      token => place_802_token,
      clk   => clk,
      reset => reset);

  place_807_preds(0) <= transition_803_symbol_out;
  place_807_succs(0) <= transition_804_symbol_out;
  place_807 : place
    generic map(marking => false)
    port map(
      preds => place_807_preds,
      succs => place_807_succs,
      token => place_807_token,
      clk   => clk,
      reset => reset);

  place_808_preds(0) <= transition_804_symbol_out;
  place_808_succs(0) <= transition_805_symbol_out;
  place_808 : place
    generic map(marking => false)
    port map(
      preds => place_808_preds,
      succs => place_808_succs,
      token => place_808_token,
      clk   => clk,
      reset => reset);

  place_809_preds(0) <= transition_805_symbol_out;
  place_809_succs(0) <= transition_806_symbol_out;
  place_809 : place
    generic map(marking => false)
    port map(
      preds => place_809_preds,
      succs => place_809_succs,
      token => place_809_token,
      clk   => clk,
      reset => reset);

  place_815_preds(0) <= transition_811_symbol_out;
  place_815_succs(0) <= transition_812_symbol_out;
  place_815 : place
    generic map(marking => false)
    port map(
      preds => place_815_preds,
      succs => place_815_succs,
      token => place_815_token,
      clk   => clk,
      reset => reset);

  place_816_preds(0) <= transition_812_symbol_out;
  place_816_succs(0) <= transition_813_symbol_out;
  place_816 : place
    generic map(marking => false)
    port map(
      preds => place_816_preds,
      succs => place_816_succs,
      token => place_816_token,
      clk   => clk,
      reset => reset);

  place_817_preds(0) <= transition_813_symbol_out;
  place_817_succs(0) <= transition_814_symbol_out;
  place_817 : place
    generic map(marking => false)
    port map(
      preds => place_817_preds,
      succs => place_817_succs,
      token => place_817_token,
      clk   => clk,
      reset => reset);

  place_822_preds(0) <= transition_818_symbol_out;
  place_822_succs(0) <= transition_819_symbol_out;
  place_822 : place
    generic map(marking => false)
    port map(
      preds => place_822_preds,
      succs => place_822_succs,
      token => place_822_token,
      clk   => clk,
      reset => reset);

  place_823_preds(0) <= transition_819_symbol_out;
  place_823_succs(0) <= transition_820_symbol_out;
  place_823 : place
    generic map(marking => false)
    port map(
      preds => place_823_preds,
      succs => place_823_succs,
      token => place_823_token,
      clk   => clk,
      reset => reset);

  place_824_preds(0) <= transition_820_symbol_out;
  place_824_succs(0) <= transition_821_symbol_out;
  place_824 : place
    generic map(marking => false)
    port map(
      preds => place_824_preds,
      succs => place_824_succs,
      token => place_824_token,
      clk   => clk,
      reset => reset);

  place_830_preds(0) <= transition_826_symbol_out;
  place_830_succs(0) <= transition_827_symbol_out;
  place_830 : place
    generic map(marking => false)
    port map(
      preds => place_830_preds,
      succs => place_830_succs,
      token => place_830_token,
      clk   => clk,
      reset => reset);

  place_831_preds(0) <= transition_827_symbol_out;
  place_831_succs(0) <= transition_828_symbol_out;
  place_831 : place
    generic map(marking => false)
    port map(
      preds => place_831_preds,
      succs => place_831_succs,
      token => place_831_token,
      clk   => clk,
      reset => reset);

  place_832_preds(0) <= transition_828_symbol_out;
  place_832_succs(0) <= transition_829_symbol_out;
  place_832 : place
    generic map(marking => false)
    port map(
      preds => place_832_preds,
      succs => place_832_succs,
      token => place_832_token,
      clk   => clk,
      reset => reset);

  place_833_preds(0) <= transition_835_symbol_out;
  place_833_succs(0) <= transition_834_symbol_out;
  place_833 : place
    generic map(marking => false)
    port map(
      preds => place_833_preds,
      succs => place_833_succs,
      token => place_833_token,
      clk   => clk,
      reset => reset);

  place_841_preds(0) <= transition_837_symbol_out;
  place_841_succs(0) <= transition_838_symbol_out;
  place_841 : place
    generic map(marking => false)
    port map(
      preds => place_841_preds,
      succs => place_841_succs,
      token => place_841_token,
      clk   => clk,
      reset => reset);

  place_842_preds(0) <= transition_838_symbol_out;
  place_842_succs(0) <= transition_839_symbol_out;
  place_842 : place
    generic map(marking => false)
    port map(
      preds => place_842_preds,
      succs => place_842_succs,
      token => place_842_token,
      clk   => clk,
      reset => reset);

  place_843_preds(0) <= transition_839_symbol_out;
  place_843_succs(0) <= transition_840_symbol_out;
  place_843 : place
    generic map(marking => false)
    port map(
      preds => place_843_preds,
      succs => place_843_succs,
      token => place_843_token,
      clk   => clk,
      reset => reset);

  place_848_preds(0) <= transition_844_symbol_out;
  place_848_succs(0) <= transition_845_symbol_out;
  place_848 : place
    generic map(marking => false)
    port map(
      preds => place_848_preds,
      succs => place_848_succs,
      token => place_848_token,
      clk   => clk,
      reset => reset);

  place_849_preds(0) <= transition_845_symbol_out;
  place_849_succs(0) <= transition_846_symbol_out;
  place_849 : place
    generic map(marking => false)
    port map(
      preds => place_849_preds,
      succs => place_849_succs,
      token => place_849_token,
      clk   => clk,
      reset => reset);

  place_850_preds(0) <= transition_846_symbol_out;
  place_850_succs(0) <= transition_847_symbol_out;
  place_850 : place
    generic map(marking => false)
    port map(
      preds => place_850_preds,
      succs => place_850_succs,
      token => place_850_token,
      clk   => clk,
      reset => reset);

  place_855_preds(0) <= transition_851_symbol_out;
  place_855_succs(0) <= transition_852_symbol_out;
  place_855 : place
    generic map(marking => false)
    port map(
      preds => place_855_preds,
      succs => place_855_succs,
      token => place_855_token,
      clk   => clk,
      reset => reset);

  place_856_preds(0) <= transition_852_symbol_out;
  place_856_succs(0) <= transition_853_symbol_out;
  place_856 : place
    generic map(marking => false)
    port map(
      preds => place_856_preds,
      succs => place_856_succs,
      token => place_856_token,
      clk   => clk,
      reset => reset);

  place_857_preds(0) <= transition_853_symbol_out;
  place_857_succs(0) <= transition_854_symbol_out;
  place_857 : place
    generic map(marking => false)
    port map(
      preds => place_857_preds,
      succs => place_857_succs,
      token => place_857_token,
      clk   => clk,
      reset => reset);

  place_863_preds(0) <= transition_859_symbol_out;
  place_863_succs(0) <= transition_860_symbol_out;
  place_863 : place
    generic map(marking => false)
    port map(
      preds => place_863_preds,
      succs => place_863_succs,
      token => place_863_token,
      clk   => clk,
      reset => reset);

  place_864_preds(0) <= transition_860_symbol_out;
  place_864_succs(0) <= transition_861_symbol_out;
  place_864 : place
    generic map(marking => false)
    port map(
      preds => place_864_preds,
      succs => place_864_succs,
      token => place_864_token,
      clk   => clk,
      reset => reset);

  place_865_preds(0) <= transition_861_symbol_out;
  place_865_succs(0) <= transition_862_symbol_out;
  place_865 : place
    generic map(marking => false)
    port map(
      preds => place_865_preds,
      succs => place_865_succs,
      token => place_865_token,
      clk   => clk,
      reset => reset);

  place_870_preds(0) <= transition_866_symbol_out;
  place_870_succs(0) <= transition_867_symbol_out;
  place_870 : place
    generic map(marking => false)
    port map(
      preds => place_870_preds,
      succs => place_870_succs,
      token => place_870_token,
      clk   => clk,
      reset => reset);

  place_871_preds(0) <= transition_867_symbol_out;
  place_871_succs(0) <= transition_868_symbol_out;
  place_871 : place
    generic map(marking => false)
    port map(
      preds => place_871_preds,
      succs => place_871_succs,
      token => place_871_token,
      clk   => clk,
      reset => reset);

  place_872_preds(0) <= transition_868_symbol_out;
  place_872_succs(0) <= transition_869_symbol_out;
  place_872 : place
    generic map(marking => false)
    port map(
      preds => place_872_preds,
      succs => place_872_succs,
      token => place_872_token,
      clk   => clk,
      reset => reset);

  place_878_preds(0) <= transition_874_symbol_out;
  place_878_succs(0) <= transition_875_symbol_out;
  place_878 : place
    generic map(marking => false)
    port map(
      preds => place_878_preds,
      succs => place_878_succs,
      token => place_878_token,
      clk   => clk,
      reset => reset);

  place_879_preds(0) <= transition_875_symbol_out;
  place_879_succs(0) <= transition_876_symbol_out;
  place_879 : place
    generic map(marking => false)
    port map(
      preds => place_879_preds,
      succs => place_879_succs,
      token => place_879_token,
      clk   => clk,
      reset => reset);

  place_880_preds(0) <= transition_876_symbol_out;
  place_880_succs(0) <= transition_877_symbol_out;
  place_880 : place
    generic map(marking => false)
    port map(
      preds => place_880_preds,
      succs => place_880_succs,
      token => place_880_token,
      clk   => clk,
      reset => reset);

  place_881_preds(0) <= transition_883_symbol_out;
  place_881_succs(0) <= transition_882_symbol_out;
  place_881 : place
    generic map(marking => false)
    port map(
      preds => place_881_preds,
      succs => place_881_succs,
      token => place_881_token,
      clk   => clk,
      reset => reset);

  place_889_preds(0) <= transition_885_symbol_out;
  place_889_succs(0) <= transition_886_symbol_out;
  place_889 : place
    generic map(marking => false)
    port map(
      preds => place_889_preds,
      succs => place_889_succs,
      token => place_889_token,
      clk   => clk,
      reset => reset);

  place_890_preds(0) <= transition_886_symbol_out;
  place_890_succs(0) <= transition_887_symbol_out;
  place_890 : place
    generic map(marking => false)
    port map(
      preds => place_890_preds,
      succs => place_890_succs,
      token => place_890_token,
      clk   => clk,
      reset => reset);

  place_891_preds(0) <= transition_887_symbol_out;
  place_891_succs(0) <= transition_888_symbol_out;
  place_891 : place
    generic map(marking => false)
    port map(
      preds => place_891_preds,
      succs => place_891_succs,
      token => place_891_token,
      clk   => clk,
      reset => reset);

  place_896_preds(0) <= transition_892_symbol_out;
  place_896_succs(0) <= transition_893_symbol_out;
  place_896 : place
    generic map(marking => false)
    port map(
      preds => place_896_preds,
      succs => place_896_succs,
      token => place_896_token,
      clk   => clk,
      reset => reset);

  place_897_preds(0) <= transition_893_symbol_out;
  place_897_succs(0) <= transition_894_symbol_out;
  place_897 : place
    generic map(marking => false)
    port map(
      preds => place_897_preds,
      succs => place_897_succs,
      token => place_897_token,
      clk   => clk,
      reset => reset);

  place_898_preds(0) <= transition_894_symbol_out;
  place_898_succs(0) <= transition_895_symbol_out;
  place_898 : place
    generic map(marking => false)
    port map(
      preds => place_898_preds,
      succs => place_898_succs,
      token => place_898_token,
      clk   => clk,
      reset => reset);

  place_903_preds(0) <= transition_899_symbol_out;
  place_903_succs(0) <= transition_900_symbol_out;
  place_903 : place
    generic map(marking => false)
    port map(
      preds => place_903_preds,
      succs => place_903_succs,
      token => place_903_token,
      clk   => clk,
      reset => reset);

  place_904_preds(0) <= transition_900_symbol_out;
  place_904_succs(0) <= transition_901_symbol_out;
  place_904 : place
    generic map(marking => false)
    port map(
      preds => place_904_preds,
      succs => place_904_succs,
      token => place_904_token,
      clk   => clk,
      reset => reset);

  place_905_preds(0) <= transition_901_symbol_out;
  place_905_succs(0) <= transition_902_symbol_out;
  place_905 : place
    generic map(marking => false)
    port map(
      preds => place_905_preds,
      succs => place_905_succs,
      token => place_905_token,
      clk   => clk,
      reset => reset);

  place_911_preds(0) <= transition_907_symbol_out;
  place_911_succs(0) <= transition_908_symbol_out;
  place_911 : place
    generic map(marking => false)
    port map(
      preds => place_911_preds,
      succs => place_911_succs,
      token => place_911_token,
      clk   => clk,
      reset => reset);

  place_912_preds(0) <= transition_908_symbol_out;
  place_912_succs(0) <= transition_909_symbol_out;
  place_912 : place
    generic map(marking => false)
    port map(
      preds => place_912_preds,
      succs => place_912_succs,
      token => place_912_token,
      clk   => clk,
      reset => reset);

  place_913_preds(0) <= transition_909_symbol_out;
  place_913_succs(0) <= transition_910_symbol_out;
  place_913 : place
    generic map(marking => false)
    port map(
      preds => place_913_preds,
      succs => place_913_succs,
      token => place_913_token,
      clk   => clk,
      reset => reset);

  place_918_preds(0) <= transition_914_symbol_out;
  place_918_succs(0) <= transition_915_symbol_out;
  place_918 : place
    generic map(marking => false)
    port map(
      preds => place_918_preds,
      succs => place_918_succs,
      token => place_918_token,
      clk   => clk,
      reset => reset);

  place_919_preds(0) <= transition_915_symbol_out;
  place_919_succs(0) <= transition_916_symbol_out;
  place_919 : place
    generic map(marking => false)
    port map(
      preds => place_919_preds,
      succs => place_919_succs,
      token => place_919_token,
      clk   => clk,
      reset => reset);

  place_920_preds(0) <= transition_916_symbol_out;
  place_920_succs(0) <= transition_917_symbol_out;
  place_920 : place
    generic map(marking => false)
    port map(
      preds => place_920_preds,
      succs => place_920_succs,
      token => place_920_token,
      clk   => clk,
      reset => reset);

  place_926_preds(0) <= transition_922_symbol_out;
  place_926_succs(0) <= transition_923_symbol_out;
  place_926 : place
    generic map(marking => false)
    port map(
      preds => place_926_preds,
      succs => place_926_succs,
      token => place_926_token,
      clk   => clk,
      reset => reset);

  place_927_preds(0) <= transition_923_symbol_out;
  place_927_succs(0) <= transition_924_symbol_out;
  place_927 : place
    generic map(marking => false)
    port map(
      preds => place_927_preds,
      succs => place_927_succs,
      token => place_927_token,
      clk   => clk,
      reset => reset);

  place_928_preds(0) <= transition_924_symbol_out;
  place_928_succs(0) <= transition_925_symbol_out;
  place_928 : place
    generic map(marking => false)
    port map(
      preds => place_928_preds,
      succs => place_928_succs,
      token => place_928_token,
      clk   => clk,
      reset => reset);

  place_929_preds(0) <= transition_931_symbol_out;
  place_929_succs(0) <= transition_930_symbol_out;
  place_929 : place
    generic map(marking => false)
    port map(
      preds => place_929_preds,
      succs => place_929_succs,
      token => place_929_token,
      clk   => clk,
      reset => reset);

  place_937_preds(0) <= transition_933_symbol_out;
  place_937_succs(0) <= transition_934_symbol_out;
  place_937 : place
    generic map(marking => false)
    port map(
      preds => place_937_preds,
      succs => place_937_succs,
      token => place_937_token,
      clk   => clk,
      reset => reset);

  place_938_preds(0) <= transition_934_symbol_out;
  place_938_succs(0) <= transition_935_symbol_out;
  place_938 : place
    generic map(marking => false)
    port map(
      preds => place_938_preds,
      succs => place_938_succs,
      token => place_938_token,
      clk   => clk,
      reset => reset);

  place_939_preds(0) <= transition_935_symbol_out;
  place_939_succs(0) <= transition_936_symbol_out;
  place_939 : place
    generic map(marking => false)
    port map(
      preds => place_939_preds,
      succs => place_939_succs,
      token => place_939_token,
      clk   => clk,
      reset => reset);

  place_944_preds(0) <= transition_940_symbol_out;
  place_944_succs(0) <= transition_941_symbol_out;
  place_944 : place
    generic map(marking => false)
    port map(
      preds => place_944_preds,
      succs => place_944_succs,
      token => place_944_token,
      clk   => clk,
      reset => reset);

  place_945_preds(0) <= transition_941_symbol_out;
  place_945_succs(0) <= transition_942_symbol_out;
  place_945 : place
    generic map(marking => false)
    port map(
      preds => place_945_preds,
      succs => place_945_succs,
      token => place_945_token,
      clk   => clk,
      reset => reset);

  place_946_preds(0) <= transition_942_symbol_out;
  place_946_succs(0) <= transition_943_symbol_out;
  place_946 : place
    generic map(marking => false)
    port map(
      preds => place_946_preds,
      succs => place_946_succs,
      token => place_946_token,
      clk   => clk,
      reset => reset);

  place_951_preds(0) <= transition_947_symbol_out;
  place_951_succs(0) <= transition_948_symbol_out;
  place_951 : place
    generic map(marking => false)
    port map(
      preds => place_951_preds,
      succs => place_951_succs,
      token => place_951_token,
      clk   => clk,
      reset => reset);

  place_952_preds(0) <= transition_948_symbol_out;
  place_952_succs(0) <= transition_949_symbol_out;
  place_952 : place
    generic map(marking => false)
    port map(
      preds => place_952_preds,
      succs => place_952_succs,
      token => place_952_token,
      clk   => clk,
      reset => reset);

  place_953_preds(0) <= transition_949_symbol_out;
  place_953_succs(0) <= transition_950_symbol_out;
  place_953 : place
    generic map(marking => false)
    port map(
      preds => place_953_preds,
      succs => place_953_succs,
      token => place_953_token,
      clk   => clk,
      reset => reset);

  place_959_preds(0) <= transition_955_symbol_out;
  place_959_succs(0) <= transition_956_symbol_out;
  place_959 : place
    generic map(marking => false)
    port map(
      preds => place_959_preds,
      succs => place_959_succs,
      token => place_959_token,
      clk   => clk,
      reset => reset);

  place_960_preds(0) <= transition_956_symbol_out;
  place_960_succs(0) <= transition_957_symbol_out;
  place_960 : place
    generic map(marking => false)
    port map(
      preds => place_960_preds,
      succs => place_960_succs,
      token => place_960_token,
      clk   => clk,
      reset => reset);

  place_961_preds(0) <= transition_957_symbol_out;
  place_961_succs(0) <= transition_958_symbol_out;
  place_961 : place
    generic map(marking => false)
    port map(
      preds => place_961_preds,
      succs => place_961_succs,
      token => place_961_token,
      clk   => clk,
      reset => reset);

  place_966_preds(0) <= transition_962_symbol_out;
  place_966_succs(0) <= transition_963_symbol_out;
  place_966 : place
    generic map(marking => false)
    port map(
      preds => place_966_preds,
      succs => place_966_succs,
      token => place_966_token,
      clk   => clk,
      reset => reset);

  place_967_preds(0) <= transition_963_symbol_out;
  place_967_succs(0) <= transition_964_symbol_out;
  place_967 : place
    generic map(marking => false)
    port map(
      preds => place_967_preds,
      succs => place_967_succs,
      token => place_967_token,
      clk   => clk,
      reset => reset);

  place_968_preds(0) <= transition_964_symbol_out;
  place_968_succs(0) <= transition_965_symbol_out;
  place_968 : place
    generic map(marking => false)
    port map(
      preds => place_968_preds,
      succs => place_968_succs,
      token => place_968_token,
      clk   => clk,
      reset => reset);

  place_974_preds(0) <= transition_970_symbol_out;
  place_974_succs(0) <= transition_971_symbol_out;
  place_974 : place
    generic map(marking => false)
    port map(
      preds => place_974_preds,
      succs => place_974_succs,
      token => place_974_token,
      clk   => clk,
      reset => reset);

  place_975_preds(0) <= transition_971_symbol_out;
  place_975_succs(0) <= transition_972_symbol_out;
  place_975 : place
    generic map(marking => false)
    port map(
      preds => place_975_preds,
      succs => place_975_succs,
      token => place_975_token,
      clk   => clk,
      reset => reset);

  place_976_preds(0) <= transition_972_symbol_out;
  place_976_succs(0) <= transition_973_symbol_out;
  place_976 : place
    generic map(marking => false)
    port map(
      preds => place_976_preds,
      succs => place_976_succs,
      token => place_976_token,
      clk   => clk,
      reset => reset);

  place_977_preds(0) <= transition_979_symbol_out;
  place_977_succs(0) <= transition_978_symbol_out;
  place_977 : place
    generic map(marking => false)
    port map(
      preds => place_977_preds,
      succs => place_977_succs,
      token => place_977_token,
      clk   => clk,
      reset => reset);

  place_985_preds(0) <= transition_981_symbol_out;
  place_985_succs(0) <= transition_982_symbol_out;
  place_985 : place
    generic map(marking => false)
    port map(
      preds => place_985_preds,
      succs => place_985_succs,
      token => place_985_token,
      clk   => clk,
      reset => reset);

  place_986_preds(0) <= transition_982_symbol_out;
  place_986_succs(0) <= transition_983_symbol_out;
  place_986 : place
    generic map(marking => false)
    port map(
      preds => place_986_preds,
      succs => place_986_succs,
      token => place_986_token,
      clk   => clk,
      reset => reset);

  place_987_preds(0) <= transition_983_symbol_out;
  place_987_succs(0) <= transition_984_symbol_out;
  place_987 : place
    generic map(marking => false)
    port map(
      preds => place_987_preds,
      succs => place_987_succs,
      token => place_987_token,
      clk   => clk,
      reset => reset);

  place_992_preds(0) <= transition_988_symbol_out;
  place_992_succs(0) <= transition_989_symbol_out;
  place_992 : place
    generic map(marking => false)
    port map(
      preds => place_992_preds,
      succs => place_992_succs,
      token => place_992_token,
      clk   => clk,
      reset => reset);

  place_993_preds(0) <= transition_989_symbol_out;
  place_993_succs(0) <= transition_990_symbol_out;
  place_993 : place
    generic map(marking => false)
    port map(
      preds => place_993_preds,
      succs => place_993_succs,
      token => place_993_token,
      clk   => clk,
      reset => reset);

  place_994_preds(0) <= transition_990_symbol_out;
  place_994_succs(0) <= transition_991_symbol_out;
  place_994 : place
    generic map(marking => false)
    port map(
      preds => place_994_preds,
      succs => place_994_succs,
      token => place_994_token,
      clk   => clk,
      reset => reset);

  place_999_preds(0) <= transition_995_symbol_out;
  place_999_succs(0) <= transition_996_symbol_out;
  place_999 : place
    generic map(marking => false)
    port map(
      preds => place_999_preds,
      succs => place_999_succs,
      token => place_999_token,
      clk   => clk,
      reset => reset);

  place_1000_preds(0) <= transition_996_symbol_out;
  place_1000_succs(0) <= transition_997_symbol_out;
  place_1000 : place
    generic map(marking => false)
    port map(
      preds => place_1000_preds,
      succs => place_1000_succs,
      token => place_1000_token,
      clk   => clk,
      reset => reset);

  place_1001_preds(0) <= transition_997_symbol_out;
  place_1001_succs(0) <= transition_998_symbol_out;
  place_1001 : place
    generic map(marking => false)
    port map(
      preds => place_1001_preds,
      succs => place_1001_succs,
      token => place_1001_token,
      clk   => clk,
      reset => reset);

  place_1007_preds(0) <= transition_1003_symbol_out;
  place_1007_succs(0) <= transition_1004_symbol_out;
  place_1007 : place
    generic map(marking => false)
    port map(
      preds => place_1007_preds,
      succs => place_1007_succs,
      token => place_1007_token,
      clk   => clk,
      reset => reset);

  place_1008_preds(0) <= transition_1004_symbol_out;
  place_1008_succs(0) <= transition_1005_symbol_out;
  place_1008 : place
    generic map(marking => false)
    port map(
      preds => place_1008_preds,
      succs => place_1008_succs,
      token => place_1008_token,
      clk   => clk,
      reset => reset);

  place_1009_preds(0) <= transition_1005_symbol_out;
  place_1009_succs(0) <= transition_1006_symbol_out;
  place_1009 : place
    generic map(marking => false)
    port map(
      preds => place_1009_preds,
      succs => place_1009_succs,
      token => place_1009_token,
      clk   => clk,
      reset => reset);

  place_1014_preds(0) <= transition_1010_symbol_out;
  place_1014_succs(0) <= transition_1011_symbol_out;
  place_1014 : place
    generic map(marking => false)
    port map(
      preds => place_1014_preds,
      succs => place_1014_succs,
      token => place_1014_token,
      clk   => clk,
      reset => reset);

  place_1015_preds(0) <= transition_1011_symbol_out;
  place_1015_succs(0) <= transition_1012_symbol_out;
  place_1015 : place
    generic map(marking => false)
    port map(
      preds => place_1015_preds,
      succs => place_1015_succs,
      token => place_1015_token,
      clk   => clk,
      reset => reset);

  place_1016_preds(0) <= transition_1012_symbol_out;
  place_1016_succs(0) <= transition_1013_symbol_out;
  place_1016 : place
    generic map(marking => false)
    port map(
      preds => place_1016_preds,
      succs => place_1016_succs,
      token => place_1016_token,
      clk   => clk,
      reset => reset);

  place_1022_preds(0) <= transition_1018_symbol_out;
  place_1022_succs(0) <= transition_1019_symbol_out;
  place_1022 : place
    generic map(marking => false)
    port map(
      preds => place_1022_preds,
      succs => place_1022_succs,
      token => place_1022_token,
      clk   => clk,
      reset => reset);

  place_1023_preds(0) <= transition_1019_symbol_out;
  place_1023_succs(0) <= transition_1020_symbol_out;
  place_1023 : place
    generic map(marking => false)
    port map(
      preds => place_1023_preds,
      succs => place_1023_succs,
      token => place_1023_token,
      clk   => clk,
      reset => reset);

  place_1024_preds(0) <= transition_1020_symbol_out;
  place_1024_succs(0) <= transition_1021_symbol_out;
  place_1024 : place
    generic map(marking => false)
    port map(
      preds => place_1024_preds,
      succs => place_1024_succs,
      token => place_1024_token,
      clk   => clk,
      reset => reset);

  place_1025_preds(0) <= transition_1027_symbol_out;
  place_1025_succs(0) <= transition_1026_symbol_out;
  place_1025 : place
    generic map(marking => false)
    port map(
      preds => place_1025_preds,
      succs => place_1025_succs,
      token => place_1025_token,
      clk   => clk,
      reset => reset);

  place_1029_preds(0) <= transition_1031_symbol_out;
  place_1029_succs(0) <= transition_1030_symbol_out;
  place_1029 : place
    generic map(marking => false)
    port map(
      preds => place_1029_preds,
      succs => place_1029_succs,
      token => place_1029_token,
      clk   => clk,
      reset => reset);

  place_1032_preds(0) <= transition_1034_symbol_out;
  place_1032_succs(0) <= transition_1033_symbol_out;
  place_1032 : place
    generic map(marking => false)
    port map(
      preds => place_1032_preds,
      succs => place_1032_succs,
      token => place_1032_token,
      clk   => clk,
      reset => reset);

  place_1036_preds(0) <= transition_1038_symbol_out;
  place_1036_succs(0) <= transition_1037_symbol_out;
  place_1036 : place
    generic map(marking => false)
    port map(
      preds => place_1036_preds,
      succs => place_1036_succs,
      token => place_1036_token,
      clk   => clk,
      reset => reset);

  place_1039_preds(0) <= transition_1041_symbol_out;
  place_1039_succs(0) <= transition_1040_symbol_out;
  place_1039 : place
    generic map(marking => false)
    port map(
      preds => place_1039_preds,
      succs => place_1039_succs,
      token => place_1039_token,
      clk   => clk,
      reset => reset);

  place_1047_preds(0) <= transition_1043_symbol_out;
  place_1047_succs(0) <= transition_1044_symbol_out;
  place_1047 : place
    generic map(marking => false)
    port map(
      preds => place_1047_preds,
      succs => place_1047_succs,
      token => place_1047_token,
      clk   => clk,
      reset => reset);

  place_1048_preds(0) <= transition_1044_symbol_out;
  place_1048_succs(0) <= transition_1045_symbol_out;
  place_1048 : place
    generic map(marking => false)
    port map(
      preds => place_1048_preds,
      succs => place_1048_succs,
      token => place_1048_token,
      clk   => clk,
      reset => reset);

  place_1049_preds(0) <= transition_1045_symbol_out;
  place_1049_succs(0) <= transition_1046_symbol_out;
  place_1049 : place
    generic map(marking => false)
    port map(
      preds => place_1049_preds,
      succs => place_1049_succs,
      token => place_1049_token,
      clk   => clk,
      reset => reset);

  place_1050_preds(0) <= transition_1052_symbol_out;
  place_1050_succs(0) <= transition_1051_symbol_out;
  place_1050 : place
    generic map(marking => false)
    port map(
      preds => place_1050_preds,
      succs => place_1050_succs,
      token => place_1050_token,
      clk   => clk,
      reset => reset);

  place_1053_preds(0) <= transition_1055_symbol_out;
  place_1053_succs(0) <= transition_1054_symbol_out;
  place_1053 : place
    generic map(marking => false)
    port map(
      preds => place_1053_preds,
      succs => place_1053_succs,
      token => place_1053_token,
      clk   => clk,
      reset => reset);

  place_1060_preds(0) <= transition_1056_symbol_out;
  place_1060_succs(0) <= transition_1057_symbol_out;
  place_1060 : place
    generic map(marking => false)
    port map(
      preds => place_1060_preds,
      succs => place_1060_succs,
      token => place_1060_token,
      clk   => clk,
      reset => reset);

  place_1061_preds(0) <= transition_1057_symbol_out;
  place_1061_succs(0) <= transition_1058_symbol_out;
  place_1061 : place
    generic map(marking => false)
    port map(
      preds => place_1061_preds,
      succs => place_1061_succs,
      token => place_1061_token,
      clk   => clk,
      reset => reset);

  place_1062_preds(0) <= transition_1058_symbol_out;
  place_1062_succs(0) <= transition_1059_symbol_out;
  place_1062 : place
    generic map(marking => false)
    port map(
      preds => place_1062_preds,
      succs => place_1062_succs,
      token => place_1062_token,
      clk   => clk,
      reset => reset);

  place_1067_preds(0) <= transition_1063_symbol_out;
  place_1067_succs(0) <= transition_1064_symbol_out;
  place_1067 : place
    generic map(marking => false)
    port map(
      preds => place_1067_preds,
      succs => place_1067_succs,
      token => place_1067_token,
      clk   => clk,
      reset => reset);

  place_1068_preds(0) <= transition_1064_symbol_out;
  place_1068_succs(0) <= transition_1065_symbol_out;
  place_1068 : place
    generic map(marking => false)
    port map(
      preds => place_1068_preds,
      succs => place_1068_succs,
      token => place_1068_token,
      clk   => clk,
      reset => reset);

  place_1069_preds(0) <= transition_1065_symbol_out;
  place_1069_succs(0) <= transition_1066_symbol_out;
  place_1069 : place
    generic map(marking => false)
    port map(
      preds => place_1069_preds,
      succs => place_1069_succs,
      token => place_1069_token,
      clk   => clk,
      reset => reset);

  place_1075_preds(0) <= transition_1071_symbol_out;
  place_1075_succs(0) <= transition_1072_symbol_out;
  place_1075 : place
    generic map(marking => false)
    port map(
      preds => place_1075_preds,
      succs => place_1075_succs,
      token => place_1075_token,
      clk   => clk,
      reset => reset);

  place_1076_preds(0) <= transition_1072_symbol_out;
  place_1076_succs(0) <= transition_1073_symbol_out;
  place_1076 : place
    generic map(marking => false)
    port map(
      preds => place_1076_preds,
      succs => place_1076_succs,
      token => place_1076_token,
      clk   => clk,
      reset => reset);

  place_1077_preds(0) <= transition_1073_symbol_out;
  place_1077_succs(0) <= transition_1074_symbol_out;
  place_1077 : place
    generic map(marking => false)
    port map(
      preds => place_1077_preds,
      succs => place_1077_succs,
      token => place_1077_token,
      clk   => clk,
      reset => reset);

  place_1079_preds(0) <= transition_1081_symbol_out;
  place_1079_succs(0) <= transition_1080_symbol_out;
  place_1079 : place
    generic map(marking => false)
    port map(
      preds => place_1079_preds,
      succs => place_1079_succs,
      token => place_1079_token,
      clk   => clk,
      reset => reset);

  place_1082_preds(0) <= transition_152_symbol_out;
  place_1082_succs(0) <= transition_163_symbol_out;
  place_1082 : place
    generic map(marking => false)
    port map(
      preds => place_1082_preds,
      succs => place_1082_succs,
      token => place_1082_token,
      clk   => clk,
      reset => reset);

  place_1083_preds(0) <= transition_4_symbol_out;
  place_1083_succs(0) <= transition_149_symbol_out;
  place_1083 : place
    generic map(marking => false)
    port map(
      preds => place_1083_preds,
      succs => place_1083_succs,
      token => place_1083_token,
      clk   => clk,
      reset => reset);

  place_1084_preds(0) <= transition_163_symbol_out;
  place_1084_succs(0) <= transition_156_symbol_out;
  place_1084 : place
    generic map(marking => false)
    port map(
      preds => place_1084_preds,
      succs => place_1084_succs,
      token => place_1084_token,
      clk   => clk,
      reset => reset);

  place_1085_preds(0) <= transition_159_symbol_out;
  place_1085_succs(0) <= transition_164_symbol_out;
  place_1085 : place
    generic map(marking => false)
    port map(
      preds => place_1085_preds,
      succs => place_1085_succs,
      token => place_1085_token,
      clk   => clk,
      reset => reset);

  place_1086_preds(0) <= transition_168_symbol_out;
  place_1086_succs(0) <= transition_167_symbol_out;
  place_1086 : place
    generic map(marking => false)
    port map(
      preds => place_1086_preds,
      succs => place_1086_succs,
      token => place_1086_token,
      clk   => clk,
      reset => reset);

  place_1087_preds(0) <= transition_166_symbol_out;
  place_1087_succs(0) <= transition_216_symbol_out;
  place_1087 : place
    generic map(marking => false)
    port map(
      preds => place_1087_preds,
      succs => place_1087_succs,
      token => place_1087_token,
      clk   => clk,
      reset => reset);

  place_1088_preds(0) <= transition_7_symbol_out;
  place_1088_succs(0) <= transition_22_symbol_out;
  place_1088 : place
    generic map(marking => false)
    port map(
      preds => place_1088_preds,
      succs => place_1088_succs,
      token => place_1088_token,
      clk   => clk,
      reset => reset);

  place_1089_preds(0) <= transition_164_symbol_out;
  place_1089_succs(0) <= transition_168_symbol_out;
  place_1089 : place
    generic map(marking => false)
    port map(
      preds => place_1089_preds,
      succs => place_1089_succs,
      token => place_1089_token,
      clk   => clk,
      reset => reset);

  place_1090_preds(0) <= transition_4_symbol_out;
  place_1090_succs(0) <= transition_168_symbol_out;
  place_1090 : place
    generic map(marking => false)
    port map(
      preds => place_1090_preds,
      succs => place_1090_succs,
      token => place_1090_token,
      clk   => clk,
      reset => reset);

  place_1091_preds(0) <= transition_172_symbol_out;
  place_1091_succs(0) <= transition_190_symbol_out;
  place_1091 : place
    generic map(marking => false)
    port map(
      preds => place_1091_preds,
      succs => place_1091_succs,
      token => place_1091_token,
      clk   => clk,
      reset => reset);

  place_1092_preds(0) <= transition_4_symbol_out;
  place_1092_succs(0) <= transition_169_symbol_out;
  place_1092 : place
    generic map(marking => false)
    port map(
      preds => place_1092_preds,
      succs => place_1092_succs,
      token => place_1092_token,
      clk   => clk,
      reset => reset);

  place_1093_preds(0) <= transition_179_symbol_out;
  place_1093_succs(0) <= transition_190_symbol_out;
  place_1093 : place
    generic map(marking => false)
    port map(
      preds => place_1093_preds,
      succs => place_1093_succs,
      token => place_1093_token,
      clk   => clk,
      reset => reset);

  place_1094_preds(0) <= transition_8_symbol_out;
  place_1094_succs(0) <= transition_23_symbol_out;
  place_1094 : place
    generic map(marking => false)
    port map(
      preds => place_1094_preds,
      succs => place_1094_succs,
      token => place_1094_token,
      clk   => clk,
      reset => reset);

  place_1095_preds(0) <= transition_4_symbol_out;
  place_1095_succs(0) <= transition_176_symbol_out;
  place_1095 : place
    generic map(marking => false)
    port map(
      preds => place_1095_preds,
      succs => place_1095_succs,
      token => place_1095_token,
      clk   => clk,
      reset => reset);

  place_1096_preds(0) <= transition_190_symbol_out;
  place_1096_succs(0) <= transition_183_symbol_out;
  place_1096 : place
    generic map(marking => false)
    port map(
      preds => place_1096_preds,
      succs => place_1096_succs,
      token => place_1096_token,
      clk   => clk,
      reset => reset);

  place_1097_preds(0) <= transition_186_symbol_out;
  place_1097_succs(0) <= transition_191_symbol_out;
  place_1097 : place
    generic map(marking => false)
    port map(
      preds => place_1097_preds,
      succs => place_1097_succs,
      token => place_1097_token,
      clk   => clk,
      reset => reset);

  place_1098_preds(0) <= transition_194_symbol_out;
  place_1098_succs(0) <= transition_212_symbol_out;
  place_1098 : place
    generic map(marking => false)
    port map(
      preds => place_1098_preds,
      succs => place_1098_succs,
      token => place_1098_token,
      clk   => clk,
      reset => reset);

  place_1099_preds(0) <= transition_201_symbol_out;
  place_1099_succs(0) <= transition_212_symbol_out;
  place_1099 : place
    generic map(marking => false)
    port map(
      preds => place_1099_preds,
      succs => place_1099_succs,
      token => place_1099_token,
      clk   => clk,
      reset => reset);

  place_1100_preds(0) <= transition_164_symbol_out;
  place_1100_succs(0) <= transition_198_symbol_out;
  place_1100 : place
    generic map(marking => false)
    port map(
      preds => place_1100_preds,
      succs => place_1100_succs,
      token => place_1100_token,
      clk   => clk,
      reset => reset);

  place_1101_preds(0) <= transition_212_symbol_out;
  place_1101_succs(0) <= transition_205_symbol_out;
  place_1101 : place
    generic map(marking => false)
    port map(
      preds => place_1101_preds,
      succs => place_1101_succs,
      token => place_1101_token,
      clk   => clk,
      reset => reset);

  place_1102_preds(0) <= transition_208_symbol_out;
  place_1102_succs(0) <= transition_216_symbol_out;
  place_1102 : place
    generic map(marking => false)
    port map(
      preds => place_1102_preds,
      succs => place_1102_succs,
      token => place_1102_token,
      clk   => clk,
      reset => reset);

  place_1103_preds(0) <= transition_22_symbol_out;
  place_1103_succs(0) <= transition_26_symbol_out;
  place_1103 : place
    generic map(marking => false)
    port map(
      preds => place_1103_preds,
      succs => place_1103_succs,
      token => place_1103_token,
      clk   => clk,
      reset => reset);

  place_1104_preds(0) <= transition_216_symbol_out;
  place_1104_succs(0) <= transition_215_symbol_out;
  place_1104 : place
    generic map(marking => false)
    port map(
      preds => place_1104_preds,
      succs => place_1104_succs,
      token => place_1104_token,
      clk   => clk,
      reset => reset);

  place_1105_preds(0) <= transition_214_symbol_out;
  place_1105_succs(0) <= transition_5_symbol_out;
  place_1105 : place
    generic map(marking => false)
    port map(
      preds => place_1105_preds,
      succs => place_1105_succs,
      token => place_1105_token,
      clk   => clk,
      reset => reset);

  place_1106_preds(0) <= transition_220_symbol_out;
  place_1106_succs(0) <= transition_224_symbol_out;
  place_1106 : place
    generic map(marking => false)
    port map(
      preds => place_1106_preds,
      succs => place_1106_succs,
      token => place_1106_token,
      clk   => clk,
      reset => reset);

  place_1107_preds(0) <= transition_4_symbol_out;
  place_1107_succs(0) <= transition_217_symbol_out;
  place_1107 : place
    generic map(marking => false)
    port map(
      preds => place_1107_preds,
      succs => place_1107_succs,
      token => place_1107_token,
      clk   => clk,
      reset => reset);

  place_1108_preds(0) <= transition_25_symbol_out;
  place_1108_succs(0) <= transition_3_symbol_out;
  place_1108 : place
    generic map(marking => false)
    port map(
      preds => place_1108_preds,
      succs => place_1108_succs,
      token => place_1108_token,
      clk   => clk,
      reset => reset);

  place_1109_preds(0) <= transition_227_symbol_out;
  place_1109_succs(0) <= transition_5_symbol_out;
  place_1109 : place
    generic map(marking => false)
    port map(
      preds => place_1109_preds,
      succs => place_1109_succs,
      token => place_1109_token,
      clk   => clk,
      reset => reset);

  place_1110_preds(0) <= transition_14_symbol_out;
  place_1110_succs(0) <= transition_231_symbol_out;
  place_1110 : place
    generic map(marking => false)
    port map(
      preds => place_1110_preds,
      succs => place_1110_succs,
      token => place_1110_token,
      clk   => clk,
      reset => reset);

  place_1111_preds(0) <= transition_15_symbol_out;
  place_1111_succs(0) <= transition_17_symbol_out;
  place_1111 : place
    generic map(marking => false)
    port map(
      preds => place_1111_preds,
      succs => place_1111_succs,
      token => place_1111_token,
      clk   => clk,
      reset => reset);

  place_1112_preds(0) <= transition_23_symbol_out;
  place_1112_succs(0) <= transition_234_symbol_out;
  place_1112 : place
    generic map(marking => false)
    port map(
      preds => place_1112_preds,
      succs => place_1112_succs,
      token => place_1112_token,
      clk   => clk,
      reset => reset);

  place_1113_preds(0) <= transition_233_symbol_out;
  place_1113_succs(0) <= transition_10_symbol_out;
  place_1113 : place
    generic map(marking => false)
    port map(
      preds => place_1113_preds,
      succs => place_1113_succs,
      token => place_1113_token,
      clk   => clk,
      reset => reset);

  place_1114_preds(0) <= transition_231_symbol_out;
  place_1114_succs(0) <= transition_235_symbol_out;
  place_1114 : place
    generic map(marking => false)
    port map(
      preds => place_1114_preds,
      succs => place_1114_succs,
      token => place_1114_token,
      clk   => clk,
      reset => reset);

  place_1115_preds(0) <= transition_23_symbol_out;
  place_1115_succs(0) <= transition_238_symbol_out;
  place_1115 : place
    generic map(marking => false)
    port map(
      preds => place_1115_preds,
      succs => place_1115_succs,
      token => place_1115_token,
      clk   => clk,
      reset => reset);

  place_1116_preds(0) <= transition_237_symbol_out;
  place_1116_succs(0) <= transition_10_symbol_out;
  place_1116 : place
    generic map(marking => false)
    port map(
      preds => place_1116_preds,
      succs => place_1116_succs,
      token => place_1116_token,
      clk   => clk,
      reset => reset);

  place_1117_preds(0) <= transition_231_symbol_out;
  place_1117_succs(0) <= transition_239_symbol_out;
  place_1117 : place
    generic map(marking => false)
    port map(
      preds => place_1117_preds,
      succs => place_1117_succs,
      token => place_1117_token,
      clk   => clk,
      reset => reset);

  place_1118_preds(0) <= transition_243_symbol_out;
  place_1118_succs(0) <= transition_261_symbol_out;
  place_1118 : place
    generic map(marking => false)
    port map(
      preds => place_1118_preds,
      succs => place_1118_succs,
      token => place_1118_token,
      clk   => clk,
      reset => reset);

  place_1119_preds(0) <= transition_21_symbol_out;
  place_1119_succs(0) <= transition_27_symbol_out;
  place_1119 : place
    generic map(marking => false)
    port map(
      preds => place_1119_preds,
      succs => place_1119_succs,
      token => place_1119_token,
      clk   => clk,
      reset => reset);

  place_1120_preds(0) <= transition_11_symbol_out;
  place_1120_succs(0) <= transition_240_symbol_out;
  place_1120 : place
    generic map(marking => false)
    port map(
      preds => place_1120_preds,
      succs => place_1120_succs,
      token => place_1120_token,
      clk   => clk,
      reset => reset);

  place_1121_preds(0) <= transition_250_symbol_out;
  place_1121_succs(0) <= transition_261_symbol_out;
  place_1121 : place
    generic map(marking => false)
    port map(
      preds => place_1121_preds,
      succs => place_1121_succs,
      token => place_1121_token,
      clk   => clk,
      reset => reset);

  place_1122_preds(0) <= transition_11_symbol_out;
  place_1122_succs(0) <= transition_247_symbol_out;
  place_1122 : place
    generic map(marking => false)
    port map(
      preds => place_1122_preds,
      succs => place_1122_succs,
      token => place_1122_token,
      clk   => clk,
      reset => reset);

  place_1123_preds(0) <= transition_261_symbol_out;
  place_1123_succs(0) <= transition_254_symbol_out;
  place_1123 : place
    generic map(marking => false)
    port map(
      preds => place_1123_preds,
      succs => place_1123_succs,
      token => place_1123_token,
      clk   => clk,
      reset => reset);

  place_1124_preds(0) <= transition_257_symbol_out;
  place_1124_succs(0) <= transition_276_symbol_out;
  place_1124 : place
    generic map(marking => false)
    port map(
      preds => place_1124_preds,
      succs => place_1124_succs,
      token => place_1124_token,
      clk   => clk,
      reset => reset);

  place_1125_preds(0) <= transition_265_symbol_out;
  place_1125_succs(0) <= transition_276_symbol_out;
  place_1125 : place
    generic map(marking => false)
    port map(
      preds => place_1125_preds,
      succs => place_1125_succs,
      token => place_1125_token,
      clk   => clk,
      reset => reset);

  place_1126_preds(0) <= transition_11_symbol_out;
  place_1126_succs(0) <= transition_262_symbol_out;
  place_1126 : place
    generic map(marking => false)
    port map(
      preds => place_1126_preds,
      succs => place_1126_succs,
      token => place_1126_token,
      clk   => clk,
      reset => reset);

  place_1127_preds(0) <= transition_276_symbol_out;
  place_1127_succs(0) <= transition_269_symbol_out;
  place_1127 : place
    generic map(marking => false)
    port map(
      preds => place_1127_preds,
      succs => place_1127_succs,
      token => place_1127_token,
      clk   => clk,
      reset => reset);

  place_1128_preds(0) <= transition_272_symbol_out;
  place_1128_succs(0) <= transition_277_symbol_out;
  place_1128 : place
    generic map(marking => false)
    port map(
      preds => place_1128_preds,
      succs => place_1128_succs,
      token => place_1128_token,
      clk   => clk,
      reset => reset);

  place_1129_preds(0) <= transition_22_symbol_out;
  place_1129_succs(0) <= transition_30_symbol_out;
  place_1129 : place
    generic map(marking => false)
    port map(
      preds => place_1129_preds,
      succs => place_1129_succs,
      token => place_1129_token,
      clk   => clk,
      reset => reset);

  place_1130_preds(0) <= transition_280_symbol_out;
  place_1130_succs(0) <= transition_383_symbol_out;
  place_1130 : place
    generic map(marking => false)
    port map(
      preds => place_1130_preds,
      succs => place_1130_succs,
      token => place_1130_token,
      clk   => clk,
      reset => reset);

  place_1131_preds(0) <= transition_287_symbol_out;
  place_1131_succs(0) <= transition_305_symbol_out;
  place_1131 : place
    generic map(marking => false)
    port map(
      preds => place_1131_preds,
      succs => place_1131_succs,
      token => place_1131_token,
      clk   => clk,
      reset => reset);

  place_1132_preds(0) <= transition_3_symbol_out;
  place_1132_succs(0) <= transition_4_symbol_out;
  place_1132 : place
    generic map(marking => false)
    port map(
      preds => place_1132_preds,
      succs => place_1132_succs,
      token => place_1132_token,
      clk   => clk,
      reset => reset);

  place_1133_preds(0) <= transition_29_symbol_out;
  place_1133_succs(0) <= transition_3_symbol_out;
  place_1133 : place
    generic map(marking => false)
    port map(
      preds => place_1133_preds,
      succs => place_1133_succs,
      token => place_1133_token,
      clk   => clk,
      reset => reset);

  place_1134_preds(0) <= transition_11_symbol_out;
  place_1134_succs(0) <= transition_284_symbol_out;
  place_1134 : place
    generic map(marking => false)
    port map(
      preds => place_1134_preds,
      succs => place_1134_succs,
      token => place_1134_token,
      clk   => clk,
      reset => reset);

  place_1135_preds(0) <= transition_294_symbol_out;
  place_1135_succs(0) <= transition_305_symbol_out;
  place_1135 : place
    generic map(marking => false)
    port map(
      preds => place_1135_preds,
      succs => place_1135_succs,
      token => place_1135_token,
      clk   => clk,
      reset => reset);

  place_1136_preds(0) <= transition_11_symbol_out;
  place_1136_succs(0) <= transition_291_symbol_out;
  place_1136 : place
    generic map(marking => false)
    port map(
      preds => place_1136_preds,
      succs => place_1136_succs,
      token => place_1136_token,
      clk   => clk,
      reset => reset);

  place_1137_preds(0) <= transition_305_symbol_out;
  place_1137_succs(0) <= transition_298_symbol_out;
  place_1137 : place
    generic map(marking => false)
    port map(
      preds => place_1137_preds,
      succs => place_1137_succs,
      token => place_1137_token,
      clk   => clk,
      reset => reset);

  place_1138_preds(0) <= transition_301_symbol_out;
  place_1138_succs(0) <= transition_320_symbol_out;
  place_1138 : place
    generic map(marking => false)
    port map(
      preds => place_1138_preds,
      succs => place_1138_succs,
      token => place_1138_token,
      clk   => clk,
      reset => reset);

  place_1139_preds(0) <= transition_309_symbol_out;
  place_1139_succs(0) <= transition_320_symbol_out;
  place_1139 : place
    generic map(marking => false)
    port map(
      preds => place_1139_preds,
      succs => place_1139_succs,
      token => place_1139_token,
      clk   => clk,
      reset => reset);

  place_1140_preds(0) <= transition_11_symbol_out;
  place_1140_succs(0) <= transition_306_symbol_out;
  place_1140 : place
    generic map(marking => false)
    port map(
      preds => place_1140_preds,
      succs => place_1140_succs,
      token => place_1140_token,
      clk   => clk,
      reset => reset);

  place_1141_preds(0) <= transition_320_symbol_out;
  place_1141_succs(0) <= transition_313_symbol_out;
  place_1141 : place
    generic map(marking => false)
    port map(
      preds => place_1141_preds,
      succs => place_1141_succs,
      token => place_1141_token,
      clk   => clk,
      reset => reset);

  place_1142_preds(0) <= transition_316_symbol_out;
  place_1142_succs(0) <= transition_321_symbol_out;
  place_1142 : place
    generic map(marking => false)
    port map(
      preds => place_1142_preds,
      succs => place_1142_succs,
      token => place_1142_token,
      clk   => clk,
      reset => reset);

  place_1143_preds(0) <= transition_21_symbol_out;
  place_1143_succs(0) <= transition_31_symbol_out;
  place_1143 : place
    generic map(marking => false)
    port map(
      preds => place_1143_preds,
      succs => place_1143_succs,
      token => place_1143_token,
      clk   => clk,
      reset => reset);

  place_1144_preds(0) <= transition_324_symbol_out;
  place_1144_succs(0) <= transition_438_symbol_out;
  place_1144 : place
    generic map(marking => false)
    port map(
      preds => place_1144_preds,
      succs => place_1144_succs,
      token => place_1144_token,
      clk   => clk,
      reset => reset);

  place_1145_preds(0) <= transition_331_symbol_out;
  place_1145_succs(0) <= transition_349_symbol_out;
  place_1145 : place
    generic map(marking => false)
    port map(
      preds => place_1145_preds,
      succs => place_1145_succs,
      token => place_1145_token,
      clk   => clk,
      reset => reset);

  place_1146_preds(0) <= transition_11_symbol_out;
  place_1146_succs(0) <= transition_328_symbol_out;
  place_1146 : place
    generic map(marking => false)
    port map(
      preds => place_1146_preds,
      succs => place_1146_succs,
      token => place_1146_token,
      clk   => clk,
      reset => reset);

  place_1147_preds(0) <= transition_338_symbol_out;
  place_1147_succs(0) <= transition_349_symbol_out;
  place_1147 : place
    generic map(marking => false)
    port map(
      preds => place_1147_preds,
      succs => place_1147_succs,
      token => place_1147_token,
      clk   => clk,
      reset => reset);

  place_1148_preds(0) <= transition_11_symbol_out;
  place_1148_succs(0) <= transition_335_symbol_out;
  place_1148 : place
    generic map(marking => false)
    port map(
      preds => place_1148_preds,
      succs => place_1148_succs,
      token => place_1148_token,
      clk   => clk,
      reset => reset);

  place_1149_preds(0) <= transition_349_symbol_out;
  place_1149_succs(0) <= transition_342_symbol_out;
  place_1149 : place
    generic map(marking => false)
    port map(
      preds => place_1149_preds,
      succs => place_1149_succs,
      token => place_1149_token,
      clk   => clk,
      reset => reset);

  place_1150_preds(0) <= transition_345_symbol_out;
  place_1150_succs(0) <= transition_350_symbol_out;
  place_1150 : place
    generic map(marking => false)
    port map(
      preds => place_1150_preds,
      succs => place_1150_succs,
      token => place_1150_token,
      clk   => clk,
      reset => reset);

  place_1151_preds(0) <= transition_353_symbol_out;
  place_1151_succs(0) <= transition_371_symbol_out;
  place_1151 : place
    generic map(marking => false)
    port map(
      preds => place_1151_preds,
      succs => place_1151_succs,
      token => place_1151_token,
      clk   => clk,
      reset => reset);

  place_1152_preds(0) <= transition_35_symbol_out;
  place_1152_succs(0) <= transition_53_symbol_out;
  place_1152 : place
    generic map(marking => false)
    port map(
      preds => place_1152_preds,
      succs => place_1152_succs,
      token => place_1152_token,
      clk   => clk,
      reset => reset);

  place_1153_preds(0) <= transition_360_symbol_out;
  place_1153_succs(0) <= transition_371_symbol_out;
  place_1153 : place
    generic map(marking => false)
    port map(
      preds => place_1153_preds,
      succs => place_1153_succs,
      token => place_1153_token,
      clk   => clk,
      reset => reset);

  place_1154_preds(0) <= transition_11_symbol_out;
  place_1154_succs(0) <= transition_357_symbol_out;
  place_1154 : place
    generic map(marking => false)
    port map(
      preds => place_1154_preds,
      succs => place_1154_succs,
      token => place_1154_token,
      clk   => clk,
      reset => reset);

  place_1155_preds(0) <= transition_371_symbol_out;
  place_1155_succs(0) <= transition_364_symbol_out;
  place_1155 : place
    generic map(marking => false)
    port map(
      preds => place_1155_preds,
      succs => place_1155_succs,
      token => place_1155_token,
      clk   => clk,
      reset => reset);

  place_1156_preds(0) <= transition_367_symbol_out;
  place_1156_succs(0) <= transition_372_symbol_out;
  place_1156 : place
    generic map(marking => false)
    port map(
      preds => place_1156_preds,
      succs => place_1156_succs,
      token => place_1156_token,
      clk   => clk,
      reset => reset);

  place_1157_preds(0) <= transition_376_symbol_out;
  place_1157_succs(0) <= transition_383_symbol_out;
  place_1157 : place
    generic map(marking => false)
    port map(
      preds => place_1157_preds,
      succs => place_1157_succs,
      token => place_1157_token,
      clk   => clk,
      reset => reset);

  place_1158_preds(0) <= transition_372_symbol_out;
  place_1158_succs(0) <= transition_373_symbol_out;
  place_1158 : place
    generic map(marking => false)
    port map(
      preds => place_1158_preds,
      succs => place_1158_succs,
      token => place_1158_token,
      clk   => clk,
      reset => reset);

  place_1159_preds(0) <= transition_383_symbol_out;
  place_1159_succs(0) <= transition_382_symbol_out;
  place_1159 : place
    generic map(marking => false)
    port map(
      preds => place_1159_preds,
      succs => place_1159_succs,
      token => place_1159_token,
      clk   => clk,
      reset => reset);

  place_1160_preds(0) <= transition_381_symbol_out;
  place_1160_succs(0) <= transition_438_symbol_out;
  place_1160 : place
    generic map(marking => false)
    port map(
      preds => place_1160_preds,
      succs => place_1160_succs,
      token => place_1160_token,
      clk   => clk,
      reset => reset);

  place_1161_preds(0) <= transition_11_symbol_out;
  place_1161_succs(0) <= transition_383_symbol_out;
  place_1161 : place
    generic map(marking => false)
    port map(
      preds => place_1161_preds,
      succs => place_1161_succs,
      token => place_1161_token,
      clk   => clk,
      reset => reset);

  place_1162_preds(0) <= transition_387_symbol_out;
  place_1162_succs(0) <= transition_405_symbol_out;
  place_1162 : place
    generic map(marking => false)
    port map(
      preds => place_1162_preds,
      succs => place_1162_succs,
      token => place_1162_token,
      clk   => clk,
      reset => reset);

  place_1163_preds(0) <= transition_11_symbol_out;
  place_1163_succs(0) <= transition_384_symbol_out;
  place_1163 : place
    generic map(marking => false)
    port map(
      preds => place_1163_preds,
      succs => place_1163_succs,
      token => place_1163_token,
      clk   => clk,
      reset => reset);

  place_1164_preds(0) <= transition_394_symbol_out;
  place_1164_succs(0) <= transition_405_symbol_out;
  place_1164 : place
    generic map(marking => false)
    port map(
      preds => place_1164_preds,
      succs => place_1164_succs,
      token => place_1164_token,
      clk   => clk,
      reset => reset);

  place_1165_preds(0) <= transition_11_symbol_out;
  place_1165_succs(0) <= transition_391_symbol_out;
  place_1165 : place
    generic map(marking => false)
    port map(
      preds => place_1165_preds,
      succs => place_1165_succs,
      token => place_1165_token,
      clk   => clk,
      reset => reset);

  place_1166_preds(0) <= transition_405_symbol_out;
  place_1166_succs(0) <= transition_398_symbol_out;
  place_1166 : place
    generic map(marking => false)
    port map(
      preds => place_1166_preds,
      succs => place_1166_succs,
      token => place_1166_token,
      clk   => clk,
      reset => reset);

  place_1167_preds(0) <= transition_401_symbol_out;
  place_1167_succs(0) <= transition_406_symbol_out;
  place_1167 : place
    generic map(marking => false)
    port map(
      preds => place_1167_preds,
      succs => place_1167_succs,
      token => place_1167_token,
      clk   => clk,
      reset => reset);

  place_1168_preds(0) <= transition_4_symbol_out;
  place_1168_succs(0) <= transition_32_symbol_out;
  place_1168 : place
    generic map(marking => false)
    port map(
      preds => place_1168_preds,
      succs => place_1168_succs,
      token => place_1168_token,
      clk   => clk,
      reset => reset);

  place_1169_preds(0) <= transition_409_symbol_out;
  place_1169_succs(0) <= transition_427_symbol_out;
  place_1169 : place
    generic map(marking => false)
    port map(
      preds => place_1169_preds,
      succs => place_1169_succs,
      token => place_1169_token,
      clk   => clk,
      reset => reset);

  place_1170_preds(0) <= transition_416_symbol_out;
  place_1170_succs(0) <= transition_427_symbol_out;
  place_1170 : place
    generic map(marking => false)
    port map(
      preds => place_1170_preds,
      succs => place_1170_succs,
      token => place_1170_token,
      clk   => clk,
      reset => reset);

  place_1171_preds(0) <= transition_372_symbol_out;
  place_1171_succs(0) <= transition_413_symbol_out;
  place_1171 : place
    generic map(marking => false)
    port map(
      preds => place_1171_preds,
      succs => place_1171_succs,
      token => place_1171_token,
      clk   => clk,
      reset => reset);

  place_1172_preds(0) <= transition_427_symbol_out;
  place_1172_succs(0) <= transition_420_symbol_out;
  place_1172 : place
    generic map(marking => false)
    port map(
      preds => place_1172_preds,
      succs => place_1172_succs,
      token => place_1172_token,
      clk   => clk,
      reset => reset);

  place_1173_preds(0) <= transition_423_symbol_out;
  place_1173_succs(0) <= transition_428_symbol_out;
  place_1173 : place
    generic map(marking => false)
    port map(
      preds => place_1173_preds,
      succs => place_1173_succs,
      token => place_1173_token,
      clk   => clk,
      reset => reset);

  place_1174_preds(0) <= transition_431_symbol_out;
  place_1174_succs(0) <= transition_438_symbol_out;
  place_1174 : place
    generic map(marking => false)
    port map(
      preds => place_1174_preds,
      succs => place_1174_succs,
      token => place_1174_token,
      clk   => clk,
      reset => reset);

  place_1175_preds(0) <= transition_438_symbol_out;
  place_1175_succs(0) <= transition_437_symbol_out;
  place_1175 : place
    generic map(marking => false)
    port map(
      preds => place_1175_preds,
      succs => place_1175_succs,
      token => place_1175_token,
      clk   => clk,
      reset => reset);

  place_1176_preds(0) <= transition_42_symbol_out;
  place_1176_succs(0) <= transition_53_symbol_out;
  place_1176 : place
    generic map(marking => false)
    port map(
      preds => place_1176_preds,
      succs => place_1176_succs,
      token => place_1176_token,
      clk   => clk,
      reset => reset);

  place_1177_preds(0) <= transition_436_symbol_out;
  place_1177_succs(0) <= transition_12_symbol_out;
  place_1177 : place
    generic map(marking => false)
    port map(
      preds => place_1177_preds,
      succs => place_1177_succs,
      token => place_1177_token,
      clk   => clk,
      reset => reset);

  place_1178_preds(0) <= transition_442_symbol_out;
  place_1178_succs(0) <= transition_446_symbol_out;
  place_1178 : place
    generic map(marking => false)
    port map(
      preds => place_1178_preds,
      succs => place_1178_succs,
      token => place_1178_token,
      clk   => clk,
      reset => reset);

  place_1179_preds(0) <= transition_11_symbol_out;
  place_1179_succs(0) <= transition_439_symbol_out;
  place_1179 : place
    generic map(marking => false)
    port map(
      preds => place_1179_preds,
      succs => place_1179_succs,
      token => place_1179_token,
      clk   => clk,
      reset => reset);

  place_1180_preds(0) <= transition_449_symbol_out;
  place_1180_succs(0) <= transition_12_symbol_out;
  place_1180 : place
    generic map(marking => false)
    port map(
      preds => place_1180_preds,
      succs => place_1180_succs,
      token => place_1180_token,
      clk   => clk,
      reset => reset);

  place_1181_preds(0) <= transition_5_symbol_out;
  place_1181_succs(0) <= transition_9_symbol_out;
  place_1181 : place
    generic map(marking => false)
    port map(
      preds => place_1181_preds,
      succs => place_1181_succs,
      token => place_1181_token,
      clk   => clk,
      reset => reset);

  place_1182_preds(0) <= transition_456_symbol_out;
  place_1182_succs(0) <= transition_474_symbol_out;
  place_1182 : place
    generic map(marking => false)
    port map(
      preds => place_1182_preds,
      succs => place_1182_succs,
      token => place_1182_token,
      clk   => clk,
      reset => reset);

  place_1183_preds(0) <= transition_17_symbol_out;
  place_1183_succs(0) <= transition_453_symbol_out;
  place_1183 : place
    generic map(marking => false)
    port map(
      preds => place_1183_preds,
      succs => place_1183_succs,
      token => place_1183_token,
      clk   => clk,
      reset => reset);

  place_1184_preds(0) <= transition_463_symbol_out;
  place_1184_succs(0) <= transition_474_symbol_out;
  place_1184 : place
    generic map(marking => false)
    port map(
      preds => place_1184_preds,
      succs => place_1184_succs,
      token => place_1184_token,
      clk   => clk,
      reset => reset);

  place_1185_preds(0) <= transition_17_symbol_out;
  place_1185_succs(0) <= transition_460_symbol_out;
  place_1185 : place
    generic map(marking => false)
    port map(
      preds => place_1185_preds,
      succs => place_1185_succs,
      token => place_1185_token,
      clk   => clk,
      reset => reset);

  place_1186_preds(0) <= transition_474_symbol_out;
  place_1186_succs(0) <= transition_467_symbol_out;
  place_1186 : place
    generic map(marking => false)
    port map(
      preds => place_1186_preds,
      succs => place_1186_succs,
      token => place_1186_token,
      clk   => clk,
      reset => reset);

  place_1187_preds(0) <= transition_470_symbol_out;
  place_1187_succs(0) <= transition_489_symbol_out;
  place_1187 : place
    generic map(marking => false)
    port map(
      preds => place_1187_preds,
      succs => place_1187_succs,
      token => place_1187_token,
      clk   => clk,
      reset => reset);

  place_1188_preds(0) <= transition_478_symbol_out;
  place_1188_succs(0) <= transition_489_symbol_out;
  place_1188 : place
    generic map(marking => false)
    port map(
      preds => place_1188_preds,
      succs => place_1188_succs,
      token => place_1188_token,
      clk   => clk,
      reset => reset);

  place_1189_preds(0) <= transition_4_symbol_out;
  place_1189_succs(0) <= transition_39_symbol_out;
  place_1189 : place
    generic map(marking => false)
    port map(
      preds => place_1189_preds,
      succs => place_1189_succs,
      token => place_1189_token,
      clk   => clk,
      reset => reset);

  place_1190_preds(0) <= transition_17_symbol_out;
  place_1190_succs(0) <= transition_475_symbol_out;
  place_1190 : place
    generic map(marking => false)
    port map(
      preds => place_1190_preds,
      succs => place_1190_succs,
      token => place_1190_token,
      clk   => clk,
      reset => reset);

  place_1191_preds(0) <= transition_489_symbol_out;
  place_1191_succs(0) <= transition_482_symbol_out;
  place_1191 : place
    generic map(marking => false)
    port map(
      preds => place_1191_preds,
      succs => place_1191_succs,
      token => place_1191_token,
      clk   => clk,
      reset => reset);

  place_1192_preds(0) <= transition_485_symbol_out;
  place_1192_succs(0) <= transition_490_symbol_out;
  place_1192 : place
    generic map(marking => false)
    port map(
      preds => place_1192_preds,
      succs => place_1192_succs,
      token => place_1192_token,
      clk   => clk,
      reset => reset);

  place_1193_preds(0) <= transition_493_symbol_out;
  place_1193_succs(0) <= transition_500_symbol_out;
  place_1193 : place
    generic map(marking => false)
    port map(
      preds => place_1193_preds,
      succs => place_1193_succs,
      token => place_1193_token,
      clk   => clk,
      reset => reset);

  place_1194_preds(0) <= transition_53_symbol_out;
  place_1194_succs(0) <= transition_46_symbol_out;
  place_1194 : place
    generic map(marking => false)
    port map(
      preds => place_1194_preds,
      succs => place_1194_succs,
      token => place_1194_token,
      clk   => clk,
      reset => reset);

  place_1195_preds(0) <= transition_500_symbol_out;
  place_1195_succs(0) <= transition_499_symbol_out;
  place_1195 : place
    generic map(marking => false)
    port map(
      preds => place_1195_preds,
      succs => place_1195_succs,
      token => place_1195_token,
      clk   => clk,
      reset => reset);

  place_1196_preds(0) <= transition_498_symbol_out;
  place_1196_succs(0) <= transition_548_symbol_out;
  place_1196 : place
    generic map(marking => false)
    port map(
      preds => place_1196_preds,
      succs => place_1196_succs,
      token => place_1196_token,
      clk   => clk,
      reset => reset);

  place_1197_preds(0) <= transition_17_symbol_out;
  place_1197_succs(0) <= transition_500_symbol_out;
  place_1197 : place
    generic map(marking => false)
    port map(
      preds => place_1197_preds,
      succs => place_1197_succs,
      token => place_1197_token,
      clk   => clk,
      reset => reset);

  place_1198_preds(0) <= transition_504_symbol_out;
  place_1198_succs(0) <= transition_522_symbol_out;
  place_1198 : place
    generic map(marking => false)
    port map(
      preds => place_1198_preds,
      succs => place_1198_succs,
      token => place_1198_token,
      clk   => clk,
      reset => reset);

  place_1199_preds(0) <= transition_17_symbol_out;
  place_1199_succs(0) <= transition_501_symbol_out;
  place_1199 : place
    generic map(marking => false)
    port map(
      preds => place_1199_preds,
      succs => place_1199_succs,
      token => place_1199_token,
      clk   => clk,
      reset => reset);

  place_1200_preds(0) <= transition_49_symbol_out;
  place_1200_succs(0) <= transition_68_symbol_out;
  place_1200 : place
    generic map(marking => false)
    port map(
      preds => place_1200_preds,
      succs => place_1200_succs,
      token => place_1200_token,
      clk   => clk,
      reset => reset);

  place_1201_preds(0) <= transition_511_symbol_out;
  place_1201_succs(0) <= transition_522_symbol_out;
  place_1201 : place
    generic map(marking => false)
    port map(
      preds => place_1201_preds,
      succs => place_1201_succs,
      token => place_1201_token,
      clk   => clk,
      reset => reset);

  place_1202_preds(0) <= transition_17_symbol_out;
  place_1202_succs(0) <= transition_508_symbol_out;
  place_1202 : place
    generic map(marking => false)
    port map(
      preds => place_1202_preds,
      succs => place_1202_succs,
      token => place_1202_token,
      clk   => clk,
      reset => reset);

  place_1203_preds(0) <= transition_522_symbol_out;
  place_1203_succs(0) <= transition_515_symbol_out;
  place_1203 : place
    generic map(marking => false)
    port map(
      preds => place_1203_preds,
      succs => place_1203_succs,
      token => place_1203_token,
      clk   => clk,
      reset => reset);

  place_1204_preds(0) <= transition_518_symbol_out;
  place_1204_succs(0) <= transition_537_symbol_out;
  place_1204 : place
    generic map(marking => false)
    port map(
      preds => place_1204_preds,
      succs => place_1204_succs,
      token => place_1204_token,
      clk   => clk,
      reset => reset);

  place_1205_preds(0) <= transition_526_symbol_out;
  place_1205_succs(0) <= transition_537_symbol_out;
  place_1205 : place
    generic map(marking => false)
    port map(
      preds => place_1205_preds,
      succs => place_1205_succs,
      token => place_1205_token,
      clk   => clk,
      reset => reset);

  place_1206_preds(0) <= transition_17_symbol_out;
  place_1206_succs(0) <= transition_523_symbol_out;
  place_1206 : place
    generic map(marking => false)
    port map(
      preds => place_1206_preds,
      succs => place_1206_succs,
      token => place_1206_token,
      clk   => clk,
      reset => reset);

  place_1207_preds(0) <= transition_537_symbol_out;
  place_1207_succs(0) <= transition_530_symbol_out;
  place_1207 : place
    generic map(marking => false)
    port map(
      preds => place_1207_preds,
      succs => place_1207_succs,
      token => place_1207_token,
      clk   => clk,
      reset => reset);

  place_1208_preds(0) <= transition_533_symbol_out;
  place_1208_succs(0) <= transition_538_symbol_out;
  place_1208 : place
    generic map(marking => false)
    port map(
      preds => place_1208_preds,
      succs => place_1208_succs,
      token => place_1208_token,
      clk   => clk,
      reset => reset);

  place_1209_preds(0) <= transition_541_symbol_out;
  place_1209_succs(0) <= transition_548_symbol_out;
  place_1209 : place
    generic map(marking => false)
    port map(
      preds => place_1209_preds,
      succs => place_1209_succs,
      token => place_1209_token,
      clk   => clk,
      reset => reset);

  place_1210_preds(0) <= transition_548_symbol_out;
  place_1210_succs(0) <= transition_547_symbol_out;
  place_1210 : place
    generic map(marking => false)
    port map(
      preds => place_1210_preds,
      succs => place_1210_succs,
      token => place_1210_token,
      clk   => clk,
      reset => reset);

  place_1211_preds(0) <= transition_546_symbol_out;
  place_1211_succs(0) <= transition_596_symbol_out;
  place_1211 : place
    generic map(marking => false)
    port map(
      preds => place_1211_preds,
      succs => place_1211_succs,
      token => place_1211_token,
      clk   => clk,
      reset => reset);

  place_1212_preds(0) <= transition_552_symbol_out;
  place_1212_succs(0) <= transition_570_symbol_out;
  place_1212 : place
    generic map(marking => false)
    port map(
      preds => place_1212_preds,
      succs => place_1212_succs,
      token => place_1212_token,
      clk   => clk,
      reset => reset);

  place_1213_preds(0) <= transition_17_symbol_out;
  place_1213_succs(0) <= transition_549_symbol_out;
  place_1213 : place
    generic map(marking => false)
    port map(
      preds => place_1213_preds,
      succs => place_1213_succs,
      token => place_1213_token,
      clk   => clk,
      reset => reset);

  place_1214_preds(0) <= transition_559_symbol_out;
  place_1214_succs(0) <= transition_570_symbol_out;
  place_1214 : place
    generic map(marking => false)
    port map(
      preds => place_1214_preds,
      succs => place_1214_succs,
      token => place_1214_token,
      clk   => clk,
      reset => reset);

  place_1215_preds(0) <= transition_17_symbol_out;
  place_1215_succs(0) <= transition_556_symbol_out;
  place_1215 : place
    generic map(marking => false)
    port map(
      preds => place_1215_preds,
      succs => place_1215_succs,
      token => place_1215_token,
      clk   => clk,
      reset => reset);

  place_1216_preds(0) <= transition_570_symbol_out;
  place_1216_succs(0) <= transition_563_symbol_out;
  place_1216 : place
    generic map(marking => false)
    port map(
      preds => place_1216_preds,
      succs => place_1216_succs,
      token => place_1216_token,
      clk   => clk,
      reset => reset);

  place_1217_preds(0) <= transition_566_symbol_out;
  place_1217_succs(0) <= transition_585_symbol_out;
  place_1217 : place
    generic map(marking => false)
    port map(
      preds => place_1217_preds,
      succs => place_1217_succs,
      token => place_1217_token,
      clk   => clk,
      reset => reset);

  place_1218_preds(0) <= transition_574_symbol_out;
  place_1218_succs(0) <= transition_585_symbol_out;
  place_1218 : place
    generic map(marking => false)
    port map(
      preds => place_1218_preds,
      succs => place_1218_succs,
      token => place_1218_token,
      clk   => clk,
      reset => reset);

  place_1219_preds(0) <= transition_17_symbol_out;
  place_1219_succs(0) <= transition_571_symbol_out;
  place_1219 : place
    generic map(marking => false)
    port map(
      preds => place_1219_preds,
      succs => place_1219_succs,
      token => place_1219_token,
      clk   => clk,
      reset => reset);

  place_1220_preds(0) <= transition_585_symbol_out;
  place_1220_succs(0) <= transition_578_symbol_out;
  place_1220 : place
    generic map(marking => false)
    port map(
      preds => place_1220_preds,
      succs => place_1220_succs,
      token => place_1220_token,
      clk   => clk,
      reset => reset);

  place_1221_preds(0) <= transition_581_symbol_out;
  place_1221_succs(0) <= transition_586_symbol_out;
  place_1221 : place
    generic map(marking => false)
    port map(
      preds => place_1221_preds,
      succs => place_1221_succs,
      token => place_1221_token,
      clk   => clk,
      reset => reset);

  place_1222_preds(0) <= transition_57_symbol_out;
  place_1222_succs(0) <= transition_68_symbol_out;
  place_1222 : place
    generic map(marking => false)
    port map(
      preds => place_1222_preds,
      succs => place_1222_succs,
      token => place_1222_token,
      clk   => clk,
      reset => reset);

  place_1223_preds(0) <= transition_589_symbol_out;
  place_1223_succs(0) <= transition_596_symbol_out;
  place_1223 : place
    generic map(marking => false)
    port map(
      preds => place_1223_preds,
      succs => place_1223_succs,
      token => place_1223_token,
      clk   => clk,
      reset => reset);

  place_1224_preds(0) <= transition_596_symbol_out;
  place_1224_succs(0) <= transition_595_symbol_out;
  place_1224 : place
    generic map(marking => false)
    port map(
      preds => place_1224_preds,
      succs => place_1224_succs,
      token => place_1224_token,
      clk   => clk,
      reset => reset);

  place_1225_preds(0) <= transition_594_symbol_out;
  place_1225_succs(0) <= transition_644_symbol_out;
  place_1225 : place
    generic map(marking => false)
    port map(
      preds => place_1225_preds,
      succs => place_1225_succs,
      token => place_1225_token,
      clk   => clk,
      reset => reset);

  place_1226_preds(0) <= transition_600_symbol_out;
  place_1226_succs(0) <= transition_618_symbol_out;
  place_1226 : place
    generic map(marking => false)
    port map(
      preds => place_1226_preds,
      succs => place_1226_succs,
      token => place_1226_token,
      clk   => clk,
      reset => reset);

  place_1227_preds(0) <= transition_10_symbol_out;
  place_1227_succs(0) <= transition_11_symbol_out;
  place_1227 : place
    generic map(marking => false)
    port map(
      preds => place_1227_preds,
      succs => place_1227_succs,
      token => place_1227_token,
      clk   => clk,
      reset => reset);

  place_1228_preds(0) <= transition_17_symbol_out;
  place_1228_succs(0) <= transition_597_symbol_out;
  place_1228 : place
    generic map(marking => false)
    port map(
      preds => place_1228_preds,
      succs => place_1228_succs,
      token => place_1228_token,
      clk   => clk,
      reset => reset);

  place_1229_preds(0) <= transition_607_symbol_out;
  place_1229_succs(0) <= transition_618_symbol_out;
  place_1229 : place
    generic map(marking => false)
    port map(
      preds => place_1229_preds,
      succs => place_1229_succs,
      token => place_1229_token,
      clk   => clk,
      reset => reset);

  place_1230_preds(0) <= transition_17_symbol_out;
  place_1230_succs(0) <= transition_604_symbol_out;
  place_1230 : place
    generic map(marking => false)
    port map(
      preds => place_1230_preds,
      succs => place_1230_succs,
      token => place_1230_token,
      clk   => clk,
      reset => reset);

  place_1231_preds(0) <= transition_618_symbol_out;
  place_1231_succs(0) <= transition_611_symbol_out;
  place_1231 : place
    generic map(marking => false)
    port map(
      preds => place_1231_preds,
      succs => place_1231_succs,
      token => place_1231_token,
      clk   => clk,
      reset => reset);

  place_1232_preds(0) <= transition_614_symbol_out;
  place_1232_succs(0) <= transition_633_symbol_out;
  place_1232 : place
    generic map(marking => false)
    port map(
      preds => place_1232_preds,
      succs => place_1232_succs,
      token => place_1232_token,
      clk   => clk,
      reset => reset);

  place_1233_preds(0) <= transition_622_symbol_out;
  place_1233_succs(0) <= transition_633_symbol_out;
  place_1233 : place
    generic map(marking => false)
    port map(
      preds => place_1233_preds,
      succs => place_1233_succs,
      token => place_1233_token,
      clk   => clk,
      reset => reset);

  place_1234_preds(0) <= transition_17_symbol_out;
  place_1234_succs(0) <= transition_619_symbol_out;
  place_1234 : place
    generic map(marking => false)
    port map(
      preds => place_1234_preds,
      succs => place_1234_succs,
      token => place_1234_token,
      clk   => clk,
      reset => reset);

  place_1235_preds(0) <= transition_633_symbol_out;
  place_1235_succs(0) <= transition_626_symbol_out;
  place_1235 : place
    generic map(marking => false)
    port map(
      preds => place_1235_preds,
      succs => place_1235_succs,
      token => place_1235_token,
      clk   => clk,
      reset => reset);

  place_1236_preds(0) <= transition_629_symbol_out;
  place_1236_succs(0) <= transition_634_symbol_out;
  place_1236 : place
    generic map(marking => false)
    port map(
      preds => place_1236_preds,
      succs => place_1236_succs,
      token => place_1236_token,
      clk   => clk,
      reset => reset);

  place_1237_preds(0) <= transition_4_symbol_out;
  place_1237_succs(0) <= transition_54_symbol_out;
  place_1237 : place
    generic map(marking => false)
    port map(
      preds => place_1237_preds,
      succs => place_1237_succs,
      token => place_1237_token,
      clk   => clk,
      reset => reset);

  place_1238_preds(0) <= transition_637_symbol_out;
  place_1238_succs(0) <= transition_644_symbol_out;
  place_1238 : place
    generic map(marking => false)
    port map(
      preds => place_1238_preds,
      succs => place_1238_succs,
      token => place_1238_token,
      clk   => clk,
      reset => reset);

  place_1239_preds(0) <= transition_644_symbol_out;
  place_1239_succs(0) <= transition_643_symbol_out;
  place_1239 : place
    generic map(marking => false)
    port map(
      preds => place_1239_preds,
      succs => place_1239_succs,
      token => place_1239_token,
      clk   => clk,
      reset => reset);

  place_1240_preds(0) <= transition_642_symbol_out;
  place_1240_succs(0) <= transition_692_symbol_out;
  place_1240 : place
    generic map(marking => false)
    port map(
      preds => place_1240_preds,
      succs => place_1240_succs,
      token => place_1240_token,
      clk   => clk,
      reset => reset);

  place_1241_preds(0) <= transition_68_symbol_out;
  place_1241_succs(0) <= transition_61_symbol_out;
  place_1241 : place
    generic map(marking => false)
    port map(
      preds => place_1241_preds,
      succs => place_1241_succs,
      token => place_1241_token,
      clk   => clk,
      reset => reset);

  place_1242_preds(0) <= transition_648_symbol_out;
  place_1242_succs(0) <= transition_666_symbol_out;
  place_1242 : place
    generic map(marking => false)
    port map(
      preds => place_1242_preds,
      succs => place_1242_succs,
      token => place_1242_token,
      clk   => clk,
      reset => reset);

  place_1243_preds(0) <= transition_17_symbol_out;
  place_1243_succs(0) <= transition_645_symbol_out;
  place_1243 : place
    generic map(marking => false)
    port map(
      preds => place_1243_preds,
      succs => place_1243_succs,
      token => place_1243_token,
      clk   => clk,
      reset => reset);

  place_1244_preds(0) <= transition_655_symbol_out;
  place_1244_succs(0) <= transition_666_symbol_out;
  place_1244 : place
    generic map(marking => false)
    port map(
      preds => place_1244_preds,
      succs => place_1244_succs,
      token => place_1244_token,
      clk   => clk,
      reset => reset);

  place_1245_preds(0) <= transition_17_symbol_out;
  place_1245_succs(0) <= transition_652_symbol_out;
  place_1245 : place
    generic map(marking => false)
    port map(
      preds => place_1245_preds,
      succs => place_1245_succs,
      token => place_1245_token,
      clk   => clk,
      reset => reset);

  place_1246_preds(0) <= transition_666_symbol_out;
  place_1246_succs(0) <= transition_659_symbol_out;
  place_1246 : place
    generic map(marking => false)
    port map(
      preds => place_1246_preds,
      succs => place_1246_succs,
      token => place_1246_token,
      clk   => clk,
      reset => reset);

  place_1247_preds(0) <= transition_662_symbol_out;
  place_1247_succs(0) <= transition_681_symbol_out;
  place_1247 : place
    generic map(marking => false)
    port map(
      preds => place_1247_preds,
      succs => place_1247_succs,
      token => place_1247_token,
      clk   => clk,
      reset => reset);

  place_1248_preds(0) <= transition_64_symbol_out;
  place_1248_succs(0) <= transition_69_symbol_out;
  place_1248 : place
    generic map(marking => false)
    port map(
      preds => place_1248_preds,
      succs => place_1248_succs,
      token => place_1248_token,
      clk   => clk,
      reset => reset);

  place_1249_preds(0) <= transition_670_symbol_out;
  place_1249_succs(0) <= transition_681_symbol_out;
  place_1249 : place
    generic map(marking => false)
    port map(
      preds => place_1249_preds,
      succs => place_1249_succs,
      token => place_1249_token,
      clk   => clk,
      reset => reset);

  place_1250_preds(0) <= transition_17_symbol_out;
  place_1250_succs(0) <= transition_667_symbol_out;
  place_1250 : place
    generic map(marking => false)
    port map(
      preds => place_1250_preds,
      succs => place_1250_succs,
      token => place_1250_token,
      clk   => clk,
      reset => reset);

  place_1251_preds(0) <= transition_681_symbol_out;
  place_1251_succs(0) <= transition_674_symbol_out;
  place_1251 : place
    generic map(marking => false)
    port map(
      preds => place_1251_preds,
      succs => place_1251_succs,
      token => place_1251_token,
      clk   => clk,
      reset => reset);

  place_1252_preds(0) <= transition_677_symbol_out;
  place_1252_succs(0) <= transition_682_symbol_out;
  place_1252 : place
    generic map(marking => false)
    port map(
      preds => place_1252_preds,
      succs => place_1252_succs,
      token => place_1252_token,
      clk   => clk,
      reset => reset);

  place_1253_preds(0) <= transition_685_symbol_out;
  place_1253_succs(0) <= transition_692_symbol_out;
  place_1253 : place
    generic map(marking => false)
    port map(
      preds => place_1253_preds,
      succs => place_1253_succs,
      token => place_1253_token,
      clk   => clk,
      reset => reset);

  place_1254_preds(0) <= transition_692_symbol_out;
  place_1254_succs(0) <= transition_691_symbol_out;
  place_1254 : place
    generic map(marking => false)
    port map(
      preds => place_1254_preds,
      succs => place_1254_succs,
      token => place_1254_token,
      clk   => clk,
      reset => reset);

  place_1255_preds(0) <= transition_690_symbol_out;
  place_1255_succs(0) <= transition_740_symbol_out;
  place_1255 : place
    generic map(marking => false)
    port map(
      preds => place_1255_preds,
      succs => place_1255_succs,
      token => place_1255_token,
      clk   => clk,
      reset => reset);

  place_1256_preds(0) <= transition_696_symbol_out;
  place_1256_succs(0) <= transition_714_symbol_out;
  place_1256 : place
    generic map(marking => false)
    port map(
      preds => place_1256_preds,
      succs => place_1256_succs,
      token => place_1256_token,
      clk   => clk,
      reset => reset);

  place_1257_preds(0) <= transition_17_symbol_out;
  place_1257_succs(0) <= transition_693_symbol_out;
  place_1257 : place
    generic map(marking => false)
    port map(
      preds => place_1257_preds,
      succs => place_1257_succs,
      token => place_1257_token,
      clk   => clk,
      reset => reset);

  place_1258_preds(0) <= transition_703_symbol_out;
  place_1258_succs(0) <= transition_714_symbol_out;
  place_1258 : place
    generic map(marking => false)
    port map(
      preds => place_1258_preds,
      succs => place_1258_succs,
      token => place_1258_token,
      clk   => clk,
      reset => reset);

  place_1259_preds(0) <= transition_17_symbol_out;
  place_1259_succs(0) <= transition_700_symbol_out;
  place_1259 : place
    generic map(marking => false)
    port map(
      preds => place_1259_preds,
      succs => place_1259_succs,
      token => place_1259_token,
      clk   => clk,
      reset => reset);

  place_1260_preds(0) <= transition_714_symbol_out;
  place_1260_succs(0) <= transition_707_symbol_out;
  place_1260 : place
    generic map(marking => false)
    port map(
      preds => place_1260_preds,
      succs => place_1260_succs,
      token => place_1260_token,
      clk   => clk,
      reset => reset);

  place_1261_preds(0) <= transition_710_symbol_out;
  place_1261_succs(0) <= transition_729_symbol_out;
  place_1261 : place
    generic map(marking => false)
    port map(
      preds => place_1261_preds,
      succs => place_1261_succs,
      token => place_1261_token,
      clk   => clk,
      reset => reset);

  place_1262_preds(0) <= transition_718_symbol_out;
  place_1262_succs(0) <= transition_729_symbol_out;
  place_1262 : place
    generic map(marking => false)
    port map(
      preds => place_1262_preds,
      succs => place_1262_succs,
      token => place_1262_token,
      clk   => clk,
      reset => reset);

  place_1263_preds(0) <= transition_17_symbol_out;
  place_1263_succs(0) <= transition_715_symbol_out;
  place_1263 : place
    generic map(marking => false)
    port map(
      preds => place_1263_preds,
      succs => place_1263_succs,
      token => place_1263_token,
      clk   => clk,
      reset => reset);

  place_1264_preds(0) <= transition_729_symbol_out;
  place_1264_succs(0) <= transition_722_symbol_out;
  place_1264 : place
    generic map(marking => false)
    port map(
      preds => place_1264_preds,
      succs => place_1264_succs,
      token => place_1264_token,
      clk   => clk,
      reset => reset);

  place_1265_preds(0) <= transition_725_symbol_out;
  place_1265_succs(0) <= transition_730_symbol_out;
  place_1265 : place
    generic map(marking => false)
    port map(
      preds => place_1265_preds,
      succs => place_1265_succs,
      token => place_1265_token,
      clk   => clk,
      reset => reset);

  place_1266_preds(0) <= transition_733_symbol_out;
  place_1266_succs(0) <= transition_740_symbol_out;
  place_1266 : place
    generic map(marking => false)
    port map(
      preds => place_1266_preds,
      succs => place_1266_succs,
      token => place_1266_token,
      clk   => clk,
      reset => reset);

  place_1267_preds(0) <= transition_740_symbol_out;
  place_1267_succs(0) <= transition_739_symbol_out;
  place_1267 : place
    generic map(marking => false)
    port map(
      preds => place_1267_preds,
      succs => place_1267_succs,
      token => place_1267_token,
      clk   => clk,
      reset => reset);

  place_1268_preds(0) <= transition_738_symbol_out;
  place_1268_succs(0) <= transition_788_symbol_out;
  place_1268 : place
    generic map(marking => false)
    port map(
      preds => place_1268_preds,
      succs => place_1268_succs,
      token => place_1268_token,
      clk   => clk,
      reset => reset);

  place_1269_preds(0) <= transition_72_symbol_out;
  place_1269_succs(0) <= transition_168_symbol_out;
  place_1269 : place
    generic map(marking => false)
    port map(
      preds => place_1269_preds,
      succs => place_1269_succs,
      token => place_1269_token,
      clk   => clk,
      reset => reset);

  place_1270_preds(0) <= transition_744_symbol_out;
  place_1270_succs(0) <= transition_762_symbol_out;
  place_1270 : place
    generic map(marking => false)
    port map(
      preds => place_1270_preds,
      succs => place_1270_succs,
      token => place_1270_token,
      clk   => clk,
      reset => reset);

  place_1271_preds(0) <= transition_17_symbol_out;
  place_1271_succs(0) <= transition_741_symbol_out;
  place_1271 : place
    generic map(marking => false)
    port map(
      preds => place_1271_preds,
      succs => place_1271_succs,
      token => place_1271_token,
      clk   => clk,
      reset => reset);

  place_1272_preds(0) <= transition_751_symbol_out;
  place_1272_succs(0) <= transition_762_symbol_out;
  place_1272 : place
    generic map(marking => false)
    port map(
      preds => place_1272_preds,
      succs => place_1272_succs,
      token => place_1272_token,
      clk   => clk,
      reset => reset);

  place_1273_preds(0) <= transition_12_symbol_out;
  place_1273_succs(0) <= transition_16_symbol_out;
  place_1273 : place
    generic map(marking => false)
    port map(
      preds => place_1273_preds,
      succs => place_1273_succs,
      token => place_1273_token,
      clk   => clk,
      reset => reset);

  place_1274_preds(0) <= transition_17_symbol_out;
  place_1274_succs(0) <= transition_748_symbol_out;
  place_1274 : place
    generic map(marking => false)
    port map(
      preds => place_1274_preds,
      succs => place_1274_succs,
      token => place_1274_token,
      clk   => clk,
      reset => reset);

  place_1275_preds(0) <= transition_762_symbol_out;
  place_1275_succs(0) <= transition_755_symbol_out;
  place_1275 : place
    generic map(marking => false)
    port map(
      preds => place_1275_preds,
      succs => place_1275_succs,
      token => place_1275_token,
      clk   => clk,
      reset => reset);

  place_1276_preds(0) <= transition_758_symbol_out;
  place_1276_succs(0) <= transition_777_symbol_out;
  place_1276 : place
    generic map(marking => false)
    port map(
      preds => place_1276_preds,
      succs => place_1276_succs,
      token => place_1276_token,
      clk   => clk,
      reset => reset);

  place_1277_preds(0) <= transition_766_symbol_out;
  place_1277_succs(0) <= transition_777_symbol_out;
  place_1277 : place
    generic map(marking => false)
    port map(
      preds => place_1277_preds,
      succs => place_1277_succs,
      token => place_1277_token,
      clk   => clk,
      reset => reset);

  place_1278_preds(0) <= transition_17_symbol_out;
  place_1278_succs(0) <= transition_763_symbol_out;
  place_1278 : place
    generic map(marking => false)
    port map(
      preds => place_1278_preds,
      succs => place_1278_succs,
      token => place_1278_token,
      clk   => clk,
      reset => reset);

  place_1279_preds(0) <= transition_777_symbol_out;
  place_1279_succs(0) <= transition_770_symbol_out;
  place_1279 : place
    generic map(marking => false)
    port map(
      preds => place_1279_preds,
      succs => place_1279_succs,
      token => place_1279_token,
      clk   => clk,
      reset => reset);

  place_1280_preds(0) <= transition_773_symbol_out;
  place_1280_succs(0) <= transition_778_symbol_out;
  place_1280 : place
    generic map(marking => false)
    port map(
      preds => place_1280_preds,
      succs => place_1280_succs,
      token => place_1280_token,
      clk   => clk,
      reset => reset);

  place_1281_preds(0) <= transition_781_symbol_out;
  place_1281_succs(0) <= transition_788_symbol_out;
  place_1281 : place
    generic map(marking => false)
    port map(
      preds => place_1281_preds,
      succs => place_1281_succs,
      token => place_1281_token,
      clk   => clk,
      reset => reset);

  place_1282_preds(0) <= transition_788_symbol_out;
  place_1282_succs(0) <= transition_787_symbol_out;
  place_1282 : place
    generic map(marking => false)
    port map(
      preds => place_1282_preds,
      succs => place_1282_succs,
      token => place_1282_token,
      clk   => clk,
      reset => reset);

  place_1283_preds(0) <= transition_786_symbol_out;
  place_1283_succs(0) <= transition_836_symbol_out;
  place_1283 : place
    generic map(marking => false)
    port map(
      preds => place_1283_preds,
      succs => place_1283_succs,
      token => place_1283_token,
      clk   => clk,
      reset => reset);

  place_1284_preds(0) <= transition_792_symbol_out;
  place_1284_succs(0) <= transition_810_symbol_out;
  place_1284 : place
    generic map(marking => false)
    port map(
      preds => place_1284_preds,
      succs => place_1284_succs,
      token => place_1284_token,
      clk   => clk,
      reset => reset);

  place_1285_preds(0) <= transition_17_symbol_out;
  place_1285_succs(0) <= transition_789_symbol_out;
  place_1285 : place
    generic map(marking => false)
    port map(
      preds => place_1285_preds,
      succs => place_1285_succs,
      token => place_1285_token,
      clk   => clk,
      reset => reset);

  place_1286_preds(0) <= transition_79_symbol_out;
  place_1286_succs(0) <= transition_97_symbol_out;
  place_1286 : place
    generic map(marking => false)
    port map(
      preds => place_1286_preds,
      succs => place_1286_succs,
      token => place_1286_token,
      clk   => clk,
      reset => reset);

  place_1287_preds(0) <= transition_799_symbol_out;
  place_1287_succs(0) <= transition_810_symbol_out;
  place_1287 : place
    generic map(marking => false)
    port map(
      preds => place_1287_preds,
      succs => place_1287_succs,
      token => place_1287_token,
      clk   => clk,
      reset => reset);

  place_1288_preds(0) <= transition_17_symbol_out;
  place_1288_succs(0) <= transition_796_symbol_out;
  place_1288 : place
    generic map(marking => false)
    port map(
      preds => place_1288_preds,
      succs => place_1288_succs,
      token => place_1288_token,
      clk   => clk,
      reset => reset);

  place_1289_preds(0) <= transition_810_symbol_out;
  place_1289_succs(0) <= transition_803_symbol_out;
  place_1289 : place
    generic map(marking => false)
    port map(
      preds => place_1289_preds,
      succs => place_1289_succs,
      token => place_1289_token,
      clk   => clk,
      reset => reset);

  place_1290_preds(0) <= transition_806_symbol_out;
  place_1290_succs(0) <= transition_825_symbol_out;
  place_1290 : place
    generic map(marking => false)
    port map(
      preds => place_1290_preds,
      succs => place_1290_succs,
      token => place_1290_token,
      clk   => clk,
      reset => reset);

  place_1291_preds(0) <= transition_814_symbol_out;
  place_1291_succs(0) <= transition_825_symbol_out;
  place_1291 : place
    generic map(marking => false)
    port map(
      preds => place_1291_preds,
      succs => place_1291_succs,
      token => place_1291_token,
      clk   => clk,
      reset => reset);

  place_1292_preds(0) <= transition_17_symbol_out;
  place_1292_succs(0) <= transition_811_symbol_out;
  place_1292 : place
    generic map(marking => false)
    port map(
      preds => place_1292_preds,
      succs => place_1292_succs,
      token => place_1292_token,
      clk   => clk,
      reset => reset);

  place_1293_preds(0) <= transition_825_symbol_out;
  place_1293_succs(0) <= transition_818_symbol_out;
  place_1293 : place
    generic map(marking => false)
    port map(
      preds => place_1293_preds,
      succs => place_1293_succs,
      token => place_1293_token,
      clk   => clk,
      reset => reset);

  place_1294_preds(0) <= transition_821_symbol_out;
  place_1294_succs(0) <= transition_826_symbol_out;
  place_1294 : place
    generic map(marking => false)
    port map(
      preds => place_1294_preds,
      succs => place_1294_succs,
      token => place_1294_token,
      clk   => clk,
      reset => reset);

  place_1295_preds(0) <= transition_829_symbol_out;
  place_1295_succs(0) <= transition_836_symbol_out;
  place_1295 : place
    generic map(marking => false)
    port map(
      preds => place_1295_preds,
      succs => place_1295_succs,
      token => place_1295_token,
      clk   => clk,
      reset => reset);

  place_1296_preds(0) <= transition_836_symbol_out;
  place_1296_succs(0) <= transition_835_symbol_out;
  place_1296 : place
    generic map(marking => false)
    port map(
      preds => place_1296_preds,
      succs => place_1296_succs,
      token => place_1296_token,
      clk   => clk,
      reset => reset);

  place_1297_preds(0) <= transition_834_symbol_out;
  place_1297_succs(0) <= transition_884_symbol_out;
  place_1297 : place
    generic map(marking => false)
    port map(
      preds => place_1297_preds,
      succs => place_1297_succs,
      token => place_1297_token,
      clk   => clk,
      reset => reset);

  place_1298_preds(0) <= transition_840_symbol_out;
  place_1298_succs(0) <= transition_858_symbol_out;
  place_1298 : place
    generic map(marking => false)
    port map(
      preds => place_1298_preds,
      succs => place_1298_succs,
      token => place_1298_token,
      clk   => clk,
      reset => reset);

  place_1299_preds(0) <= transition_17_symbol_out;
  place_1299_succs(0) <= transition_837_symbol_out;
  place_1299 : place
    generic map(marking => false)
    port map(
      preds => place_1299_preds,
      succs => place_1299_succs,
      token => place_1299_token,
      clk   => clk,
      reset => reset);

  place_1300_preds(0) <= transition_4_symbol_out;
  place_1300_succs(0) <= transition_76_symbol_out;
  place_1300 : place
    generic map(marking => false)
    port map(
      preds => place_1300_preds,
      succs => place_1300_succs,
      token => place_1300_token,
      clk   => clk,
      reset => reset);

  place_1301_preds(0) <= transition_847_symbol_out;
  place_1301_succs(0) <= transition_858_symbol_out;
  place_1301 : place
    generic map(marking => false)
    port map(
      preds => place_1301_preds,
      succs => place_1301_succs,
      token => place_1301_token,
      clk   => clk,
      reset => reset);

  place_1302_preds(0) <= transition_17_symbol_out;
  place_1302_succs(0) <= transition_844_symbol_out;
  place_1302 : place
    generic map(marking => false)
    port map(
      preds => place_1302_preds,
      succs => place_1302_succs,
      token => place_1302_token,
      clk   => clk,
      reset => reset);

  place_1303_preds(0) <= transition_858_symbol_out;
  place_1303_succs(0) <= transition_851_symbol_out;
  place_1303 : place
    generic map(marking => false)
    port map(
      preds => place_1303_preds,
      succs => place_1303_succs,
      token => place_1303_token,
      clk   => clk,
      reset => reset);

  place_1304_preds(0) <= transition_854_symbol_out;
  place_1304_succs(0) <= transition_873_symbol_out;
  place_1304 : place
    generic map(marking => false)
    port map(
      preds => place_1304_preds,
      succs => place_1304_succs,
      token => place_1304_token,
      clk   => clk,
      reset => reset);

  place_1305_preds(0) <= transition_862_symbol_out;
  place_1305_succs(0) <= transition_873_symbol_out;
  place_1305 : place
    generic map(marking => false)
    port map(
      preds => place_1305_preds,
      succs => place_1305_succs,
      token => place_1305_token,
      clk   => clk,
      reset => reset);

  place_1306_preds(0) <= transition_17_symbol_out;
  place_1306_succs(0) <= transition_859_symbol_out;
  place_1306 : place
    generic map(marking => false)
    port map(
      preds => place_1306_preds,
      succs => place_1306_succs,
      token => place_1306_token,
      clk   => clk,
      reset => reset);

  place_1307_preds(0) <= transition_873_symbol_out;
  place_1307_succs(0) <= transition_866_symbol_out;
  place_1307 : place
    generic map(marking => false)
    port map(
      preds => place_1307_preds,
      succs => place_1307_succs,
      token => place_1307_token,
      clk   => clk,
      reset => reset);

  place_1308_preds(0) <= transition_869_symbol_out;
  place_1308_succs(0) <= transition_874_symbol_out;
  place_1308 : place
    generic map(marking => false)
    port map(
      preds => place_1308_preds,
      succs => place_1308_succs,
      token => place_1308_token,
      clk   => clk,
      reset => reset);

  place_1309_preds(0) <= transition_877_symbol_out;
  place_1309_succs(0) <= transition_884_symbol_out;
  place_1309 : place
    generic map(marking => false)
    port map(
      preds => place_1309_preds,
      succs => place_1309_succs,
      token => place_1309_token,
      clk   => clk,
      reset => reset);

  place_1310_preds(0) <= transition_86_symbol_out;
  place_1310_succs(0) <= transition_97_symbol_out;
  place_1310 : place
    generic map(marking => false)
    port map(
      preds => place_1310_preds,
      succs => place_1310_succs,
      token => place_1310_token,
      clk   => clk,
      reset => reset);

  place_1311_preds(0) <= transition_884_symbol_out;
  place_1311_succs(0) <= transition_883_symbol_out;
  place_1311 : place
    generic map(marking => false)
    port map(
      preds => place_1311_preds,
      succs => place_1311_succs,
      token => place_1311_token,
      clk   => clk,
      reset => reset);

  place_1312_preds(0) <= transition_882_symbol_out;
  place_1312_succs(0) <= transition_932_symbol_out;
  place_1312 : place
    generic map(marking => false)
    port map(
      preds => place_1312_preds,
      succs => place_1312_succs,
      token => place_1312_token,
      clk   => clk,
      reset => reset);

  place_1313_preds(0) <= transition_888_symbol_out;
  place_1313_succs(0) <= transition_906_symbol_out;
  place_1313 : place
    generic map(marking => false)
    port map(
      preds => place_1313_preds,
      succs => place_1313_succs,
      token => place_1313_token,
      clk   => clk,
      reset => reset);

  place_1314_preds(0) <= transition_17_symbol_out;
  place_1314_succs(0) <= transition_885_symbol_out;
  place_1314 : place
    generic map(marking => false)
    port map(
      preds => place_1314_preds,
      succs => place_1314_succs,
      token => place_1314_token,
      clk   => clk,
      reset => reset);

  place_1315_preds(0) <= transition_895_symbol_out;
  place_1315_succs(0) <= transition_906_symbol_out;
  place_1315 : place
    generic map(marking => false)
    port map(
      preds => place_1315_preds,
      succs => place_1315_succs,
      token => place_1315_token,
      clk   => clk,
      reset => reset);

  place_1316_preds(0) <= transition_17_symbol_out;
  place_1316_succs(0) <= transition_892_symbol_out;
  place_1316 : place
    generic map(marking => false)
    port map(
      preds => place_1316_preds,
      succs => place_1316_succs,
      token => place_1316_token,
      clk   => clk,
      reset => reset);

  place_1317_preds(0) <= transition_906_symbol_out;
  place_1317_succs(0) <= transition_899_symbol_out;
  place_1317 : place
    generic map(marking => false)
    port map(
      preds => place_1317_preds,
      succs => place_1317_succs,
      token => place_1317_token,
      clk   => clk,
      reset => reset);

  place_1318_preds(0) <= transition_902_symbol_out;
  place_1318_succs(0) <= transition_921_symbol_out;
  place_1318 : place
    generic map(marking => false)
    port map(
      preds => place_1318_preds,
      succs => place_1318_succs,
      token => place_1318_token,
      clk   => clk,
      reset => reset);

  place_1319_preds(0) <= transition_4_symbol_out;
  place_1319_succs(0) <= transition_83_symbol_out;
  place_1319 : place
    generic map(marking => false)
    port map(
      preds => place_1319_preds,
      succs => place_1319_succs,
      token => place_1319_token,
      clk   => clk,
      reset => reset);

  place_1320_preds(0) <= transition_910_symbol_out;
  place_1320_succs(0) <= transition_921_symbol_out;
  place_1320 : place
    generic map(marking => false)
    port map(
      preds => place_1320_preds,
      succs => place_1320_succs,
      token => place_1320_token,
      clk   => clk,
      reset => reset);

  place_1321_preds(0) <= transition_17_symbol_out;
  place_1321_succs(0) <= transition_907_symbol_out;
  place_1321 : place
    generic map(marking => false)
    port map(
      preds => place_1321_preds,
      succs => place_1321_succs,
      token => place_1321_token,
      clk   => clk,
      reset => reset);

  place_1322_preds(0) <= transition_921_symbol_out;
  place_1322_succs(0) <= transition_914_symbol_out;
  place_1322 : place
    generic map(marking => false)
    port map(
      preds => place_1322_preds,
      succs => place_1322_succs,
      token => place_1322_token,
      clk   => clk,
      reset => reset);

  place_1323_preds(0) <= transition_917_symbol_out;
  place_1323_succs(0) <= transition_922_symbol_out;
  place_1323 : place
    generic map(marking => false)
    port map(
      preds => place_1323_preds,
      succs => place_1323_succs,
      token => place_1323_token,
      clk   => clk,
      reset => reset);

  place_1324_preds(0) <= transition_97_symbol_out;
  place_1324_succs(0) <= transition_90_symbol_out;
  place_1324 : place
    generic map(marking => false)
    port map(
      preds => place_1324_preds,
      succs => place_1324_succs,
      token => place_1324_token,
      clk   => clk,
      reset => reset);

  place_1325_preds(0) <= transition_925_symbol_out;
  place_1325_succs(0) <= transition_932_symbol_out;
  place_1325 : place
    generic map(marking => false)
    port map(
      preds => place_1325_preds,
      succs => place_1325_succs,
      token => place_1325_token,
      clk   => clk,
      reset => reset);

  place_1326_preds(0) <= transition_932_symbol_out;
  place_1326_succs(0) <= transition_931_symbol_out;
  place_1326 : place
    generic map(marking => false)
    port map(
      preds => place_1326_preds,
      succs => place_1326_succs,
      token => place_1326_token,
      clk   => clk,
      reset => reset);

  place_1327_preds(0) <= transition_930_symbol_out;
  place_1327_succs(0) <= transition_980_symbol_out;
  place_1327 : place
    generic map(marking => false)
    port map(
      preds => place_1327_preds,
      succs => place_1327_succs,
      token => place_1327_token,
      clk   => clk,
      reset => reset);

  place_1328_preds(0) <= transition_936_symbol_out;
  place_1328_succs(0) <= transition_954_symbol_out;
  place_1328 : place
    generic map(marking => false)
    port map(
      preds => place_1328_preds,
      succs => place_1328_succs,
      token => place_1328_token,
      clk   => clk,
      reset => reset);

  place_1329_preds(0) <= transition_93_symbol_out;
  place_1329_succs(0) <= transition_112_symbol_out;
  place_1329 : place
    generic map(marking => false)
    port map(
      preds => place_1329_preds,
      succs => place_1329_succs,
      token => place_1329_token,
      clk   => clk,
      reset => reset);

  place_1330_preds(0) <= transition_17_symbol_out;
  place_1330_succs(0) <= transition_933_symbol_out;
  place_1330 : place
    generic map(marking => false)
    port map(
      preds => place_1330_preds,
      succs => place_1330_succs,
      token => place_1330_token,
      clk   => clk,
      reset => reset);

  place_1331_preds(0) <= transition_943_symbol_out;
  place_1331_succs(0) <= transition_954_symbol_out;
  place_1331 : place
    generic map(marking => false)
    port map(
      preds => place_1331_preds,
      succs => place_1331_succs,
      token => place_1331_token,
      clk   => clk,
      reset => reset);

  place_1332_preds(0) <= transition_17_symbol_out;
  place_1332_succs(0) <= transition_940_symbol_out;
  place_1332 : place
    generic map(marking => false)
    port map(
      preds => place_1332_preds,
      succs => place_1332_succs,
      token => place_1332_token,
      clk   => clk,
      reset => reset);

  place_1333_preds(0) <= transition_954_symbol_out;
  place_1333_succs(0) <= transition_947_symbol_out;
  place_1333 : place
    generic map(marking => false)
    port map(
      preds => place_1333_preds,
      succs => place_1333_succs,
      token => place_1333_token,
      clk   => clk,
      reset => reset);

  place_1334_preds(0) <= transition_950_symbol_out;
  place_1334_succs(0) <= transition_969_symbol_out;
  place_1334 : place
    generic map(marking => false)
    port map(
      preds => place_1334_preds,
      succs => place_1334_succs,
      token => place_1334_token,
      clk   => clk,
      reset => reset);

  place_1335_preds(0) <= transition_958_symbol_out;
  place_1335_succs(0) <= transition_969_symbol_out;
  place_1335 : place
    generic map(marking => false)
    port map(
      preds => place_1335_preds,
      succs => place_1335_succs,
      token => place_1335_token,
      clk   => clk,
      reset => reset);

  place_1336_preds(0) <= transition_17_symbol_out;
  place_1336_succs(0) <= transition_955_symbol_out;
  place_1336 : place
    generic map(marking => false)
    port map(
      preds => place_1336_preds,
      succs => place_1336_succs,
      token => place_1336_token,
      clk   => clk,
      reset => reset);

  place_1337_preds(0) <= transition_969_symbol_out;
  place_1337_succs(0) <= transition_962_symbol_out;
  place_1337 : place
    generic map(marking => false)
    port map(
      preds => place_1337_preds,
      succs => place_1337_succs,
      token => place_1337_token,
      clk   => clk,
      reset => reset);

  place_1338_preds(0) <= transition_965_symbol_out;
  place_1338_succs(0) <= transition_970_symbol_out;
  place_1338 : place
    generic map(marking => false)
    port map(
      preds => place_1338_preds,
      succs => place_1338_succs,
      token => place_1338_token,
      clk   => clk,
      reset => reset);

  place_1339_preds(0) <= transition_973_symbol_out;
  place_1339_succs(0) <= transition_980_symbol_out;
  place_1339 : place
    generic map(marking => false)
    port map(
      preds => place_1339_preds,
      succs => place_1339_succs,
      token => place_1339_token,
      clk   => clk,
      reset => reset);

  place_1340_preds(0) <= transition_980_symbol_out;
  place_1340_succs(0) <= transition_979_symbol_out;
  place_1340 : place
    generic map(marking => false)
    port map(
      preds => place_1340_preds,
      succs => place_1340_succs,
      token => place_1340_token,
      clk   => clk,
      reset => reset);

  place_1341_preds(0) <= transition_978_symbol_out;
  place_1341_succs(0) <= transition_1028_symbol_out;
  place_1341 : place
    generic map(marking => false)
    port map(
      preds => place_1341_preds,
      succs => place_1341_succs,
      token => place_1341_token,
      clk   => clk,
      reset => reset);

  place_1342_preds(0) <= transition_984_symbol_out;
  place_1342_succs(0) <= transition_1002_symbol_out;
  place_1342 : place
    generic map(marking => false)
    port map(
      preds => place_1342_preds,
      succs => place_1342_succs,
      token => place_1342_token,
      clk   => clk,
      reset => reset);

  place_1343_preds(0) <= transition_17_symbol_out;
  place_1343_succs(0) <= transition_981_symbol_out;
  place_1343 : place
    generic map(marking => false)
    port map(
      preds => place_1343_preds,
      succs => place_1343_succs,
      token => place_1343_token,
      clk   => clk,
      reset => reset);

  place_1344_preds(0) <= transition_991_symbol_out;
  place_1344_succs(0) <= transition_1002_symbol_out;
  place_1344 : place
    generic map(marking => false)
    port map(
      preds => place_1344_preds,
      succs => place_1344_succs,
      token => place_1344_token,
      clk   => clk,
      reset => reset);

  place_1345_preds(0) <= transition_17_symbol_out;
  place_1345_succs(0) <= transition_988_symbol_out;
  place_1345 : place
    generic map(marking => false)
    port map(
      preds => place_1345_preds,
      succs => place_1345_succs,
      token => place_1345_token,
      clk   => clk,
      reset => reset);

  place_1346_preds(0) <= transition_1002_symbol_out;
  place_1346_succs(0) <= transition_995_symbol_out;
  place_1346 : place
    generic map(marking => false)
    port map(
      preds => place_1346_preds,
      succs => place_1346_succs,
      token => place_1346_token,
      clk   => clk,
      reset => reset);

  place_1347_preds(0) <= transition_998_symbol_out;
  place_1347_succs(0) <= transition_1017_symbol_out;
  place_1347 : place
    generic map(marking => false)
    port map(
      preds => place_1347_preds,
      succs => place_1347_succs,
      token => place_1347_token,
      clk   => clk,
      reset => reset);

  place_1348_preds(0) <= transition_1006_symbol_out;
  place_1348_succs(0) <= transition_1017_symbol_out;
  place_1348 : place
    generic map(marking => false)
    port map(
      preds => place_1348_preds,
      succs => place_1348_succs,
      token => place_1348_token,
      clk   => clk,
      reset => reset);

  place_1349_preds(0) <= transition_17_symbol_out;
  place_1349_succs(0) <= transition_1003_symbol_out;
  place_1349 : place
    generic map(marking => false)
    port map(
      preds => place_1349_preds,
      succs => place_1349_succs,
      token => place_1349_token,
      clk   => clk,
      reset => reset);

  place_1350_preds(0) <= transition_1017_symbol_out;
  place_1350_succs(0) <= transition_1010_symbol_out;
  place_1350 : place
    generic map(marking => false)
    port map(
      preds => place_1350_preds,
      succs => place_1350_succs,
      token => place_1350_token,
      clk   => clk,
      reset => reset);

  place_1351_preds(0) <= transition_1013_symbol_out;
  place_1351_succs(0) <= transition_1018_symbol_out;
  place_1351 : place
    generic map(marking => false)
    port map(
      preds => place_1351_preds,
      succs => place_1351_succs,
      token => place_1351_token,
      clk   => clk,
      reset => reset);

  place_1352_preds(0) <= transition_101_symbol_out;
  place_1352_succs(0) <= transition_112_symbol_out;
  place_1352 : place
    generic map(marking => false)
    port map(
      preds => place_1352_preds,
      succs => place_1352_succs,
      token => place_1352_token,
      clk   => clk,
      reset => reset);

  place_1353_preds(0) <= transition_1021_symbol_out;
  place_1353_succs(0) <= transition_1028_symbol_out;
  place_1353 : place
    generic map(marking => false)
    port map(
      preds => place_1353_preds,
      succs => place_1353_succs,
      token => place_1353_token,
      clk   => clk,
      reset => reset);

  place_1354_preds(0) <= transition_1028_symbol_out;
  place_1354_succs(0) <= transition_1027_symbol_out;
  place_1354 : place
    generic map(marking => false)
    port map(
      preds => place_1354_preds,
      succs => place_1354_succs,
      token => place_1354_token,
      clk   => clk,
      reset => reset);

  place_1355_preds(0) <= transition_1026_symbol_out;
  place_1355_succs(0) <= transition_1031_symbol_out;
  place_1355 : place
    generic map(marking => false)
    port map(
      preds => place_1355_preds,
      succs => place_1355_succs,
      token => place_1355_token,
      clk   => clk,
      reset => reset);

  place_1356_preds(0) <= transition_1030_symbol_out;
  place_1356_succs(0) <= transition_1034_symbol_out;
  place_1356 : place
    generic map(marking => false)
    port map(
      preds => place_1356_preds,
      succs => place_1356_succs,
      token => place_1356_token,
      clk   => clk,
      reset => reset);

  place_1357_preds(0) <= transition_1033_symbol_out;
  place_1357_succs(0) <= transition_1035_symbol_out;
  place_1357 : place
    generic map(marking => false)
    port map(
      preds => place_1357_preds,
      succs => place_1357_succs,
      token => place_1357_token,
      clk   => clk,
      reset => reset);

  place_1358_preds(0) <= transition_1037_symbol_out;
  place_1358_succs(0) <= transition_1041_symbol_out;
  place_1358 : place
    generic map(marking => false)
    port map(
      preds => place_1358_preds,
      succs => place_1358_succs,
      token => place_1358_token,
      clk   => clk,
      reset => reset);

  place_1359_preds(0) <= transition_4_symbol_out;
  place_1359_succs(0) <= transition_98_symbol_out;
  place_1359 : place
    generic map(marking => false)
    port map(
      preds => place_1359_preds,
      succs => place_1359_succs,
      token => place_1359_token,
      clk   => clk,
      reset => reset);

  place_1360_preds(0) <= transition_1040_symbol_out;
  place_1360_succs(0) <= transition_1042_symbol_out;
  place_1360 : place
    generic map(marking => false)
    port map(
      preds => place_1360_preds,
      succs => place_1360_succs,
      token => place_1360_token,
      clk   => clk,
      reset => reset);

  place_1361_preds(0) <= transition_1035_symbol_out;
  place_1361_succs(0) <= transition_1038_symbol_out;
  place_1361 : place
    generic map(marking => false)
    port map(
      preds => place_1361_preds,
      succs => place_1361_succs,
      token => place_1361_token,
      clk   => clk,
      reset => reset);

  place_1362_preds(0) <= transition_1046_symbol_out;
  place_1362_succs(0) <= transition_1070_symbol_out;
  place_1362 : place
    generic map(marking => false)
    port map(
      preds => place_1362_preds,
      succs => place_1362_succs,
      token => place_1362_token,
      clk   => clk,
      reset => reset);

  place_1363_preds(0) <= transition_1042_symbol_out;
  place_1363_succs(0) <= transition_1043_symbol_out;
  place_1363 : place
    generic map(marking => false)
    port map(
      preds => place_1363_preds,
      succs => place_1363_succs,
      token => place_1363_token,
      clk   => clk,
      reset => reset);

  place_1364_preds(0) <= transition_1051_symbol_out;
  place_1364_succs(0) <= transition_1055_symbol_out;
  place_1364 : place
    generic map(marking => false)
    port map(
      preds => place_1364_preds,
      succs => place_1364_succs,
      token => place_1364_token,
      clk   => clk,
      reset => reset);

  place_1365_preds(0) <= transition_1_symbol_out;
  place_1365_succs(0) <= transition_20_symbol_out;
  place_1365 : place
    generic map(marking => false)
    port map(
      preds => place_1365_preds,
      succs => place_1365_succs,
      token => place_1365_token,
      clk   => clk,
      reset => reset);

  place_1366_preds(0) <= transition_112_symbol_out;
  place_1366_succs(0) <= transition_105_symbol_out;
  place_1366 : place
    generic map(marking => false)
    port map(
      preds => place_1366_preds,
      succs => place_1366_succs,
      token => place_1366_token,
      clk   => clk,
      reset => reset);

  place_1367_preds(0) <= transition_1054_symbol_out;
  place_1367_succs(0) <= transition_1056_symbol_out;
  place_1367 : place
    generic map(marking => false)
    port map(
      preds => place_1367_preds,
      succs => place_1367_succs,
      token => place_1367_token,
      clk   => clk,
      reset => reset);

  place_1368_preds(0) <= transition_1042_symbol_out;
  place_1368_succs(0) <= transition_1052_symbol_out;
  place_1368 : place
    generic map(marking => false)
    port map(
      preds => place_1368_preds,
      succs => place_1368_succs,
      token => place_1368_token,
      clk   => clk,
      reset => reset);

  place_1369_preds(0) <= transition_1059_symbol_out;
  place_1369_succs(0) <= transition_1078_symbol_out;
  place_1369 : place
    generic map(marking => false)
    port map(
      preds => place_1369_preds,
      succs => place_1369_succs,
      token => place_1369_token,
      clk   => clk,
      reset => reset);

  place_1370_preds(0) <= transition_1070_symbol_out;
  place_1370_succs(0) <= transition_1063_symbol_out;
  place_1370 : place
    generic map(marking => false)
    port map(
      preds => place_1370_preds,
      succs => place_1370_succs,
      token => place_1370_token,
      clk   => clk,
      reset => reset);

  place_1371_preds(0) <= transition_108_symbol_out;
  place_1371_succs(0) <= transition_113_symbol_out;
  place_1371 : place
    generic map(marking => false)
    port map(
      preds => place_1371_preds,
      succs => place_1371_succs,
      token => place_1371_token,
      clk   => clk,
      reset => reset);

  place_1372_preds(0) <= transition_1066_symbol_out;
  place_1372_succs(0) <= transition_1078_symbol_out;
  place_1372 : place
    generic map(marking => false)
    port map(
      preds => place_1372_preds,
      succs => place_1372_succs,
      token => place_1372_token,
      clk   => clk,
      reset => reset);

  place_1373_preds(0) <= transition_1035_symbol_out;
  place_1373_succs(0) <= transition_1070_symbol_out;
  place_1373 : place
    generic map(marking => false)
    port map(
      preds => place_1373_preds,
      succs => place_1373_succs,
      token => place_1373_token,
      clk   => clk,
      reset => reset);

  place_1374_preds(0) <= transition_1078_symbol_out;
  place_1374_succs(0) <= transition_1071_symbol_out;
  place_1374 : place
    generic map(marking => false)
    port map(
      preds => place_1374_preds,
      succs => place_1374_succs,
      token => place_1374_token,
      clk   => clk,
      reset => reset);

  place_1375_preds(0) <= transition_1074_symbol_out;
  place_1375_succs(0) <= transition_1081_symbol_out;
  place_1375 : place
    generic map(marking => false)
    port map(
      preds => place_1375_preds,
      succs => place_1375_succs,
      token => place_1375_token,
      clk   => clk,
      reset => reset);

  place_1376_preds(0) <= transition_1080_symbol_out;
  place_1376_succs(0) <= transition_2_symbol_out;
  place_1376 : place
    generic map(marking => false)
    port map(
      preds => place_1376_preds,
      succs => place_1376_succs,
      token => place_1376_token,
      clk   => clk,
      reset => reset);

  place_1377_preds(0) <= transition_116_symbol_out;
  place_1377_succs(0) <= transition_216_symbol_out;
  place_1377 : place
    generic map(marking => false)
    port map(
      preds => place_1377_preds,
      succs => place_1377_succs,
      token => place_1377_token,
      clk   => clk,
      reset => reset);

  place_1378_preds(0) <= transition_19_symbol_out;
  place_1378_succs(0) <= transition_21_symbol_out;
  place_1378 : place
    generic map(marking => false)
    port map(
      preds => place_1378_preds,
      succs => place_1378_succs,
      token => place_1378_token,
      clk   => clk,
      reset => reset);

  place_1379_preds(0) <= transition_123_symbol_out;
  place_1379_succs(0) <= transition_141_symbol_out;
  place_1379 : place
    generic map(marking => false)
    port map(
      preds => place_1379_preds,
      succs => place_1379_succs,
      token => place_1379_token,
      clk   => clk,
      reset => reset);

  place_1380_preds(0) <= transition_4_symbol_out;
  place_1380_succs(0) <= transition_120_symbol_out;
  place_1380 : place
    generic map(marking => false)
    port map(
      preds => place_1380_preds,
      succs => place_1380_succs,
      token => place_1380_token,
      clk   => clk,
      reset => reset);

  place_1381_preds(0) <= transition_130_symbol_out;
  place_1381_succs(0) <= transition_141_symbol_out;
  place_1381 : place
    generic map(marking => false)
    port map(
      preds => place_1381_preds,
      succs => place_1381_succs,
      token => place_1381_token,
      clk   => clk,
      reset => reset);

  place_1382_preds(0) <= transition_4_symbol_out;
  place_1382_succs(0) <= transition_127_symbol_out;
  place_1382 : place
    generic map(marking => false)
    port map(
      preds => place_1382_preds,
      succs => place_1382_succs,
      token => place_1382_token,
      clk   => clk,
      reset => reset);

  place_1383_preds(0) <= transition_141_symbol_out;
  place_1383_succs(0) <= transition_134_symbol_out;
  place_1383 : place
    generic map(marking => false)
    port map(
      preds => place_1383_preds,
      succs => place_1383_succs,
      token => place_1383_token,
      clk   => clk,
      reset => reset);

  place_1384_preds(0) <= transition_137_symbol_out;
  place_1384_succs(0) <= transition_142_symbol_out;
  place_1384 : place
    generic map(marking => false)
    port map(
      preds => place_1384_preds,
      succs => place_1384_succs,
      token => place_1384_token,
      clk   => clk,
      reset => reset);

  place_1385_preds(0) <= transition_145_symbol_out;
  place_1385_succs(0) <= transition_163_symbol_out;
  place_1385 : place
    generic map(marking => false)
    port map(
      preds => place_1385_preds,
      succs => place_1385_succs,
      token => place_1385_token,
      clk   => clk,
      reset => reset);

  transition_1_preds(0) <= place_0_token;
  transition_1 : transition
    port map(
      preds      => transition_1_preds,
      symbol_out => transition_1_symbol_out,
      symbol_in  => true);

  transition_2_preds(0) <= place_1376_token;
  transition_2 : transition
    port map(
      preds      => transition_2_preds,
      symbol_out => transition_2_symbol_out,
      symbol_in  => true);

  transition_3_preds(0) <= place_1108_token;
  transition_3_preds(1) <= place_1133_token;
  transition_3 : transition
    port map(
      preds      => transition_3_preds,
      symbol_out => transition_3_symbol_out,
      symbol_in  => true);

  transition_4_preds(0) <= place_1132_token;
  transition_4 : transition
    port map(
      preds      => transition_4_preds,
      symbol_out => transition_4_symbol_out,
      symbol_in  => true);

  transition_5_preds(0) <= place_1105_token;
  transition_5_preds(1) <= place_1109_token;
  transition_5 : transition
    port map(
      preds      => transition_5_preds,
      symbol_out => transition_5_symbol_out,
      symbol_in  => true);

  transition_7_preds(0) <= place_6_token;
  transition_7 : transition
    port map(
      preds      => transition_7_preds,
      symbol_out => transition_7_symbol_out,
      symbol_in  => LambdaIn(1));

  transition_8_preds(0) <= place_6_token;
  transition_8 : transition
    port map(
      preds      => transition_8_preds,
      symbol_out => transition_8_symbol_out,
      symbol_in  => LambdaIn(2));

  transition_9_preds(0) <= place_1181_token;
  LambdaOut(1) <= transition_9_symbol_out;
  transition_9 : transition
    port map(
      preds      => transition_9_preds,
      symbol_out => transition_9_symbol_out,
      symbol_in  => true);

  transition_10_preds(0) <= place_1113_token;
  transition_10_preds(1) <= place_1116_token;
  transition_10 : transition
    port map(
      preds      => transition_10_preds,
      symbol_out => transition_10_symbol_out,
      symbol_in  => true);

  transition_11_preds(0) <= place_1227_token;
  transition_11 : transition
    port map(
      preds      => transition_11_preds,
      symbol_out => transition_11_symbol_out,
      symbol_in  => true);

  transition_12_preds(0) <= place_1177_token;
  transition_12_preds(1) <= place_1180_token;
  transition_12 : transition
    port map(
      preds      => transition_12_preds,
      symbol_out => transition_12_symbol_out,
      symbol_in  => true);

  transition_14_preds(0) <= place_13_token;
  transition_14 : transition
    port map(
      preds      => transition_14_preds,
      symbol_out => transition_14_symbol_out,
      symbol_in  => LambdaIn(3));

  transition_15_preds(0) <= place_13_token;
  transition_15 : transition
    port map(
      preds      => transition_15_preds,
      symbol_out => transition_15_symbol_out,
      symbol_in  => LambdaIn(4));

  transition_16_preds(0) <= place_1273_token;
  LambdaOut(2) <= transition_16_symbol_out;
  transition_16 : transition
    port map(
      preds      => transition_16_preds,
      symbol_out => transition_16_symbol_out,
      symbol_in  => true);

  transition_17_preds(0) <= place_1111_token;
  transition_17 : transition
    port map(
      preds      => transition_17_preds,
      symbol_out => transition_17_symbol_out,
      symbol_in  => true);

  transition_19_preds(0) <= place_18_token;
  transition_19 : transition
    port map(
      preds      => transition_19_preds,
      symbol_out => transition_19_symbol_out,
      symbol_in  => LambdaIn(5));

  transition_20_preds(0) <= place_1365_token;
  LambdaOut(3) <= transition_20_symbol_out;
  transition_20 : transition
    port map(
      preds      => transition_20_preds,
      symbol_out => transition_20_symbol_out,
      symbol_in  => true);

  transition_21_preds(0) <= place_1378_token;
  transition_21 : transition
    port map(
      preds      => transition_21_preds,
      symbol_out => transition_21_symbol_out,
      symbol_in  => true);

  transition_22_preds(0) <= place_1088_token;
  transition_22 : transition
    port map(
      preds      => transition_22_preds,
      symbol_out => transition_22_symbol_out,
      symbol_in  => true);

  transition_23_preds(0) <= place_1094_token;
  transition_23 : transition
    port map(
      preds      => transition_23_preds,
      symbol_out => transition_23_symbol_out,
      symbol_in  => true);

  transition_25_preds(0) <= place_24_token;
  transition_25 : transition
    port map(
      preds      => transition_25_preds,
      symbol_out => transition_25_symbol_out,
      symbol_in  => LambdaIn(6));

  transition_26_preds(0) <= place_1103_token;
  LambdaOut(4) <= transition_26_symbol_out;
  transition_26 : transition
    port map(
      preds      => transition_26_preds,
      symbol_out => transition_26_symbol_out,
      symbol_in  => true);

  transition_27_preds(0) <= place_1119_token;
  LambdaOut(5) <= transition_27_symbol_out;
  transition_27 : transition
    port map(
      preds      => transition_27_preds,
      symbol_out => transition_27_symbol_out,
      symbol_in  => true);

  transition_29_preds(0) <= place_28_token;
  transition_29 : transition
    port map(
      preds      => transition_29_preds,
      symbol_out => transition_29_symbol_out,
      symbol_in  => LambdaIn(7));

  transition_30_preds(0) <= place_1129_token;
  LambdaOut(6) <= transition_30_symbol_out;
  transition_30 : transition
    port map(
      preds      => transition_30_preds,
      symbol_out => transition_30_symbol_out,
      symbol_in  => true);

  transition_31_preds(0) <= place_1143_token;
  LambdaOut(7) <= transition_31_symbol_out;
  transition_31 : transition
    port map(
      preds      => transition_31_preds,
      symbol_out => transition_31_symbol_out,
      symbol_in  => true);

  transition_32_preds(0) <= place_1168_token;
  LambdaOut(8) <= transition_32_symbol_out;
  transition_32 : transition
    port map(
      preds      => transition_32_preds,
      symbol_out => transition_32_symbol_out,
      symbol_in  => true);

  transition_33_preds(0) <= place_36_token;
  transition_33 : transition
    port map(
      preds      => transition_33_preds,
      symbol_out => transition_33_symbol_out,
      symbol_in  => LambdaIn(8));

  transition_34_preds(0) <= place_37_token;
  LambdaOut(9) <= transition_34_symbol_out;
  transition_34 : transition
    port map(
      preds      => transition_34_preds,
      symbol_out => transition_34_symbol_out,
      symbol_in  => true);

  transition_35_preds(0) <= place_38_token;
  transition_35 : transition
    port map(
      preds      => transition_35_preds,
      symbol_out => transition_35_symbol_out,
      symbol_in  => LambdaIn(9));

  transition_39_preds(0) <= place_1189_token;
  LambdaOut(10) <= transition_39_symbol_out;
  transition_39 : transition
    port map(
      preds      => transition_39_preds,
      symbol_out => transition_39_symbol_out,
      symbol_in  => true);

  transition_40_preds(0) <= place_43_token;
  transition_40 : transition
    port map(
      preds      => transition_40_preds,
      symbol_out => transition_40_symbol_out,
      symbol_in  => LambdaIn(10));

  transition_41_preds(0) <= place_44_token;
  LambdaOut(11) <= transition_41_symbol_out;
  transition_41 : transition
    port map(
      preds      => transition_41_preds,
      symbol_out => transition_41_symbol_out,
      symbol_in  => true);

  transition_42_preds(0) <= place_45_token;
  transition_42 : transition
    port map(
      preds      => transition_42_preds,
      symbol_out => transition_42_symbol_out,
      symbol_in  => LambdaIn(11));

  transition_46_preds(0) <= place_1194_token;
  LambdaOut(12) <= transition_46_symbol_out;
  transition_46 : transition
    port map(
      preds      => transition_46_preds,
      symbol_out => transition_46_symbol_out,
      symbol_in  => true);

  transition_47_preds(0) <= place_50_token;
  transition_47 : transition
    port map(
      preds      => transition_47_preds,
      symbol_out => transition_47_symbol_out,
      symbol_in  => LambdaIn(12));

  transition_48_preds(0) <= place_51_token;
  LambdaOut(13) <= transition_48_symbol_out;
  transition_48 : transition
    port map(
      preds      => transition_48_preds,
      symbol_out => transition_48_symbol_out,
      symbol_in  => true);

  transition_49_preds(0) <= place_52_token;
  transition_49 : transition
    port map(
      preds      => transition_49_preds,
      symbol_out => transition_49_symbol_out,
      symbol_in  => LambdaIn(13));

  transition_53_preds(0) <= place_1152_token;
  transition_53_preds(1) <= place_1176_token;
  transition_53 : transition
    port map(
      preds      => transition_53_preds,
      symbol_out => transition_53_symbol_out,
      symbol_in  => true);

  transition_54_preds(0) <= place_1237_token;
  LambdaOut(14) <= transition_54_symbol_out;
  transition_54 : transition
    port map(
      preds      => transition_54_preds,
      symbol_out => transition_54_symbol_out,
      symbol_in  => true);

  transition_55_preds(0) <= place_58_token;
  transition_55 : transition
    port map(
      preds      => transition_55_preds,
      symbol_out => transition_55_symbol_out,
      symbol_in  => LambdaIn(14));

  transition_56_preds(0) <= place_59_token;
  LambdaOut(15) <= transition_56_symbol_out;
  transition_56 : transition
    port map(
      preds      => transition_56_preds,
      symbol_out => transition_56_symbol_out,
      symbol_in  => true);

  transition_57_preds(0) <= place_60_token;
  transition_57 : transition
    port map(
      preds      => transition_57_preds,
      symbol_out => transition_57_symbol_out,
      symbol_in  => LambdaIn(15));

  transition_61_preds(0) <= place_1241_token;
  LambdaOut(16) <= transition_61_symbol_out;
  transition_61 : transition
    port map(
      preds      => transition_61_preds,
      symbol_out => transition_61_symbol_out,
      symbol_in  => true);

  transition_62_preds(0) <= place_65_token;
  transition_62 : transition
    port map(
      preds      => transition_62_preds,
      symbol_out => transition_62_symbol_out,
      symbol_in  => LambdaIn(16));

  transition_63_preds(0) <= place_66_token;
  LambdaOut(17) <= transition_63_symbol_out;
  transition_63 : transition
    port map(
      preds      => transition_63_preds,
      symbol_out => transition_63_symbol_out,
      symbol_in  => true);

  transition_64_preds(0) <= place_67_token;
  transition_64 : transition
    port map(
      preds      => transition_64_preds,
      symbol_out => transition_64_symbol_out,
      symbol_in  => LambdaIn(17));

  transition_68_preds(0) <= place_1200_token;
  transition_68_preds(1) <= place_1222_token;
  transition_68 : transition
    port map(
      preds      => transition_68_preds,
      symbol_out => transition_68_symbol_out,
      symbol_in  => true);

  transition_69_preds(0) <= place_1248_token;
  LambdaOut(18) <= transition_69_symbol_out;
  transition_69 : transition
    port map(
      preds      => transition_69_preds,
      symbol_out => transition_69_symbol_out,
      symbol_in  => true);

  transition_70_preds(0) <= place_73_token;
  transition_70 : transition
    port map(
      preds      => transition_70_preds,
      symbol_out => transition_70_symbol_out,
      symbol_in  => LambdaIn(18));

  transition_71_preds(0) <= place_74_token;
  LambdaOut(19) <= transition_71_symbol_out;
  transition_71 : transition
    port map(
      preds      => transition_71_preds,
      symbol_out => transition_71_symbol_out,
      symbol_in  => true);

  transition_72_preds(0) <= place_75_token;
  transition_72 : transition
    port map(
      preds      => transition_72_preds,
      symbol_out => transition_72_symbol_out,
      symbol_in  => LambdaIn(19));

  transition_76_preds(0) <= place_1300_token;
  LambdaOut(20) <= transition_76_symbol_out;
  transition_76 : transition
    port map(
      preds      => transition_76_preds,
      symbol_out => transition_76_symbol_out,
      symbol_in  => true);

  transition_77_preds(0) <= place_80_token;
  transition_77 : transition
    port map(
      preds      => transition_77_preds,
      symbol_out => transition_77_symbol_out,
      symbol_in  => LambdaIn(20));

  transition_78_preds(0) <= place_81_token;
  LambdaOut(21) <= transition_78_symbol_out;
  transition_78 : transition
    port map(
      preds      => transition_78_preds,
      symbol_out => transition_78_symbol_out,
      symbol_in  => true);

  transition_79_preds(0) <= place_82_token;
  transition_79 : transition
    port map(
      preds      => transition_79_preds,
      symbol_out => transition_79_symbol_out,
      symbol_in  => LambdaIn(21));

  transition_83_preds(0) <= place_1319_token;
  LambdaOut(22) <= transition_83_symbol_out;
  transition_83 : transition
    port map(
      preds      => transition_83_preds,
      symbol_out => transition_83_symbol_out,
      symbol_in  => true);

  transition_84_preds(0) <= place_87_token;
  transition_84 : transition
    port map(
      preds      => transition_84_preds,
      symbol_out => transition_84_symbol_out,
      symbol_in  => LambdaIn(22));

  transition_85_preds(0) <= place_88_token;
  LambdaOut(23) <= transition_85_symbol_out;
  transition_85 : transition
    port map(
      preds      => transition_85_preds,
      symbol_out => transition_85_symbol_out,
      symbol_in  => true);

  transition_86_preds(0) <= place_89_token;
  transition_86 : transition
    port map(
      preds      => transition_86_preds,
      symbol_out => transition_86_symbol_out,
      symbol_in  => LambdaIn(23));

  transition_90_preds(0) <= place_1324_token;
  LambdaOut(24) <= transition_90_symbol_out;
  transition_90 : transition
    port map(
      preds      => transition_90_preds,
      symbol_out => transition_90_symbol_out,
      symbol_in  => true);

  transition_91_preds(0) <= place_94_token;
  transition_91 : transition
    port map(
      preds      => transition_91_preds,
      symbol_out => transition_91_symbol_out,
      symbol_in  => LambdaIn(24));

  transition_92_preds(0) <= place_95_token;
  LambdaOut(25) <= transition_92_symbol_out;
  transition_92 : transition
    port map(
      preds      => transition_92_preds,
      symbol_out => transition_92_symbol_out,
      symbol_in  => true);

  transition_93_preds(0) <= place_96_token;
  transition_93 : transition
    port map(
      preds      => transition_93_preds,
      symbol_out => transition_93_symbol_out,
      symbol_in  => LambdaIn(25));

  transition_97_preds(0) <= place_1286_token;
  transition_97_preds(1) <= place_1310_token;
  transition_97 : transition
    port map(
      preds      => transition_97_preds,
      symbol_out => transition_97_symbol_out,
      symbol_in  => true);

  transition_98_preds(0) <= place_1359_token;
  LambdaOut(26) <= transition_98_symbol_out;
  transition_98 : transition
    port map(
      preds      => transition_98_preds,
      symbol_out => transition_98_symbol_out,
      symbol_in  => true);

  transition_99_preds(0) <= place_102_token;
  transition_99 : transition
    port map(
      preds      => transition_99_preds,
      symbol_out => transition_99_symbol_out,
      symbol_in  => LambdaIn(26));

  transition_100_preds(0) <= place_103_token;
  LambdaOut(27) <= transition_100_symbol_out;
  transition_100 : transition
    port map(
      preds      => transition_100_preds,
      symbol_out => transition_100_symbol_out,
      symbol_in  => true);

  transition_101_preds(0) <= place_104_token;
  transition_101 : transition
    port map(
      preds      => transition_101_preds,
      symbol_out => transition_101_symbol_out,
      symbol_in  => LambdaIn(27));

  transition_105_preds(0) <= place_1366_token;
  LambdaOut(28) <= transition_105_symbol_out;
  transition_105 : transition
    port map(
      preds      => transition_105_preds,
      symbol_out => transition_105_symbol_out,
      symbol_in  => true);

  transition_106_preds(0) <= place_109_token;
  transition_106 : transition
    port map(
      preds      => transition_106_preds,
      symbol_out => transition_106_symbol_out,
      symbol_in  => LambdaIn(28));

  transition_107_preds(0) <= place_110_token;
  LambdaOut(29) <= transition_107_symbol_out;
  transition_107 : transition
    port map(
      preds      => transition_107_preds,
      symbol_out => transition_107_symbol_out,
      symbol_in  => true);

  transition_108_preds(0) <= place_111_token;
  transition_108 : transition
    port map(
      preds      => transition_108_preds,
      symbol_out => transition_108_symbol_out,
      symbol_in  => LambdaIn(29));

  transition_112_preds(0) <= place_1329_token;
  transition_112_preds(1) <= place_1352_token;
  transition_112 : transition
    port map(
      preds      => transition_112_preds,
      symbol_out => transition_112_symbol_out,
      symbol_in  => true);

  transition_113_preds(0) <= place_1371_token;
  LambdaOut(30) <= transition_113_symbol_out;
  transition_113 : transition
    port map(
      preds      => transition_113_preds,
      symbol_out => transition_113_symbol_out,
      symbol_in  => true);

  transition_114_preds(0) <= place_117_token;
  transition_114 : transition
    port map(
      preds      => transition_114_preds,
      symbol_out => transition_114_symbol_out,
      symbol_in  => LambdaIn(30));

  transition_115_preds(0) <= place_118_token;
  LambdaOut(31) <= transition_115_symbol_out;
  transition_115 : transition
    port map(
      preds      => transition_115_preds,
      symbol_out => transition_115_symbol_out,
      symbol_in  => true);

  transition_116_preds(0) <= place_119_token;
  transition_116 : transition
    port map(
      preds      => transition_116_preds,
      symbol_out => transition_116_symbol_out,
      symbol_in  => LambdaIn(31));

  transition_120_preds(0) <= place_1380_token;
  LambdaOut(32) <= transition_120_symbol_out;
  transition_120 : transition
    port map(
      preds      => transition_120_preds,
      symbol_out => transition_120_symbol_out,
      symbol_in  => true);

  transition_121_preds(0) <= place_124_token;
  transition_121 : transition
    port map(
      preds      => transition_121_preds,
      symbol_out => transition_121_symbol_out,
      symbol_in  => LambdaIn(32));

  transition_122_preds(0) <= place_125_token;
  LambdaOut(33) <= transition_122_symbol_out;
  transition_122 : transition
    port map(
      preds      => transition_122_preds,
      symbol_out => transition_122_symbol_out,
      symbol_in  => true);

  transition_123_preds(0) <= place_126_token;
  transition_123 : transition
    port map(
      preds      => transition_123_preds,
      symbol_out => transition_123_symbol_out,
      symbol_in  => LambdaIn(33));

  transition_127_preds(0) <= place_1382_token;
  LambdaOut(34) <= transition_127_symbol_out;
  transition_127 : transition
    port map(
      preds      => transition_127_preds,
      symbol_out => transition_127_symbol_out,
      symbol_in  => true);

  transition_128_preds(0) <= place_131_token;
  transition_128 : transition
    port map(
      preds      => transition_128_preds,
      symbol_out => transition_128_symbol_out,
      symbol_in  => LambdaIn(34));

  transition_129_preds(0) <= place_132_token;
  LambdaOut(35) <= transition_129_symbol_out;
  transition_129 : transition
    port map(
      preds      => transition_129_preds,
      symbol_out => transition_129_symbol_out,
      symbol_in  => true);

  transition_130_preds(0) <= place_133_token;
  transition_130 : transition
    port map(
      preds      => transition_130_preds,
      symbol_out => transition_130_symbol_out,
      symbol_in  => LambdaIn(35));

  transition_134_preds(0) <= place_1383_token;
  LambdaOut(36) <= transition_134_symbol_out;
  transition_134 : transition
    port map(
      preds      => transition_134_preds,
      symbol_out => transition_134_symbol_out,
      symbol_in  => true);

  transition_135_preds(0) <= place_138_token;
  transition_135 : transition
    port map(
      preds      => transition_135_preds,
      symbol_out => transition_135_symbol_out,
      symbol_in  => LambdaIn(36));

  transition_136_preds(0) <= place_139_token;
  LambdaOut(37) <= transition_136_symbol_out;
  transition_136 : transition
    port map(
      preds      => transition_136_preds,
      symbol_out => transition_136_symbol_out,
      symbol_in  => true);

  transition_137_preds(0) <= place_140_token;
  transition_137 : transition
    port map(
      preds      => transition_137_preds,
      symbol_out => transition_137_symbol_out,
      symbol_in  => LambdaIn(37));

  transition_141_preds(0) <= place_1379_token;
  transition_141_preds(1) <= place_1381_token;
  transition_141 : transition
    port map(
      preds      => transition_141_preds,
      symbol_out => transition_141_symbol_out,
      symbol_in  => true);

  transition_142_preds(0) <= place_1384_token;
  LambdaOut(38) <= transition_142_symbol_out;
  transition_142 : transition
    port map(
      preds      => transition_142_preds,
      symbol_out => transition_142_symbol_out,
      symbol_in  => true);

  transition_143_preds(0) <= place_146_token;
  transition_143 : transition
    port map(
      preds      => transition_143_preds,
      symbol_out => transition_143_symbol_out,
      symbol_in  => LambdaIn(38));

  transition_144_preds(0) <= place_147_token;
  LambdaOut(39) <= transition_144_symbol_out;
  transition_144 : transition
    port map(
      preds      => transition_144_preds,
      symbol_out => transition_144_symbol_out,
      symbol_in  => true);

  transition_145_preds(0) <= place_148_token;
  transition_145 : transition
    port map(
      preds      => transition_145_preds,
      symbol_out => transition_145_symbol_out,
      symbol_in  => LambdaIn(39));

  transition_149_preds(0) <= place_1083_token;
  LambdaOut(40) <= transition_149_symbol_out;
  transition_149 : transition
    port map(
      preds      => transition_149_preds,
      symbol_out => transition_149_symbol_out,
      symbol_in  => true);

  transition_150_preds(0) <= place_153_token;
  transition_150 : transition
    port map(
      preds      => transition_150_preds,
      symbol_out => transition_150_symbol_out,
      symbol_in  => LambdaIn(40));

  transition_151_preds(0) <= place_154_token;
  LambdaOut(41) <= transition_151_symbol_out;
  transition_151 : transition
    port map(
      preds      => transition_151_preds,
      symbol_out => transition_151_symbol_out,
      symbol_in  => true);

  transition_152_preds(0) <= place_155_token;
  transition_152 : transition
    port map(
      preds      => transition_152_preds,
      symbol_out => transition_152_symbol_out,
      symbol_in  => LambdaIn(41));

  transition_156_preds(0) <= place_1084_token;
  LambdaOut(42) <= transition_156_symbol_out;
  transition_156 : transition
    port map(
      preds      => transition_156_preds,
      symbol_out => transition_156_symbol_out,
      symbol_in  => true);

  transition_157_preds(0) <= place_160_token;
  transition_157 : transition
    port map(
      preds      => transition_157_preds,
      symbol_out => transition_157_symbol_out,
      symbol_in  => LambdaIn(42));

  transition_158_preds(0) <= place_161_token;
  LambdaOut(43) <= transition_158_symbol_out;
  transition_158 : transition
    port map(
      preds      => transition_158_preds,
      symbol_out => transition_158_symbol_out,
      symbol_in  => true);

  transition_159_preds(0) <= place_162_token;
  transition_159 : transition
    port map(
      preds      => transition_159_preds,
      symbol_out => transition_159_symbol_out,
      symbol_in  => LambdaIn(43));

  transition_163_preds(0) <= place_1082_token;
  transition_163_preds(1) <= place_1385_token;
  transition_163 : transition
    port map(
      preds      => transition_163_preds,
      symbol_out => transition_163_symbol_out,
      symbol_in  => true);

  transition_164_preds(0) <= place_1085_token;
  transition_164 : transition
    port map(
      preds      => transition_164_preds,
      symbol_out => transition_164_symbol_out,
      symbol_in  => true);

  transition_166_preds(0) <= place_165_token;
  transition_166 : transition
    port map(
      preds      => transition_166_preds,
      symbol_out => transition_166_symbol_out,
      symbol_in  => LambdaIn(44));

  transition_167_preds(0) <= place_1086_token;
  LambdaOut(44) <= transition_167_symbol_out;
  transition_167 : transition
    port map(
      preds      => transition_167_preds,
      symbol_out => transition_167_symbol_out,
      symbol_in  => true);

  transition_168_preds(0) <= place_1089_token;
  transition_168_preds(1) <= place_1090_token;
  transition_168_preds(2) <= place_1269_token;
  transition_168 : transition
    port map(
      preds      => transition_168_preds,
      symbol_out => transition_168_symbol_out,
      symbol_in  => true);

  transition_169_preds(0) <= place_1092_token;
  LambdaOut(45) <= transition_169_symbol_out;
  transition_169 : transition
    port map(
      preds      => transition_169_preds,
      symbol_out => transition_169_symbol_out,
      symbol_in  => true);

  transition_170_preds(0) <= place_173_token;
  transition_170 : transition
    port map(
      preds      => transition_170_preds,
      symbol_out => transition_170_symbol_out,
      symbol_in  => LambdaIn(45));

  transition_171_preds(0) <= place_174_token;
  LambdaOut(46) <= transition_171_symbol_out;
  transition_171 : transition
    port map(
      preds      => transition_171_preds,
      symbol_out => transition_171_symbol_out,
      symbol_in  => true);

  transition_172_preds(0) <= place_175_token;
  transition_172 : transition
    port map(
      preds      => transition_172_preds,
      symbol_out => transition_172_symbol_out,
      symbol_in  => LambdaIn(46));

  transition_176_preds(0) <= place_1095_token;
  LambdaOut(47) <= transition_176_symbol_out;
  transition_176 : transition
    port map(
      preds      => transition_176_preds,
      symbol_out => transition_176_symbol_out,
      symbol_in  => true);

  transition_177_preds(0) <= place_180_token;
  transition_177 : transition
    port map(
      preds      => transition_177_preds,
      symbol_out => transition_177_symbol_out,
      symbol_in  => LambdaIn(47));

  transition_178_preds(0) <= place_181_token;
  LambdaOut(48) <= transition_178_symbol_out;
  transition_178 : transition
    port map(
      preds      => transition_178_preds,
      symbol_out => transition_178_symbol_out,
      symbol_in  => true);

  transition_179_preds(0) <= place_182_token;
  transition_179 : transition
    port map(
      preds      => transition_179_preds,
      symbol_out => transition_179_symbol_out,
      symbol_in  => LambdaIn(48));

  transition_183_preds(0) <= place_1096_token;
  LambdaOut(49) <= transition_183_symbol_out;
  transition_183 : transition
    port map(
      preds      => transition_183_preds,
      symbol_out => transition_183_symbol_out,
      symbol_in  => true);

  transition_184_preds(0) <= place_187_token;
  transition_184 : transition
    port map(
      preds      => transition_184_preds,
      symbol_out => transition_184_symbol_out,
      symbol_in  => LambdaIn(49));

  transition_185_preds(0) <= place_188_token;
  LambdaOut(50) <= transition_185_symbol_out;
  transition_185 : transition
    port map(
      preds      => transition_185_preds,
      symbol_out => transition_185_symbol_out,
      symbol_in  => true);

  transition_186_preds(0) <= place_189_token;
  transition_186 : transition
    port map(
      preds      => transition_186_preds,
      symbol_out => transition_186_symbol_out,
      symbol_in  => LambdaIn(50));

  transition_190_preds(0) <= place_1091_token;
  transition_190_preds(1) <= place_1093_token;
  transition_190 : transition
    port map(
      preds      => transition_190_preds,
      symbol_out => transition_190_symbol_out,
      symbol_in  => true);

  transition_191_preds(0) <= place_1097_token;
  LambdaOut(51) <= transition_191_symbol_out;
  transition_191 : transition
    port map(
      preds      => transition_191_preds,
      symbol_out => transition_191_symbol_out,
      symbol_in  => true);

  transition_192_preds(0) <= place_195_token;
  transition_192 : transition
    port map(
      preds      => transition_192_preds,
      symbol_out => transition_192_symbol_out,
      symbol_in  => LambdaIn(51));

  transition_193_preds(0) <= place_196_token;
  LambdaOut(52) <= transition_193_symbol_out;
  transition_193 : transition
    port map(
      preds      => transition_193_preds,
      symbol_out => transition_193_symbol_out,
      symbol_in  => true);

  transition_194_preds(0) <= place_197_token;
  transition_194 : transition
    port map(
      preds      => transition_194_preds,
      symbol_out => transition_194_symbol_out,
      symbol_in  => LambdaIn(52));

  transition_198_preds(0) <= place_1100_token;
  LambdaOut(53) <= transition_198_symbol_out;
  transition_198 : transition
    port map(
      preds      => transition_198_preds,
      symbol_out => transition_198_symbol_out,
      symbol_in  => true);

  transition_199_preds(0) <= place_202_token;
  transition_199 : transition
    port map(
      preds      => transition_199_preds,
      symbol_out => transition_199_symbol_out,
      symbol_in  => LambdaIn(53));

  transition_200_preds(0) <= place_203_token;
  LambdaOut(54) <= transition_200_symbol_out;
  transition_200 : transition
    port map(
      preds      => transition_200_preds,
      symbol_out => transition_200_symbol_out,
      symbol_in  => true);

  transition_201_preds(0) <= place_204_token;
  transition_201 : transition
    port map(
      preds      => transition_201_preds,
      symbol_out => transition_201_symbol_out,
      symbol_in  => LambdaIn(54));

  transition_205_preds(0) <= place_1101_token;
  LambdaOut(55) <= transition_205_symbol_out;
  transition_205 : transition
    port map(
      preds      => transition_205_preds,
      symbol_out => transition_205_symbol_out,
      symbol_in  => true);

  transition_206_preds(0) <= place_209_token;
  transition_206 : transition
    port map(
      preds      => transition_206_preds,
      symbol_out => transition_206_symbol_out,
      symbol_in  => LambdaIn(55));

  transition_207_preds(0) <= place_210_token;
  LambdaOut(56) <= transition_207_symbol_out;
  transition_207 : transition
    port map(
      preds      => transition_207_preds,
      symbol_out => transition_207_symbol_out,
      symbol_in  => true);

  transition_208_preds(0) <= place_211_token;
  transition_208 : transition
    port map(
      preds      => transition_208_preds,
      symbol_out => transition_208_symbol_out,
      symbol_in  => LambdaIn(56));

  transition_212_preds(0) <= place_1098_token;
  transition_212_preds(1) <= place_1099_token;
  transition_212 : transition
    port map(
      preds      => transition_212_preds,
      symbol_out => transition_212_symbol_out,
      symbol_in  => true);

  transition_214_preds(0) <= place_213_token;
  transition_214 : transition
    port map(
      preds      => transition_214_preds,
      symbol_out => transition_214_symbol_out,
      symbol_in  => LambdaIn(57));

  transition_215_preds(0) <= place_1104_token;
  LambdaOut(57) <= transition_215_symbol_out;
  transition_215 : transition
    port map(
      preds      => transition_215_preds,
      symbol_out => transition_215_symbol_out,
      symbol_in  => true);

  transition_216_preds(0) <= place_1087_token;
  transition_216_preds(1) <= place_1102_token;
  transition_216_preds(2) <= place_1377_token;
  transition_216 : transition
    port map(
      preds      => transition_216_preds,
      symbol_out => transition_216_symbol_out,
      symbol_in  => true);

  transition_217_preds(0) <= place_1107_token;
  LambdaOut(58) <= transition_217_symbol_out;
  transition_217 : transition
    port map(
      preds      => transition_217_preds,
      symbol_out => transition_217_symbol_out,
      symbol_in  => true);

  transition_218_preds(0) <= place_221_token;
  transition_218 : transition
    port map(
      preds      => transition_218_preds,
      symbol_out => transition_218_symbol_out,
      symbol_in  => LambdaIn(58));

  transition_219_preds(0) <= place_222_token;
  LambdaOut(59) <= transition_219_symbol_out;
  transition_219 : transition
    port map(
      preds      => transition_219_preds,
      symbol_out => transition_219_symbol_out,
      symbol_in  => true);

  transition_220_preds(0) <= place_223_token;
  transition_220 : transition
    port map(
      preds      => transition_220_preds,
      symbol_out => transition_220_symbol_out,
      symbol_in  => LambdaIn(59));

  transition_224_preds(0) <= place_1106_token;
  LambdaOut(60) <= transition_224_symbol_out;
  transition_224 : transition
    port map(
      preds      => transition_224_preds,
      symbol_out => transition_224_symbol_out,
      symbol_in  => true);

  transition_225_preds(0) <= place_228_token;
  transition_225 : transition
    port map(
      preds      => transition_225_preds,
      symbol_out => transition_225_symbol_out,
      symbol_in  => LambdaIn(60));

  transition_226_preds(0) <= place_229_token;
  LambdaOut(61) <= transition_226_symbol_out;
  transition_226 : transition
    port map(
      preds      => transition_226_preds,
      symbol_out => transition_226_symbol_out,
      symbol_in  => true);

  transition_227_preds(0) <= place_230_token;
  transition_227 : transition
    port map(
      preds      => transition_227_preds,
      symbol_out => transition_227_symbol_out,
      symbol_in  => LambdaIn(61));

  transition_231_preds(0) <= place_1110_token;
  transition_231 : transition
    port map(
      preds      => transition_231_preds,
      symbol_out => transition_231_symbol_out,
      symbol_in  => true);

  transition_233_preds(0) <= place_232_token;
  transition_233 : transition
    port map(
      preds      => transition_233_preds,
      symbol_out => transition_233_symbol_out,
      symbol_in  => LambdaIn(62));

  transition_234_preds(0) <= place_1112_token;
  LambdaOut(62) <= transition_234_symbol_out;
  transition_234 : transition
    port map(
      preds      => transition_234_preds,
      symbol_out => transition_234_symbol_out,
      symbol_in  => true);

  transition_235_preds(0) <= place_1114_token;
  LambdaOut(63) <= transition_235_symbol_out;
  transition_235 : transition
    port map(
      preds      => transition_235_preds,
      symbol_out => transition_235_symbol_out,
      symbol_in  => true);

  transition_237_preds(0) <= place_236_token;
  transition_237 : transition
    port map(
      preds      => transition_237_preds,
      symbol_out => transition_237_symbol_out,
      symbol_in  => LambdaIn(63));

  transition_238_preds(0) <= place_1115_token;
  LambdaOut(64) <= transition_238_symbol_out;
  transition_238 : transition
    port map(
      preds      => transition_238_preds,
      symbol_out => transition_238_symbol_out,
      symbol_in  => true);

  transition_239_preds(0) <= place_1117_token;
  LambdaOut(65) <= transition_239_symbol_out;
  transition_239 : transition
    port map(
      preds      => transition_239_preds,
      symbol_out => transition_239_symbol_out,
      symbol_in  => true);

  transition_240_preds(0) <= place_1120_token;
  LambdaOut(66) <= transition_240_symbol_out;
  transition_240 : transition
    port map(
      preds      => transition_240_preds,
      symbol_out => transition_240_symbol_out,
      symbol_in  => true);

  transition_241_preds(0) <= place_244_token;
  transition_241 : transition
    port map(
      preds      => transition_241_preds,
      symbol_out => transition_241_symbol_out,
      symbol_in  => LambdaIn(64));

  transition_242_preds(0) <= place_245_token;
  LambdaOut(67) <= transition_242_symbol_out;
  transition_242 : transition
    port map(
      preds      => transition_242_preds,
      symbol_out => transition_242_symbol_out,
      symbol_in  => true);

  transition_243_preds(0) <= place_246_token;
  transition_243 : transition
    port map(
      preds      => transition_243_preds,
      symbol_out => transition_243_symbol_out,
      symbol_in  => LambdaIn(65));

  transition_247_preds(0) <= place_1122_token;
  LambdaOut(68) <= transition_247_symbol_out;
  transition_247 : transition
    port map(
      preds      => transition_247_preds,
      symbol_out => transition_247_symbol_out,
      symbol_in  => true);

  transition_248_preds(0) <= place_251_token;
  transition_248 : transition
    port map(
      preds      => transition_248_preds,
      symbol_out => transition_248_symbol_out,
      symbol_in  => LambdaIn(66));

  transition_249_preds(0) <= place_252_token;
  LambdaOut(69) <= transition_249_symbol_out;
  transition_249 : transition
    port map(
      preds      => transition_249_preds,
      symbol_out => transition_249_symbol_out,
      symbol_in  => true);

  transition_250_preds(0) <= place_253_token;
  transition_250 : transition
    port map(
      preds      => transition_250_preds,
      symbol_out => transition_250_symbol_out,
      symbol_in  => LambdaIn(67));

  transition_254_preds(0) <= place_1123_token;
  LambdaOut(70) <= transition_254_symbol_out;
  transition_254 : transition
    port map(
      preds      => transition_254_preds,
      symbol_out => transition_254_symbol_out,
      symbol_in  => true);

  transition_255_preds(0) <= place_258_token;
  transition_255 : transition
    port map(
      preds      => transition_255_preds,
      symbol_out => transition_255_symbol_out,
      symbol_in  => LambdaIn(68));

  transition_256_preds(0) <= place_259_token;
  LambdaOut(71) <= transition_256_symbol_out;
  transition_256 : transition
    port map(
      preds      => transition_256_preds,
      symbol_out => transition_256_symbol_out,
      symbol_in  => true);

  transition_257_preds(0) <= place_260_token;
  transition_257 : transition
    port map(
      preds      => transition_257_preds,
      symbol_out => transition_257_symbol_out,
      symbol_in  => LambdaIn(69));

  transition_261_preds(0) <= place_1118_token;
  transition_261_preds(1) <= place_1121_token;
  transition_261 : transition
    port map(
      preds      => transition_261_preds,
      symbol_out => transition_261_symbol_out,
      symbol_in  => true);

  transition_262_preds(0) <= place_1126_token;
  LambdaOut(72) <= transition_262_symbol_out;
  transition_262 : transition
    port map(
      preds      => transition_262_preds,
      symbol_out => transition_262_symbol_out,
      symbol_in  => true);

  transition_263_preds(0) <= place_266_token;
  transition_263 : transition
    port map(
      preds      => transition_263_preds,
      symbol_out => transition_263_symbol_out,
      symbol_in  => LambdaIn(70));

  transition_264_preds(0) <= place_267_token;
  LambdaOut(73) <= transition_264_symbol_out;
  transition_264 : transition
    port map(
      preds      => transition_264_preds,
      symbol_out => transition_264_symbol_out,
      symbol_in  => true);

  transition_265_preds(0) <= place_268_token;
  transition_265 : transition
    port map(
      preds      => transition_265_preds,
      symbol_out => transition_265_symbol_out,
      symbol_in  => LambdaIn(71));

  transition_269_preds(0) <= place_1127_token;
  LambdaOut(74) <= transition_269_symbol_out;
  transition_269 : transition
    port map(
      preds      => transition_269_preds,
      symbol_out => transition_269_symbol_out,
      symbol_in  => true);

  transition_270_preds(0) <= place_273_token;
  transition_270 : transition
    port map(
      preds      => transition_270_preds,
      symbol_out => transition_270_symbol_out,
      symbol_in  => LambdaIn(72));

  transition_271_preds(0) <= place_274_token;
  LambdaOut(75) <= transition_271_symbol_out;
  transition_271 : transition
    port map(
      preds      => transition_271_preds,
      symbol_out => transition_271_symbol_out,
      symbol_in  => true);

  transition_272_preds(0) <= place_275_token;
  transition_272 : transition
    port map(
      preds      => transition_272_preds,
      symbol_out => transition_272_symbol_out,
      symbol_in  => LambdaIn(73));

  transition_276_preds(0) <= place_1124_token;
  transition_276_preds(1) <= place_1125_token;
  transition_276 : transition
    port map(
      preds      => transition_276_preds,
      symbol_out => transition_276_symbol_out,
      symbol_in  => true);

  transition_277_preds(0) <= place_1128_token;
  LambdaOut(76) <= transition_277_symbol_out;
  transition_277 : transition
    port map(
      preds      => transition_277_preds,
      symbol_out => transition_277_symbol_out,
      symbol_in  => true);

  transition_278_preds(0) <= place_281_token;
  transition_278 : transition
    port map(
      preds      => transition_278_preds,
      symbol_out => transition_278_symbol_out,
      symbol_in  => LambdaIn(74));

  transition_279_preds(0) <= place_282_token;
  LambdaOut(77) <= transition_279_symbol_out;
  transition_279 : transition
    port map(
      preds      => transition_279_preds,
      symbol_out => transition_279_symbol_out,
      symbol_in  => true);

  transition_280_preds(0) <= place_283_token;
  transition_280 : transition
    port map(
      preds      => transition_280_preds,
      symbol_out => transition_280_symbol_out,
      symbol_in  => LambdaIn(75));

  transition_284_preds(0) <= place_1134_token;
  LambdaOut(78) <= transition_284_symbol_out;
  transition_284 : transition
    port map(
      preds      => transition_284_preds,
      symbol_out => transition_284_symbol_out,
      symbol_in  => true);

  transition_285_preds(0) <= place_288_token;
  transition_285 : transition
    port map(
      preds      => transition_285_preds,
      symbol_out => transition_285_symbol_out,
      symbol_in  => LambdaIn(76));

  transition_286_preds(0) <= place_289_token;
  LambdaOut(79) <= transition_286_symbol_out;
  transition_286 : transition
    port map(
      preds      => transition_286_preds,
      symbol_out => transition_286_symbol_out,
      symbol_in  => true);

  transition_287_preds(0) <= place_290_token;
  transition_287 : transition
    port map(
      preds      => transition_287_preds,
      symbol_out => transition_287_symbol_out,
      symbol_in  => LambdaIn(77));

  transition_291_preds(0) <= place_1136_token;
  LambdaOut(80) <= transition_291_symbol_out;
  transition_291 : transition
    port map(
      preds      => transition_291_preds,
      symbol_out => transition_291_symbol_out,
      symbol_in  => true);

  transition_292_preds(0) <= place_295_token;
  transition_292 : transition
    port map(
      preds      => transition_292_preds,
      symbol_out => transition_292_symbol_out,
      symbol_in  => LambdaIn(78));

  transition_293_preds(0) <= place_296_token;
  LambdaOut(81) <= transition_293_symbol_out;
  transition_293 : transition
    port map(
      preds      => transition_293_preds,
      symbol_out => transition_293_symbol_out,
      symbol_in  => true);

  transition_294_preds(0) <= place_297_token;
  transition_294 : transition
    port map(
      preds      => transition_294_preds,
      symbol_out => transition_294_symbol_out,
      symbol_in  => LambdaIn(79));

  transition_298_preds(0) <= place_1137_token;
  LambdaOut(82) <= transition_298_symbol_out;
  transition_298 : transition
    port map(
      preds      => transition_298_preds,
      symbol_out => transition_298_symbol_out,
      symbol_in  => true);

  transition_299_preds(0) <= place_302_token;
  transition_299 : transition
    port map(
      preds      => transition_299_preds,
      symbol_out => transition_299_symbol_out,
      symbol_in  => LambdaIn(80));

  transition_300_preds(0) <= place_303_token;
  LambdaOut(83) <= transition_300_symbol_out;
  transition_300 : transition
    port map(
      preds      => transition_300_preds,
      symbol_out => transition_300_symbol_out,
      symbol_in  => true);

  transition_301_preds(0) <= place_304_token;
  transition_301 : transition
    port map(
      preds      => transition_301_preds,
      symbol_out => transition_301_symbol_out,
      symbol_in  => LambdaIn(81));

  transition_305_preds(0) <= place_1131_token;
  transition_305_preds(1) <= place_1135_token;
  transition_305 : transition
    port map(
      preds      => transition_305_preds,
      symbol_out => transition_305_symbol_out,
      symbol_in  => true);

  transition_306_preds(0) <= place_1140_token;
  LambdaOut(84) <= transition_306_symbol_out;
  transition_306 : transition
    port map(
      preds      => transition_306_preds,
      symbol_out => transition_306_symbol_out,
      symbol_in  => true);

  transition_307_preds(0) <= place_310_token;
  transition_307 : transition
    port map(
      preds      => transition_307_preds,
      symbol_out => transition_307_symbol_out,
      symbol_in  => LambdaIn(82));

  transition_308_preds(0) <= place_311_token;
  LambdaOut(85) <= transition_308_symbol_out;
  transition_308 : transition
    port map(
      preds      => transition_308_preds,
      symbol_out => transition_308_symbol_out,
      symbol_in  => true);

  transition_309_preds(0) <= place_312_token;
  transition_309 : transition
    port map(
      preds      => transition_309_preds,
      symbol_out => transition_309_symbol_out,
      symbol_in  => LambdaIn(83));

  transition_313_preds(0) <= place_1141_token;
  LambdaOut(86) <= transition_313_symbol_out;
  transition_313 : transition
    port map(
      preds      => transition_313_preds,
      symbol_out => transition_313_symbol_out,
      symbol_in  => true);

  transition_314_preds(0) <= place_317_token;
  transition_314 : transition
    port map(
      preds      => transition_314_preds,
      symbol_out => transition_314_symbol_out,
      symbol_in  => LambdaIn(84));

  transition_315_preds(0) <= place_318_token;
  LambdaOut(87) <= transition_315_symbol_out;
  transition_315 : transition
    port map(
      preds      => transition_315_preds,
      symbol_out => transition_315_symbol_out,
      symbol_in  => true);

  transition_316_preds(0) <= place_319_token;
  transition_316 : transition
    port map(
      preds      => transition_316_preds,
      symbol_out => transition_316_symbol_out,
      symbol_in  => LambdaIn(85));

  transition_320_preds(0) <= place_1138_token;
  transition_320_preds(1) <= place_1139_token;
  transition_320 : transition
    port map(
      preds      => transition_320_preds,
      symbol_out => transition_320_symbol_out,
      symbol_in  => true);

  transition_321_preds(0) <= place_1142_token;
  LambdaOut(88) <= transition_321_symbol_out;
  transition_321 : transition
    port map(
      preds      => transition_321_preds,
      symbol_out => transition_321_symbol_out,
      symbol_in  => true);

  transition_322_preds(0) <= place_325_token;
  transition_322 : transition
    port map(
      preds      => transition_322_preds,
      symbol_out => transition_322_symbol_out,
      symbol_in  => LambdaIn(86));

  transition_323_preds(0) <= place_326_token;
  LambdaOut(89) <= transition_323_symbol_out;
  transition_323 : transition
    port map(
      preds      => transition_323_preds,
      symbol_out => transition_323_symbol_out,
      symbol_in  => true);

  transition_324_preds(0) <= place_327_token;
  transition_324 : transition
    port map(
      preds      => transition_324_preds,
      symbol_out => transition_324_symbol_out,
      symbol_in  => LambdaIn(87));

  transition_328_preds(0) <= place_1146_token;
  LambdaOut(90) <= transition_328_symbol_out;
  transition_328 : transition
    port map(
      preds      => transition_328_preds,
      symbol_out => transition_328_symbol_out,
      symbol_in  => true);

  transition_329_preds(0) <= place_332_token;
  transition_329 : transition
    port map(
      preds      => transition_329_preds,
      symbol_out => transition_329_symbol_out,
      symbol_in  => LambdaIn(88));

  transition_330_preds(0) <= place_333_token;
  LambdaOut(91) <= transition_330_symbol_out;
  transition_330 : transition
    port map(
      preds      => transition_330_preds,
      symbol_out => transition_330_symbol_out,
      symbol_in  => true);

  transition_331_preds(0) <= place_334_token;
  transition_331 : transition
    port map(
      preds      => transition_331_preds,
      symbol_out => transition_331_symbol_out,
      symbol_in  => LambdaIn(89));

  transition_335_preds(0) <= place_1148_token;
  LambdaOut(92) <= transition_335_symbol_out;
  transition_335 : transition
    port map(
      preds      => transition_335_preds,
      symbol_out => transition_335_symbol_out,
      symbol_in  => true);

  transition_336_preds(0) <= place_339_token;
  transition_336 : transition
    port map(
      preds      => transition_336_preds,
      symbol_out => transition_336_symbol_out,
      symbol_in  => LambdaIn(90));

  transition_337_preds(0) <= place_340_token;
  LambdaOut(93) <= transition_337_symbol_out;
  transition_337 : transition
    port map(
      preds      => transition_337_preds,
      symbol_out => transition_337_symbol_out,
      symbol_in  => true);

  transition_338_preds(0) <= place_341_token;
  transition_338 : transition
    port map(
      preds      => transition_338_preds,
      symbol_out => transition_338_symbol_out,
      symbol_in  => LambdaIn(91));

  transition_342_preds(0) <= place_1149_token;
  LambdaOut(94) <= transition_342_symbol_out;
  transition_342 : transition
    port map(
      preds      => transition_342_preds,
      symbol_out => transition_342_symbol_out,
      symbol_in  => true);

  transition_343_preds(0) <= place_346_token;
  transition_343 : transition
    port map(
      preds      => transition_343_preds,
      symbol_out => transition_343_symbol_out,
      symbol_in  => LambdaIn(92));

  transition_344_preds(0) <= place_347_token;
  LambdaOut(95) <= transition_344_symbol_out;
  transition_344 : transition
    port map(
      preds      => transition_344_preds,
      symbol_out => transition_344_symbol_out,
      symbol_in  => true);

  transition_345_preds(0) <= place_348_token;
  transition_345 : transition
    port map(
      preds      => transition_345_preds,
      symbol_out => transition_345_symbol_out,
      symbol_in  => LambdaIn(93));

  transition_349_preds(0) <= place_1145_token;
  transition_349_preds(1) <= place_1147_token;
  transition_349 : transition
    port map(
      preds      => transition_349_preds,
      symbol_out => transition_349_symbol_out,
      symbol_in  => true);

  transition_350_preds(0) <= place_1150_token;
  LambdaOut(96) <= transition_350_symbol_out;
  transition_350 : transition
    port map(
      preds      => transition_350_preds,
      symbol_out => transition_350_symbol_out,
      symbol_in  => true);

  transition_351_preds(0) <= place_354_token;
  transition_351 : transition
    port map(
      preds      => transition_351_preds,
      symbol_out => transition_351_symbol_out,
      symbol_in  => LambdaIn(94));

  transition_352_preds(0) <= place_355_token;
  LambdaOut(97) <= transition_352_symbol_out;
  transition_352 : transition
    port map(
      preds      => transition_352_preds,
      symbol_out => transition_352_symbol_out,
      symbol_in  => true);

  transition_353_preds(0) <= place_356_token;
  transition_353 : transition
    port map(
      preds      => transition_353_preds,
      symbol_out => transition_353_symbol_out,
      symbol_in  => LambdaIn(95));

  transition_357_preds(0) <= place_1154_token;
  LambdaOut(98) <= transition_357_symbol_out;
  transition_357 : transition
    port map(
      preds      => transition_357_preds,
      symbol_out => transition_357_symbol_out,
      symbol_in  => true);

  transition_358_preds(0) <= place_361_token;
  transition_358 : transition
    port map(
      preds      => transition_358_preds,
      symbol_out => transition_358_symbol_out,
      symbol_in  => LambdaIn(96));

  transition_359_preds(0) <= place_362_token;
  LambdaOut(99) <= transition_359_symbol_out;
  transition_359 : transition
    port map(
      preds      => transition_359_preds,
      symbol_out => transition_359_symbol_out,
      symbol_in  => true);

  transition_360_preds(0) <= place_363_token;
  transition_360 : transition
    port map(
      preds      => transition_360_preds,
      symbol_out => transition_360_symbol_out,
      symbol_in  => LambdaIn(97));

  transition_364_preds(0) <= place_1155_token;
  LambdaOut(100) <= transition_364_symbol_out;
  transition_364 : transition
    port map(
      preds      => transition_364_preds,
      symbol_out => transition_364_symbol_out,
      symbol_in  => true);

  transition_365_preds(0) <= place_368_token;
  transition_365 : transition
    port map(
      preds      => transition_365_preds,
      symbol_out => transition_365_symbol_out,
      symbol_in  => LambdaIn(98));

  transition_366_preds(0) <= place_369_token;
  LambdaOut(101) <= transition_366_symbol_out;
  transition_366 : transition
    port map(
      preds      => transition_366_preds,
      symbol_out => transition_366_symbol_out,
      symbol_in  => true);

  transition_367_preds(0) <= place_370_token;
  transition_367 : transition
    port map(
      preds      => transition_367_preds,
      symbol_out => transition_367_symbol_out,
      symbol_in  => LambdaIn(99));

  transition_371_preds(0) <= place_1153_token;
  transition_371_preds(1) <= place_1151_token;
  transition_371 : transition
    port map(
      preds      => transition_371_preds,
      symbol_out => transition_371_symbol_out,
      symbol_in  => true);

  transition_372_preds(0) <= place_1156_token;
  transition_372 : transition
    port map(
      preds      => transition_372_preds,
      symbol_out => transition_372_symbol_out,
      symbol_in  => true);

  transition_373_preds(0) <= place_1158_token;
  LambdaOut(102) <= transition_373_symbol_out;
  transition_373 : transition
    port map(
      preds      => transition_373_preds,
      symbol_out => transition_373_symbol_out,
      symbol_in  => true);

  transition_374_preds(0) <= place_377_token;
  transition_374 : transition
    port map(
      preds      => transition_374_preds,
      symbol_out => transition_374_symbol_out,
      symbol_in  => LambdaIn(100));

  transition_375_preds(0) <= place_378_token;
  LambdaOut(103) <= transition_375_symbol_out;
  transition_375 : transition
    port map(
      preds      => transition_375_preds,
      symbol_out => transition_375_symbol_out,
      symbol_in  => true);

  transition_376_preds(0) <= place_379_token;
  transition_376 : transition
    port map(
      preds      => transition_376_preds,
      symbol_out => transition_376_symbol_out,
      symbol_in  => LambdaIn(101));

  transition_381_preds(0) <= place_380_token;
  transition_381 : transition
    port map(
      preds      => transition_381_preds,
      symbol_out => transition_381_symbol_out,
      symbol_in  => LambdaIn(102));

  transition_382_preds(0) <= place_1159_token;
  LambdaOut(104) <= transition_382_symbol_out;
  transition_382 : transition
    port map(
      preds      => transition_382_preds,
      symbol_out => transition_382_symbol_out,
      symbol_in  => true);

  transition_383_preds(0) <= place_1130_token;
  transition_383_preds(1) <= place_1157_token;
  transition_383_preds(2) <= place_1161_token;
  transition_383 : transition
    port map(
      preds      => transition_383_preds,
      symbol_out => transition_383_symbol_out,
      symbol_in  => true);

  transition_384_preds(0) <= place_1163_token;
  LambdaOut(105) <= transition_384_symbol_out;
  transition_384 : transition
    port map(
      preds      => transition_384_preds,
      symbol_out => transition_384_symbol_out,
      symbol_in  => true);

  transition_385_preds(0) <= place_388_token;
  transition_385 : transition
    port map(
      preds      => transition_385_preds,
      symbol_out => transition_385_symbol_out,
      symbol_in  => LambdaIn(103));

  transition_386_preds(0) <= place_389_token;
  LambdaOut(106) <= transition_386_symbol_out;
  transition_386 : transition
    port map(
      preds      => transition_386_preds,
      symbol_out => transition_386_symbol_out,
      symbol_in  => true);

  transition_387_preds(0) <= place_390_token;
  transition_387 : transition
    port map(
      preds      => transition_387_preds,
      symbol_out => transition_387_symbol_out,
      symbol_in  => LambdaIn(104));

  transition_391_preds(0) <= place_1165_token;
  LambdaOut(107) <= transition_391_symbol_out;
  transition_391 : transition
    port map(
      preds      => transition_391_preds,
      symbol_out => transition_391_symbol_out,
      symbol_in  => true);

  transition_392_preds(0) <= place_395_token;
  transition_392 : transition
    port map(
      preds      => transition_392_preds,
      symbol_out => transition_392_symbol_out,
      symbol_in  => LambdaIn(105));

  transition_393_preds(0) <= place_396_token;
  LambdaOut(108) <= transition_393_symbol_out;
  transition_393 : transition
    port map(
      preds      => transition_393_preds,
      symbol_out => transition_393_symbol_out,
      symbol_in  => true);

  transition_394_preds(0) <= place_397_token;
  transition_394 : transition
    port map(
      preds      => transition_394_preds,
      symbol_out => transition_394_symbol_out,
      symbol_in  => LambdaIn(106));

  transition_398_preds(0) <= place_1166_token;
  LambdaOut(109) <= transition_398_symbol_out;
  transition_398 : transition
    port map(
      preds      => transition_398_preds,
      symbol_out => transition_398_symbol_out,
      symbol_in  => true);

  transition_399_preds(0) <= place_402_token;
  transition_399 : transition
    port map(
      preds      => transition_399_preds,
      symbol_out => transition_399_symbol_out,
      symbol_in  => LambdaIn(107));

  transition_400_preds(0) <= place_403_token;
  LambdaOut(110) <= transition_400_symbol_out;
  transition_400 : transition
    port map(
      preds      => transition_400_preds,
      symbol_out => transition_400_symbol_out,
      symbol_in  => true);

  transition_401_preds(0) <= place_404_token;
  transition_401 : transition
    port map(
      preds      => transition_401_preds,
      symbol_out => transition_401_symbol_out,
      symbol_in  => LambdaIn(108));

  transition_405_preds(0) <= place_1162_token;
  transition_405_preds(1) <= place_1164_token;
  transition_405 : transition
    port map(
      preds      => transition_405_preds,
      symbol_out => transition_405_symbol_out,
      symbol_in  => true);

  transition_406_preds(0) <= place_1167_token;
  LambdaOut(111) <= transition_406_symbol_out;
  transition_406 : transition
    port map(
      preds      => transition_406_preds,
      symbol_out => transition_406_symbol_out,
      symbol_in  => true);

  transition_407_preds(0) <= place_410_token;
  transition_407 : transition
    port map(
      preds      => transition_407_preds,
      symbol_out => transition_407_symbol_out,
      symbol_in  => LambdaIn(109));

  transition_408_preds(0) <= place_411_token;
  LambdaOut(112) <= transition_408_symbol_out;
  transition_408 : transition
    port map(
      preds      => transition_408_preds,
      symbol_out => transition_408_symbol_out,
      symbol_in  => true);

  transition_409_preds(0) <= place_412_token;
  transition_409 : transition
    port map(
      preds      => transition_409_preds,
      symbol_out => transition_409_symbol_out,
      symbol_in  => LambdaIn(110));

  transition_413_preds(0) <= place_1171_token;
  LambdaOut(113) <= transition_413_symbol_out;
  transition_413 : transition
    port map(
      preds      => transition_413_preds,
      symbol_out => transition_413_symbol_out,
      symbol_in  => true);

  transition_414_preds(0) <= place_417_token;
  transition_414 : transition
    port map(
      preds      => transition_414_preds,
      symbol_out => transition_414_symbol_out,
      symbol_in  => LambdaIn(111));

  transition_415_preds(0) <= place_418_token;
  LambdaOut(114) <= transition_415_symbol_out;
  transition_415 : transition
    port map(
      preds      => transition_415_preds,
      symbol_out => transition_415_symbol_out,
      symbol_in  => true);

  transition_416_preds(0) <= place_419_token;
  transition_416 : transition
    port map(
      preds      => transition_416_preds,
      symbol_out => transition_416_symbol_out,
      symbol_in  => LambdaIn(112));

  transition_420_preds(0) <= place_1172_token;
  LambdaOut(115) <= transition_420_symbol_out;
  transition_420 : transition
    port map(
      preds      => transition_420_preds,
      symbol_out => transition_420_symbol_out,
      symbol_in  => true);

  transition_421_preds(0) <= place_424_token;
  transition_421 : transition
    port map(
      preds      => transition_421_preds,
      symbol_out => transition_421_symbol_out,
      symbol_in  => LambdaIn(113));

  transition_422_preds(0) <= place_425_token;
  LambdaOut(116) <= transition_422_symbol_out;
  transition_422 : transition
    port map(
      preds      => transition_422_preds,
      symbol_out => transition_422_symbol_out,
      symbol_in  => true);

  transition_423_preds(0) <= place_426_token;
  transition_423 : transition
    port map(
      preds      => transition_423_preds,
      symbol_out => transition_423_symbol_out,
      symbol_in  => LambdaIn(114));

  transition_427_preds(0) <= place_1169_token;
  transition_427_preds(1) <= place_1170_token;
  transition_427 : transition
    port map(
      preds      => transition_427_preds,
      symbol_out => transition_427_symbol_out,
      symbol_in  => true);

  transition_428_preds(0) <= place_1173_token;
  LambdaOut(117) <= transition_428_symbol_out;
  transition_428 : transition
    port map(
      preds      => transition_428_preds,
      symbol_out => transition_428_symbol_out,
      symbol_in  => true);

  transition_429_preds(0) <= place_432_token;
  transition_429 : transition
    port map(
      preds      => transition_429_preds,
      symbol_out => transition_429_symbol_out,
      symbol_in  => LambdaIn(115));

  transition_430_preds(0) <= place_433_token;
  LambdaOut(118) <= transition_430_symbol_out;
  transition_430 : transition
    port map(
      preds      => transition_430_preds,
      symbol_out => transition_430_symbol_out,
      symbol_in  => true);

  transition_431_preds(0) <= place_434_token;
  transition_431 : transition
    port map(
      preds      => transition_431_preds,
      symbol_out => transition_431_symbol_out,
      symbol_in  => LambdaIn(116));

  transition_436_preds(0) <= place_435_token;
  transition_436 : transition
    port map(
      preds      => transition_436_preds,
      symbol_out => transition_436_symbol_out,
      symbol_in  => LambdaIn(117));

  transition_437_preds(0) <= place_1175_token;
  LambdaOut(119) <= transition_437_symbol_out;
  transition_437 : transition
    port map(
      preds      => transition_437_preds,
      symbol_out => transition_437_symbol_out,
      symbol_in  => true);

  transition_438_preds(0) <= place_1144_token;
  transition_438_preds(1) <= place_1160_token;
  transition_438_preds(2) <= place_1174_token;
  transition_438 : transition
    port map(
      preds      => transition_438_preds,
      symbol_out => transition_438_symbol_out,
      symbol_in  => true);

  transition_439_preds(0) <= place_1179_token;
  LambdaOut(120) <= transition_439_symbol_out;
  transition_439 : transition
    port map(
      preds      => transition_439_preds,
      symbol_out => transition_439_symbol_out,
      symbol_in  => true);

  transition_440_preds(0) <= place_443_token;
  transition_440 : transition
    port map(
      preds      => transition_440_preds,
      symbol_out => transition_440_symbol_out,
      symbol_in  => LambdaIn(118));

  transition_441_preds(0) <= place_444_token;
  LambdaOut(121) <= transition_441_symbol_out;
  transition_441 : transition
    port map(
      preds      => transition_441_preds,
      symbol_out => transition_441_symbol_out,
      symbol_in  => true);

  transition_442_preds(0) <= place_445_token;
  transition_442 : transition
    port map(
      preds      => transition_442_preds,
      symbol_out => transition_442_symbol_out,
      symbol_in  => LambdaIn(119));

  transition_446_preds(0) <= place_1178_token;
  LambdaOut(122) <= transition_446_symbol_out;
  transition_446 : transition
    port map(
      preds      => transition_446_preds,
      symbol_out => transition_446_symbol_out,
      symbol_in  => true);

  transition_447_preds(0) <= place_450_token;
  transition_447 : transition
    port map(
      preds      => transition_447_preds,
      symbol_out => transition_447_symbol_out,
      symbol_in  => LambdaIn(120));

  transition_448_preds(0) <= place_451_token;
  LambdaOut(123) <= transition_448_symbol_out;
  transition_448 : transition
    port map(
      preds      => transition_448_preds,
      symbol_out => transition_448_symbol_out,
      symbol_in  => true);

  transition_449_preds(0) <= place_452_token;
  transition_449 : transition
    port map(
      preds      => transition_449_preds,
      symbol_out => transition_449_symbol_out,
      symbol_in  => LambdaIn(121));

  transition_453_preds(0) <= place_1183_token;
  LambdaOut(124) <= transition_453_symbol_out;
  transition_453 : transition
    port map(
      preds      => transition_453_preds,
      symbol_out => transition_453_symbol_out,
      symbol_in  => true);

  transition_454_preds(0) <= place_457_token;
  transition_454 : transition
    port map(
      preds      => transition_454_preds,
      symbol_out => transition_454_symbol_out,
      symbol_in  => LambdaIn(122));

  transition_455_preds(0) <= place_458_token;
  LambdaOut(125) <= transition_455_symbol_out;
  transition_455 : transition
    port map(
      preds      => transition_455_preds,
      symbol_out => transition_455_symbol_out,
      symbol_in  => true);

  transition_456_preds(0) <= place_459_token;
  transition_456 : transition
    port map(
      preds      => transition_456_preds,
      symbol_out => transition_456_symbol_out,
      symbol_in  => LambdaIn(123));

  transition_460_preds(0) <= place_1185_token;
  LambdaOut(126) <= transition_460_symbol_out;
  transition_460 : transition
    port map(
      preds      => transition_460_preds,
      symbol_out => transition_460_symbol_out,
      symbol_in  => true);

  transition_461_preds(0) <= place_464_token;
  transition_461 : transition
    port map(
      preds      => transition_461_preds,
      symbol_out => transition_461_symbol_out,
      symbol_in  => LambdaIn(124));

  transition_462_preds(0) <= place_465_token;
  LambdaOut(127) <= transition_462_symbol_out;
  transition_462 : transition
    port map(
      preds      => transition_462_preds,
      symbol_out => transition_462_symbol_out,
      symbol_in  => true);

  transition_463_preds(0) <= place_466_token;
  transition_463 : transition
    port map(
      preds      => transition_463_preds,
      symbol_out => transition_463_symbol_out,
      symbol_in  => LambdaIn(125));

  transition_467_preds(0) <= place_1186_token;
  LambdaOut(128) <= transition_467_symbol_out;
  transition_467 : transition
    port map(
      preds      => transition_467_preds,
      symbol_out => transition_467_symbol_out,
      symbol_in  => true);

  transition_468_preds(0) <= place_471_token;
  transition_468 : transition
    port map(
      preds      => transition_468_preds,
      symbol_out => transition_468_symbol_out,
      symbol_in  => LambdaIn(126));

  transition_469_preds(0) <= place_472_token;
  LambdaOut(129) <= transition_469_symbol_out;
  transition_469 : transition
    port map(
      preds      => transition_469_preds,
      symbol_out => transition_469_symbol_out,
      symbol_in  => true);

  transition_470_preds(0) <= place_473_token;
  transition_470 : transition
    port map(
      preds      => transition_470_preds,
      symbol_out => transition_470_symbol_out,
      symbol_in  => LambdaIn(127));

  transition_474_preds(0) <= place_1184_token;
  transition_474_preds(1) <= place_1182_token;
  transition_474 : transition
    port map(
      preds      => transition_474_preds,
      symbol_out => transition_474_symbol_out,
      symbol_in  => true);

  transition_475_preds(0) <= place_1190_token;
  LambdaOut(130) <= transition_475_symbol_out;
  transition_475 : transition
    port map(
      preds      => transition_475_preds,
      symbol_out => transition_475_symbol_out,
      symbol_in  => true);

  transition_476_preds(0) <= place_479_token;
  transition_476 : transition
    port map(
      preds      => transition_476_preds,
      symbol_out => transition_476_symbol_out,
      symbol_in  => LambdaIn(128));

  transition_477_preds(0) <= place_480_token;
  LambdaOut(131) <= transition_477_symbol_out;
  transition_477 : transition
    port map(
      preds      => transition_477_preds,
      symbol_out => transition_477_symbol_out,
      symbol_in  => true);

  transition_478_preds(0) <= place_481_token;
  transition_478 : transition
    port map(
      preds      => transition_478_preds,
      symbol_out => transition_478_symbol_out,
      symbol_in  => LambdaIn(129));

  transition_482_preds(0) <= place_1191_token;
  LambdaOut(132) <= transition_482_symbol_out;
  transition_482 : transition
    port map(
      preds      => transition_482_preds,
      symbol_out => transition_482_symbol_out,
      symbol_in  => true);

  transition_483_preds(0) <= place_486_token;
  transition_483 : transition
    port map(
      preds      => transition_483_preds,
      symbol_out => transition_483_symbol_out,
      symbol_in  => LambdaIn(130));

  transition_484_preds(0) <= place_487_token;
  LambdaOut(133) <= transition_484_symbol_out;
  transition_484 : transition
    port map(
      preds      => transition_484_preds,
      symbol_out => transition_484_symbol_out,
      symbol_in  => true);

  transition_485_preds(0) <= place_488_token;
  transition_485 : transition
    port map(
      preds      => transition_485_preds,
      symbol_out => transition_485_symbol_out,
      symbol_in  => LambdaIn(131));

  transition_489_preds(0) <= place_1187_token;
  transition_489_preds(1) <= place_1188_token;
  transition_489 : transition
    port map(
      preds      => transition_489_preds,
      symbol_out => transition_489_symbol_out,
      symbol_in  => true);

  transition_490_preds(0) <= place_1192_token;
  LambdaOut(134) <= transition_490_symbol_out;
  transition_490 : transition
    port map(
      preds      => transition_490_preds,
      symbol_out => transition_490_symbol_out,
      symbol_in  => true);

  transition_491_preds(0) <= place_494_token;
  transition_491 : transition
    port map(
      preds      => transition_491_preds,
      symbol_out => transition_491_symbol_out,
      symbol_in  => LambdaIn(132));

  transition_492_preds(0) <= place_495_token;
  LambdaOut(135) <= transition_492_symbol_out;
  transition_492 : transition
    port map(
      preds      => transition_492_preds,
      symbol_out => transition_492_symbol_out,
      symbol_in  => true);

  transition_493_preds(0) <= place_496_token;
  transition_493 : transition
    port map(
      preds      => transition_493_preds,
      symbol_out => transition_493_symbol_out,
      symbol_in  => LambdaIn(133));

  transition_498_preds(0) <= place_497_token;
  transition_498 : transition
    port map(
      preds      => transition_498_preds,
      symbol_out => transition_498_symbol_out,
      symbol_in  => LambdaIn(134));

  transition_499_preds(0) <= place_1195_token;
  LambdaOut(136) <= transition_499_symbol_out;
  transition_499 : transition
    port map(
      preds      => transition_499_preds,
      symbol_out => transition_499_symbol_out,
      symbol_in  => true);

  transition_500_preds(0) <= place_1193_token;
  transition_500_preds(1) <= place_1197_token;
  transition_500 : transition
    port map(
      preds      => transition_500_preds,
      symbol_out => transition_500_symbol_out,
      symbol_in  => true);

  transition_501_preds(0) <= place_1199_token;
  LambdaOut(137) <= transition_501_symbol_out;
  transition_501 : transition
    port map(
      preds      => transition_501_preds,
      symbol_out => transition_501_symbol_out,
      symbol_in  => true);

  transition_502_preds(0) <= place_505_token;
  transition_502 : transition
    port map(
      preds      => transition_502_preds,
      symbol_out => transition_502_symbol_out,
      symbol_in  => LambdaIn(135));

  transition_503_preds(0) <= place_506_token;
  LambdaOut(138) <= transition_503_symbol_out;
  transition_503 : transition
    port map(
      preds      => transition_503_preds,
      symbol_out => transition_503_symbol_out,
      symbol_in  => true);

  transition_504_preds(0) <= place_507_token;
  transition_504 : transition
    port map(
      preds      => transition_504_preds,
      symbol_out => transition_504_symbol_out,
      symbol_in  => LambdaIn(136));

  transition_508_preds(0) <= place_1202_token;
  LambdaOut(139) <= transition_508_symbol_out;
  transition_508 : transition
    port map(
      preds      => transition_508_preds,
      symbol_out => transition_508_symbol_out,
      symbol_in  => true);

  transition_509_preds(0) <= place_512_token;
  transition_509 : transition
    port map(
      preds      => transition_509_preds,
      symbol_out => transition_509_symbol_out,
      symbol_in  => LambdaIn(137));

  transition_510_preds(0) <= place_513_token;
  LambdaOut(140) <= transition_510_symbol_out;
  transition_510 : transition
    port map(
      preds      => transition_510_preds,
      symbol_out => transition_510_symbol_out,
      symbol_in  => true);

  transition_511_preds(0) <= place_514_token;
  transition_511 : transition
    port map(
      preds      => transition_511_preds,
      symbol_out => transition_511_symbol_out,
      symbol_in  => LambdaIn(138));

  transition_515_preds(0) <= place_1203_token;
  LambdaOut(141) <= transition_515_symbol_out;
  transition_515 : transition
    port map(
      preds      => transition_515_preds,
      symbol_out => transition_515_symbol_out,
      symbol_in  => true);

  transition_516_preds(0) <= place_519_token;
  transition_516 : transition
    port map(
      preds      => transition_516_preds,
      symbol_out => transition_516_symbol_out,
      symbol_in  => LambdaIn(139));

  transition_517_preds(0) <= place_520_token;
  LambdaOut(142) <= transition_517_symbol_out;
  transition_517 : transition
    port map(
      preds      => transition_517_preds,
      symbol_out => transition_517_symbol_out,
      symbol_in  => true);

  transition_518_preds(0) <= place_521_token;
  transition_518 : transition
    port map(
      preds      => transition_518_preds,
      symbol_out => transition_518_symbol_out,
      symbol_in  => LambdaIn(140));

  transition_522_preds(0) <= place_1198_token;
  transition_522_preds(1) <= place_1201_token;
  transition_522 : transition
    port map(
      preds      => transition_522_preds,
      symbol_out => transition_522_symbol_out,
      symbol_in  => true);

  transition_523_preds(0) <= place_1206_token;
  LambdaOut(143) <= transition_523_symbol_out;
  transition_523 : transition
    port map(
      preds      => transition_523_preds,
      symbol_out => transition_523_symbol_out,
      symbol_in  => true);

  transition_524_preds(0) <= place_527_token;
  transition_524 : transition
    port map(
      preds      => transition_524_preds,
      symbol_out => transition_524_symbol_out,
      symbol_in  => LambdaIn(141));

  transition_525_preds(0) <= place_528_token;
  LambdaOut(144) <= transition_525_symbol_out;
  transition_525 : transition
    port map(
      preds      => transition_525_preds,
      symbol_out => transition_525_symbol_out,
      symbol_in  => true);

  transition_526_preds(0) <= place_529_token;
  transition_526 : transition
    port map(
      preds      => transition_526_preds,
      symbol_out => transition_526_symbol_out,
      symbol_in  => LambdaIn(142));

  transition_530_preds(0) <= place_1207_token;
  LambdaOut(145) <= transition_530_symbol_out;
  transition_530 : transition
    port map(
      preds      => transition_530_preds,
      symbol_out => transition_530_symbol_out,
      symbol_in  => true);

  transition_531_preds(0) <= place_534_token;
  transition_531 : transition
    port map(
      preds      => transition_531_preds,
      symbol_out => transition_531_symbol_out,
      symbol_in  => LambdaIn(143));

  transition_532_preds(0) <= place_535_token;
  LambdaOut(146) <= transition_532_symbol_out;
  transition_532 : transition
    port map(
      preds      => transition_532_preds,
      symbol_out => transition_532_symbol_out,
      symbol_in  => true);

  transition_533_preds(0) <= place_536_token;
  transition_533 : transition
    port map(
      preds      => transition_533_preds,
      symbol_out => transition_533_symbol_out,
      symbol_in  => LambdaIn(144));

  transition_537_preds(0) <= place_1204_token;
  transition_537_preds(1) <= place_1205_token;
  transition_537 : transition
    port map(
      preds      => transition_537_preds,
      symbol_out => transition_537_symbol_out,
      symbol_in  => true);

  transition_538_preds(0) <= place_1208_token;
  LambdaOut(147) <= transition_538_symbol_out;
  transition_538 : transition
    port map(
      preds      => transition_538_preds,
      symbol_out => transition_538_symbol_out,
      symbol_in  => true);

  transition_539_preds(0) <= place_542_token;
  transition_539 : transition
    port map(
      preds      => transition_539_preds,
      symbol_out => transition_539_symbol_out,
      symbol_in  => LambdaIn(145));

  transition_540_preds(0) <= place_543_token;
  LambdaOut(148) <= transition_540_symbol_out;
  transition_540 : transition
    port map(
      preds      => transition_540_preds,
      symbol_out => transition_540_symbol_out,
      symbol_in  => true);

  transition_541_preds(0) <= place_544_token;
  transition_541 : transition
    port map(
      preds      => transition_541_preds,
      symbol_out => transition_541_symbol_out,
      symbol_in  => LambdaIn(146));

  transition_546_preds(0) <= place_545_token;
  transition_546 : transition
    port map(
      preds      => transition_546_preds,
      symbol_out => transition_546_symbol_out,
      symbol_in  => LambdaIn(147));

  transition_547_preds(0) <= place_1210_token;
  LambdaOut(149) <= transition_547_symbol_out;
  transition_547 : transition
    port map(
      preds      => transition_547_preds,
      symbol_out => transition_547_symbol_out,
      symbol_in  => true);

  transition_548_preds(0) <= place_1196_token;
  transition_548_preds(1) <= place_1209_token;
  transition_548 : transition
    port map(
      preds      => transition_548_preds,
      symbol_out => transition_548_symbol_out,
      symbol_in  => true);

  transition_549_preds(0) <= place_1213_token;
  LambdaOut(150) <= transition_549_symbol_out;
  transition_549 : transition
    port map(
      preds      => transition_549_preds,
      symbol_out => transition_549_symbol_out,
      symbol_in  => true);

  transition_550_preds(0) <= place_553_token;
  transition_550 : transition
    port map(
      preds      => transition_550_preds,
      symbol_out => transition_550_symbol_out,
      symbol_in  => LambdaIn(148));

  transition_551_preds(0) <= place_554_token;
  LambdaOut(151) <= transition_551_symbol_out;
  transition_551 : transition
    port map(
      preds      => transition_551_preds,
      symbol_out => transition_551_symbol_out,
      symbol_in  => true);

  transition_552_preds(0) <= place_555_token;
  transition_552 : transition
    port map(
      preds      => transition_552_preds,
      symbol_out => transition_552_symbol_out,
      symbol_in  => LambdaIn(149));

  transition_556_preds(0) <= place_1215_token;
  LambdaOut(152) <= transition_556_symbol_out;
  transition_556 : transition
    port map(
      preds      => transition_556_preds,
      symbol_out => transition_556_symbol_out,
      symbol_in  => true);

  transition_557_preds(0) <= place_560_token;
  transition_557 : transition
    port map(
      preds      => transition_557_preds,
      symbol_out => transition_557_symbol_out,
      symbol_in  => LambdaIn(150));

  transition_558_preds(0) <= place_561_token;
  LambdaOut(153) <= transition_558_symbol_out;
  transition_558 : transition
    port map(
      preds      => transition_558_preds,
      symbol_out => transition_558_symbol_out,
      symbol_in  => true);

  transition_559_preds(0) <= place_562_token;
  transition_559 : transition
    port map(
      preds      => transition_559_preds,
      symbol_out => transition_559_symbol_out,
      symbol_in  => LambdaIn(151));

  transition_563_preds(0) <= place_1216_token;
  LambdaOut(154) <= transition_563_symbol_out;
  transition_563 : transition
    port map(
      preds      => transition_563_preds,
      symbol_out => transition_563_symbol_out,
      symbol_in  => true);

  transition_564_preds(0) <= place_567_token;
  transition_564 : transition
    port map(
      preds      => transition_564_preds,
      symbol_out => transition_564_symbol_out,
      symbol_in  => LambdaIn(152));

  transition_565_preds(0) <= place_568_token;
  LambdaOut(155) <= transition_565_symbol_out;
  transition_565 : transition
    port map(
      preds      => transition_565_preds,
      symbol_out => transition_565_symbol_out,
      symbol_in  => true);

  transition_566_preds(0) <= place_569_token;
  transition_566 : transition
    port map(
      preds      => transition_566_preds,
      symbol_out => transition_566_symbol_out,
      symbol_in  => LambdaIn(153));

  transition_570_preds(0) <= place_1214_token;
  transition_570_preds(1) <= place_1212_token;
  transition_570 : transition
    port map(
      preds      => transition_570_preds,
      symbol_out => transition_570_symbol_out,
      symbol_in  => true);

  transition_571_preds(0) <= place_1219_token;
  LambdaOut(156) <= transition_571_symbol_out;
  transition_571 : transition
    port map(
      preds      => transition_571_preds,
      symbol_out => transition_571_symbol_out,
      symbol_in  => true);

  transition_572_preds(0) <= place_575_token;
  transition_572 : transition
    port map(
      preds      => transition_572_preds,
      symbol_out => transition_572_symbol_out,
      symbol_in  => LambdaIn(154));

  transition_573_preds(0) <= place_576_token;
  LambdaOut(157) <= transition_573_symbol_out;
  transition_573 : transition
    port map(
      preds      => transition_573_preds,
      symbol_out => transition_573_symbol_out,
      symbol_in  => true);

  transition_574_preds(0) <= place_577_token;
  transition_574 : transition
    port map(
      preds      => transition_574_preds,
      symbol_out => transition_574_symbol_out,
      symbol_in  => LambdaIn(155));

  transition_578_preds(0) <= place_1220_token;
  LambdaOut(158) <= transition_578_symbol_out;
  transition_578 : transition
    port map(
      preds      => transition_578_preds,
      symbol_out => transition_578_symbol_out,
      symbol_in  => true);

  transition_579_preds(0) <= place_582_token;
  transition_579 : transition
    port map(
      preds      => transition_579_preds,
      symbol_out => transition_579_symbol_out,
      symbol_in  => LambdaIn(156));

  transition_580_preds(0) <= place_583_token;
  LambdaOut(159) <= transition_580_symbol_out;
  transition_580 : transition
    port map(
      preds      => transition_580_preds,
      symbol_out => transition_580_symbol_out,
      symbol_in  => true);

  transition_581_preds(0) <= place_584_token;
  transition_581 : transition
    port map(
      preds      => transition_581_preds,
      symbol_out => transition_581_symbol_out,
      symbol_in  => LambdaIn(157));

  transition_585_preds(0) <= place_1217_token;
  transition_585_preds(1) <= place_1218_token;
  transition_585 : transition
    port map(
      preds      => transition_585_preds,
      symbol_out => transition_585_symbol_out,
      symbol_in  => true);

  transition_586_preds(0) <= place_1221_token;
  LambdaOut(160) <= transition_586_symbol_out;
  transition_586 : transition
    port map(
      preds      => transition_586_preds,
      symbol_out => transition_586_symbol_out,
      symbol_in  => true);

  transition_587_preds(0) <= place_590_token;
  transition_587 : transition
    port map(
      preds      => transition_587_preds,
      symbol_out => transition_587_symbol_out,
      symbol_in  => LambdaIn(158));

  transition_588_preds(0) <= place_591_token;
  LambdaOut(161) <= transition_588_symbol_out;
  transition_588 : transition
    port map(
      preds      => transition_588_preds,
      symbol_out => transition_588_symbol_out,
      symbol_in  => true);

  transition_589_preds(0) <= place_592_token;
  transition_589 : transition
    port map(
      preds      => transition_589_preds,
      symbol_out => transition_589_symbol_out,
      symbol_in  => LambdaIn(159));

  transition_594_preds(0) <= place_593_token;
  transition_594 : transition
    port map(
      preds      => transition_594_preds,
      symbol_out => transition_594_symbol_out,
      symbol_in  => LambdaIn(160));

  transition_595_preds(0) <= place_1224_token;
  LambdaOut(162) <= transition_595_symbol_out;
  transition_595 : transition
    port map(
      preds      => transition_595_preds,
      symbol_out => transition_595_symbol_out,
      symbol_in  => true);

  transition_596_preds(0) <= place_1211_token;
  transition_596_preds(1) <= place_1223_token;
  transition_596 : transition
    port map(
      preds      => transition_596_preds,
      symbol_out => transition_596_symbol_out,
      symbol_in  => true);

  transition_597_preds(0) <= place_1228_token;
  LambdaOut(163) <= transition_597_symbol_out;
  transition_597 : transition
    port map(
      preds      => transition_597_preds,
      symbol_out => transition_597_symbol_out,
      symbol_in  => true);

  transition_598_preds(0) <= place_601_token;
  transition_598 : transition
    port map(
      preds      => transition_598_preds,
      symbol_out => transition_598_symbol_out,
      symbol_in  => LambdaIn(161));

  transition_599_preds(0) <= place_602_token;
  LambdaOut(164) <= transition_599_symbol_out;
  transition_599 : transition
    port map(
      preds      => transition_599_preds,
      symbol_out => transition_599_symbol_out,
      symbol_in  => true);

  transition_600_preds(0) <= place_603_token;
  transition_600 : transition
    port map(
      preds      => transition_600_preds,
      symbol_out => transition_600_symbol_out,
      symbol_in  => LambdaIn(162));

  transition_604_preds(0) <= place_1230_token;
  LambdaOut(165) <= transition_604_symbol_out;
  transition_604 : transition
    port map(
      preds      => transition_604_preds,
      symbol_out => transition_604_symbol_out,
      symbol_in  => true);

  transition_605_preds(0) <= place_608_token;
  transition_605 : transition
    port map(
      preds      => transition_605_preds,
      symbol_out => transition_605_symbol_out,
      symbol_in  => LambdaIn(163));

  transition_606_preds(0) <= place_609_token;
  LambdaOut(166) <= transition_606_symbol_out;
  transition_606 : transition
    port map(
      preds      => transition_606_preds,
      symbol_out => transition_606_symbol_out,
      symbol_in  => true);

  transition_607_preds(0) <= place_610_token;
  transition_607 : transition
    port map(
      preds      => transition_607_preds,
      symbol_out => transition_607_symbol_out,
      symbol_in  => LambdaIn(164));

  transition_611_preds(0) <= place_1231_token;
  LambdaOut(167) <= transition_611_symbol_out;
  transition_611 : transition
    port map(
      preds      => transition_611_preds,
      symbol_out => transition_611_symbol_out,
      symbol_in  => true);

  transition_612_preds(0) <= place_615_token;
  transition_612 : transition
    port map(
      preds      => transition_612_preds,
      symbol_out => transition_612_symbol_out,
      symbol_in  => LambdaIn(165));

  transition_613_preds(0) <= place_616_token;
  LambdaOut(168) <= transition_613_symbol_out;
  transition_613 : transition
    port map(
      preds      => transition_613_preds,
      symbol_out => transition_613_symbol_out,
      symbol_in  => true);

  transition_614_preds(0) <= place_617_token;
  transition_614 : transition
    port map(
      preds      => transition_614_preds,
      symbol_out => transition_614_symbol_out,
      symbol_in  => LambdaIn(166));

  transition_618_preds(0) <= place_1226_token;
  transition_618_preds(1) <= place_1229_token;
  transition_618 : transition
    port map(
      preds      => transition_618_preds,
      symbol_out => transition_618_symbol_out,
      symbol_in  => true);

  transition_619_preds(0) <= place_1234_token;
  LambdaOut(169) <= transition_619_symbol_out;
  transition_619 : transition
    port map(
      preds      => transition_619_preds,
      symbol_out => transition_619_symbol_out,
      symbol_in  => true);

  transition_620_preds(0) <= place_623_token;
  transition_620 : transition
    port map(
      preds      => transition_620_preds,
      symbol_out => transition_620_symbol_out,
      symbol_in  => LambdaIn(167));

  transition_621_preds(0) <= place_624_token;
  LambdaOut(170) <= transition_621_symbol_out;
  transition_621 : transition
    port map(
      preds      => transition_621_preds,
      symbol_out => transition_621_symbol_out,
      symbol_in  => true);

  transition_622_preds(0) <= place_625_token;
  transition_622 : transition
    port map(
      preds      => transition_622_preds,
      symbol_out => transition_622_symbol_out,
      symbol_in  => LambdaIn(168));

  transition_626_preds(0) <= place_1235_token;
  LambdaOut(171) <= transition_626_symbol_out;
  transition_626 : transition
    port map(
      preds      => transition_626_preds,
      symbol_out => transition_626_symbol_out,
      symbol_in  => true);

  transition_627_preds(0) <= place_630_token;
  transition_627 : transition
    port map(
      preds      => transition_627_preds,
      symbol_out => transition_627_symbol_out,
      symbol_in  => LambdaIn(169));

  transition_628_preds(0) <= place_631_token;
  LambdaOut(172) <= transition_628_symbol_out;
  transition_628 : transition
    port map(
      preds      => transition_628_preds,
      symbol_out => transition_628_symbol_out,
      symbol_in  => true);

  transition_629_preds(0) <= place_632_token;
  transition_629 : transition
    port map(
      preds      => transition_629_preds,
      symbol_out => transition_629_symbol_out,
      symbol_in  => LambdaIn(170));

  transition_633_preds(0) <= place_1232_token;
  transition_633_preds(1) <= place_1233_token;
  transition_633 : transition
    port map(
      preds      => transition_633_preds,
      symbol_out => transition_633_symbol_out,
      symbol_in  => true);

  transition_634_preds(0) <= place_1236_token;
  LambdaOut(173) <= transition_634_symbol_out;
  transition_634 : transition
    port map(
      preds      => transition_634_preds,
      symbol_out => transition_634_symbol_out,
      symbol_in  => true);

  transition_635_preds(0) <= place_638_token;
  transition_635 : transition
    port map(
      preds      => transition_635_preds,
      symbol_out => transition_635_symbol_out,
      symbol_in  => LambdaIn(171));

  transition_636_preds(0) <= place_639_token;
  LambdaOut(174) <= transition_636_symbol_out;
  transition_636 : transition
    port map(
      preds      => transition_636_preds,
      symbol_out => transition_636_symbol_out,
      symbol_in  => true);

  transition_637_preds(0) <= place_640_token;
  transition_637 : transition
    port map(
      preds      => transition_637_preds,
      symbol_out => transition_637_symbol_out,
      symbol_in  => LambdaIn(172));

  transition_642_preds(0) <= place_641_token;
  transition_642 : transition
    port map(
      preds      => transition_642_preds,
      symbol_out => transition_642_symbol_out,
      symbol_in  => LambdaIn(173));

  transition_643_preds(0) <= place_1239_token;
  LambdaOut(175) <= transition_643_symbol_out;
  transition_643 : transition
    port map(
      preds      => transition_643_preds,
      symbol_out => transition_643_symbol_out,
      symbol_in  => true);

  transition_644_preds(0) <= place_1225_token;
  transition_644_preds(1) <= place_1238_token;
  transition_644 : transition
    port map(
      preds      => transition_644_preds,
      symbol_out => transition_644_symbol_out,
      symbol_in  => true);

  transition_645_preds(0) <= place_1243_token;
  LambdaOut(176) <= transition_645_symbol_out;
  transition_645 : transition
    port map(
      preds      => transition_645_preds,
      symbol_out => transition_645_symbol_out,
      symbol_in  => true);

  transition_646_preds(0) <= place_649_token;
  transition_646 : transition
    port map(
      preds      => transition_646_preds,
      symbol_out => transition_646_symbol_out,
      symbol_in  => LambdaIn(174));

  transition_647_preds(0) <= place_650_token;
  LambdaOut(177) <= transition_647_symbol_out;
  transition_647 : transition
    port map(
      preds      => transition_647_preds,
      symbol_out => transition_647_symbol_out,
      symbol_in  => true);

  transition_648_preds(0) <= place_651_token;
  transition_648 : transition
    port map(
      preds      => transition_648_preds,
      symbol_out => transition_648_symbol_out,
      symbol_in  => LambdaIn(175));

  transition_652_preds(0) <= place_1245_token;
  LambdaOut(178) <= transition_652_symbol_out;
  transition_652 : transition
    port map(
      preds      => transition_652_preds,
      symbol_out => transition_652_symbol_out,
      symbol_in  => true);

  transition_653_preds(0) <= place_656_token;
  transition_653 : transition
    port map(
      preds      => transition_653_preds,
      symbol_out => transition_653_symbol_out,
      symbol_in  => LambdaIn(176));

  transition_654_preds(0) <= place_657_token;
  LambdaOut(179) <= transition_654_symbol_out;
  transition_654 : transition
    port map(
      preds      => transition_654_preds,
      symbol_out => transition_654_symbol_out,
      symbol_in  => true);

  transition_655_preds(0) <= place_658_token;
  transition_655 : transition
    port map(
      preds      => transition_655_preds,
      symbol_out => transition_655_symbol_out,
      symbol_in  => LambdaIn(177));

  transition_659_preds(0) <= place_1246_token;
  LambdaOut(180) <= transition_659_symbol_out;
  transition_659 : transition
    port map(
      preds      => transition_659_preds,
      symbol_out => transition_659_symbol_out,
      symbol_in  => true);

  transition_660_preds(0) <= place_663_token;
  transition_660 : transition
    port map(
      preds      => transition_660_preds,
      symbol_out => transition_660_symbol_out,
      symbol_in  => LambdaIn(178));

  transition_661_preds(0) <= place_664_token;
  LambdaOut(181) <= transition_661_symbol_out;
  transition_661 : transition
    port map(
      preds      => transition_661_preds,
      symbol_out => transition_661_symbol_out,
      symbol_in  => true);

  transition_662_preds(0) <= place_665_token;
  transition_662 : transition
    port map(
      preds      => transition_662_preds,
      symbol_out => transition_662_symbol_out,
      symbol_in  => LambdaIn(179));

  transition_666_preds(0) <= place_1242_token;
  transition_666_preds(1) <= place_1244_token;
  transition_666 : transition
    port map(
      preds      => transition_666_preds,
      symbol_out => transition_666_symbol_out,
      symbol_in  => true);

  transition_667_preds(0) <= place_1250_token;
  LambdaOut(182) <= transition_667_symbol_out;
  transition_667 : transition
    port map(
      preds      => transition_667_preds,
      symbol_out => transition_667_symbol_out,
      symbol_in  => true);

  transition_668_preds(0) <= place_671_token;
  transition_668 : transition
    port map(
      preds      => transition_668_preds,
      symbol_out => transition_668_symbol_out,
      symbol_in  => LambdaIn(180));

  transition_669_preds(0) <= place_672_token;
  LambdaOut(183) <= transition_669_symbol_out;
  transition_669 : transition
    port map(
      preds      => transition_669_preds,
      symbol_out => transition_669_symbol_out,
      symbol_in  => true);

  transition_670_preds(0) <= place_673_token;
  transition_670 : transition
    port map(
      preds      => transition_670_preds,
      symbol_out => transition_670_symbol_out,
      symbol_in  => LambdaIn(181));

  transition_674_preds(0) <= place_1251_token;
  LambdaOut(184) <= transition_674_symbol_out;
  transition_674 : transition
    port map(
      preds      => transition_674_preds,
      symbol_out => transition_674_symbol_out,
      symbol_in  => true);

  transition_675_preds(0) <= place_678_token;
  transition_675 : transition
    port map(
      preds      => transition_675_preds,
      symbol_out => transition_675_symbol_out,
      symbol_in  => LambdaIn(182));

  transition_676_preds(0) <= place_679_token;
  LambdaOut(185) <= transition_676_symbol_out;
  transition_676 : transition
    port map(
      preds      => transition_676_preds,
      symbol_out => transition_676_symbol_out,
      symbol_in  => true);

  transition_677_preds(0) <= place_680_token;
  transition_677 : transition
    port map(
      preds      => transition_677_preds,
      symbol_out => transition_677_symbol_out,
      symbol_in  => LambdaIn(183));

  transition_681_preds(0) <= place_1247_token;
  transition_681_preds(1) <= place_1249_token;
  transition_681 : transition
    port map(
      preds      => transition_681_preds,
      symbol_out => transition_681_symbol_out,
      symbol_in  => true);

  transition_682_preds(0) <= place_1252_token;
  LambdaOut(186) <= transition_682_symbol_out;
  transition_682 : transition
    port map(
      preds      => transition_682_preds,
      symbol_out => transition_682_symbol_out,
      symbol_in  => true);

  transition_683_preds(0) <= place_686_token;
  transition_683 : transition
    port map(
      preds      => transition_683_preds,
      symbol_out => transition_683_symbol_out,
      symbol_in  => LambdaIn(184));

  transition_684_preds(0) <= place_687_token;
  LambdaOut(187) <= transition_684_symbol_out;
  transition_684 : transition
    port map(
      preds      => transition_684_preds,
      symbol_out => transition_684_symbol_out,
      symbol_in  => true);

  transition_685_preds(0) <= place_688_token;
  transition_685 : transition
    port map(
      preds      => transition_685_preds,
      symbol_out => transition_685_symbol_out,
      symbol_in  => LambdaIn(185));

  transition_690_preds(0) <= place_689_token;
  transition_690 : transition
    port map(
      preds      => transition_690_preds,
      symbol_out => transition_690_symbol_out,
      symbol_in  => LambdaIn(186));

  transition_691_preds(0) <= place_1254_token;
  LambdaOut(188) <= transition_691_symbol_out;
  transition_691 : transition
    port map(
      preds      => transition_691_preds,
      symbol_out => transition_691_symbol_out,
      symbol_in  => true);

  transition_692_preds(0) <= place_1240_token;
  transition_692_preds(1) <= place_1253_token;
  transition_692 : transition
    port map(
      preds      => transition_692_preds,
      symbol_out => transition_692_symbol_out,
      symbol_in  => true);

  transition_693_preds(0) <= place_1257_token;
  LambdaOut(189) <= transition_693_symbol_out;
  transition_693 : transition
    port map(
      preds      => transition_693_preds,
      symbol_out => transition_693_symbol_out,
      symbol_in  => true);

  transition_694_preds(0) <= place_697_token;
  transition_694 : transition
    port map(
      preds      => transition_694_preds,
      symbol_out => transition_694_symbol_out,
      symbol_in  => LambdaIn(187));

  transition_695_preds(0) <= place_698_token;
  LambdaOut(190) <= transition_695_symbol_out;
  transition_695 : transition
    port map(
      preds      => transition_695_preds,
      symbol_out => transition_695_symbol_out,
      symbol_in  => true);

  transition_696_preds(0) <= place_699_token;
  transition_696 : transition
    port map(
      preds      => transition_696_preds,
      symbol_out => transition_696_symbol_out,
      symbol_in  => LambdaIn(188));

  transition_700_preds(0) <= place_1259_token;
  LambdaOut(191) <= transition_700_symbol_out;
  transition_700 : transition
    port map(
      preds      => transition_700_preds,
      symbol_out => transition_700_symbol_out,
      symbol_in  => true);

  transition_701_preds(0) <= place_704_token;
  transition_701 : transition
    port map(
      preds      => transition_701_preds,
      symbol_out => transition_701_symbol_out,
      symbol_in  => LambdaIn(189));

  transition_702_preds(0) <= place_705_token;
  LambdaOut(192) <= transition_702_symbol_out;
  transition_702 : transition
    port map(
      preds      => transition_702_preds,
      symbol_out => transition_702_symbol_out,
      symbol_in  => true);

  transition_703_preds(0) <= place_706_token;
  transition_703 : transition
    port map(
      preds      => transition_703_preds,
      symbol_out => transition_703_symbol_out,
      symbol_in  => LambdaIn(190));

  transition_707_preds(0) <= place_1260_token;
  LambdaOut(193) <= transition_707_symbol_out;
  transition_707 : transition
    port map(
      preds      => transition_707_preds,
      symbol_out => transition_707_symbol_out,
      symbol_in  => true);

  transition_708_preds(0) <= place_711_token;
  transition_708 : transition
    port map(
      preds      => transition_708_preds,
      symbol_out => transition_708_symbol_out,
      symbol_in  => LambdaIn(191));

  transition_709_preds(0) <= place_712_token;
  LambdaOut(194) <= transition_709_symbol_out;
  transition_709 : transition
    port map(
      preds      => transition_709_preds,
      symbol_out => transition_709_symbol_out,
      symbol_in  => true);

  transition_710_preds(0) <= place_713_token;
  transition_710 : transition
    port map(
      preds      => transition_710_preds,
      symbol_out => transition_710_symbol_out,
      symbol_in  => LambdaIn(192));

  transition_714_preds(0) <= place_1258_token;
  transition_714_preds(1) <= place_1256_token;
  transition_714 : transition
    port map(
      preds      => transition_714_preds,
      symbol_out => transition_714_symbol_out,
      symbol_in  => true);

  transition_715_preds(0) <= place_1263_token;
  LambdaOut(195) <= transition_715_symbol_out;
  transition_715 : transition
    port map(
      preds      => transition_715_preds,
      symbol_out => transition_715_symbol_out,
      symbol_in  => true);

  transition_716_preds(0) <= place_719_token;
  transition_716 : transition
    port map(
      preds      => transition_716_preds,
      symbol_out => transition_716_symbol_out,
      symbol_in  => LambdaIn(193));

  transition_717_preds(0) <= place_720_token;
  LambdaOut(196) <= transition_717_symbol_out;
  transition_717 : transition
    port map(
      preds      => transition_717_preds,
      symbol_out => transition_717_symbol_out,
      symbol_in  => true);

  transition_718_preds(0) <= place_721_token;
  transition_718 : transition
    port map(
      preds      => transition_718_preds,
      symbol_out => transition_718_symbol_out,
      symbol_in  => LambdaIn(194));

  transition_722_preds(0) <= place_1264_token;
  LambdaOut(197) <= transition_722_symbol_out;
  transition_722 : transition
    port map(
      preds      => transition_722_preds,
      symbol_out => transition_722_symbol_out,
      symbol_in  => true);

  transition_723_preds(0) <= place_726_token;
  transition_723 : transition
    port map(
      preds      => transition_723_preds,
      symbol_out => transition_723_symbol_out,
      symbol_in  => LambdaIn(195));

  transition_724_preds(0) <= place_727_token;
  LambdaOut(198) <= transition_724_symbol_out;
  transition_724 : transition
    port map(
      preds      => transition_724_preds,
      symbol_out => transition_724_symbol_out,
      symbol_in  => true);

  transition_725_preds(0) <= place_728_token;
  transition_725 : transition
    port map(
      preds      => transition_725_preds,
      symbol_out => transition_725_symbol_out,
      symbol_in  => LambdaIn(196));

  transition_729_preds(0) <= place_1261_token;
  transition_729_preds(1) <= place_1262_token;
  transition_729 : transition
    port map(
      preds      => transition_729_preds,
      symbol_out => transition_729_symbol_out,
      symbol_in  => true);

  transition_730_preds(0) <= place_1265_token;
  LambdaOut(199) <= transition_730_symbol_out;
  transition_730 : transition
    port map(
      preds      => transition_730_preds,
      symbol_out => transition_730_symbol_out,
      symbol_in  => true);

  transition_731_preds(0) <= place_734_token;
  transition_731 : transition
    port map(
      preds      => transition_731_preds,
      symbol_out => transition_731_symbol_out,
      symbol_in  => LambdaIn(197));

  transition_732_preds(0) <= place_735_token;
  LambdaOut(200) <= transition_732_symbol_out;
  transition_732 : transition
    port map(
      preds      => transition_732_preds,
      symbol_out => transition_732_symbol_out,
      symbol_in  => true);

  transition_733_preds(0) <= place_736_token;
  transition_733 : transition
    port map(
      preds      => transition_733_preds,
      symbol_out => transition_733_symbol_out,
      symbol_in  => LambdaIn(198));

  transition_738_preds(0) <= place_737_token;
  transition_738 : transition
    port map(
      preds      => transition_738_preds,
      symbol_out => transition_738_symbol_out,
      symbol_in  => LambdaIn(199));

  transition_739_preds(0) <= place_1267_token;
  LambdaOut(201) <= transition_739_symbol_out;
  transition_739 : transition
    port map(
      preds      => transition_739_preds,
      symbol_out => transition_739_symbol_out,
      symbol_in  => true);

  transition_740_preds(0) <= place_1255_token;
  transition_740_preds(1) <= place_1266_token;
  transition_740 : transition
    port map(
      preds      => transition_740_preds,
      symbol_out => transition_740_symbol_out,
      symbol_in  => true);

  transition_741_preds(0) <= place_1271_token;
  LambdaOut(202) <= transition_741_symbol_out;
  transition_741 : transition
    port map(
      preds      => transition_741_preds,
      symbol_out => transition_741_symbol_out,
      symbol_in  => true);

  transition_742_preds(0) <= place_745_token;
  transition_742 : transition
    port map(
      preds      => transition_742_preds,
      symbol_out => transition_742_symbol_out,
      symbol_in  => LambdaIn(200));

  transition_743_preds(0) <= place_746_token;
  LambdaOut(203) <= transition_743_symbol_out;
  transition_743 : transition
    port map(
      preds      => transition_743_preds,
      symbol_out => transition_743_symbol_out,
      symbol_in  => true);

  transition_744_preds(0) <= place_747_token;
  transition_744 : transition
    port map(
      preds      => transition_744_preds,
      symbol_out => transition_744_symbol_out,
      symbol_in  => LambdaIn(201));

  transition_748_preds(0) <= place_1274_token;
  LambdaOut(204) <= transition_748_symbol_out;
  transition_748 : transition
    port map(
      preds      => transition_748_preds,
      symbol_out => transition_748_symbol_out,
      symbol_in  => true);

  transition_749_preds(0) <= place_752_token;
  transition_749 : transition
    port map(
      preds      => transition_749_preds,
      symbol_out => transition_749_symbol_out,
      symbol_in  => LambdaIn(202));

  transition_750_preds(0) <= place_753_token;
  LambdaOut(205) <= transition_750_symbol_out;
  transition_750 : transition
    port map(
      preds      => transition_750_preds,
      symbol_out => transition_750_symbol_out,
      symbol_in  => true);

  transition_751_preds(0) <= place_754_token;
  transition_751 : transition
    port map(
      preds      => transition_751_preds,
      symbol_out => transition_751_symbol_out,
      symbol_in  => LambdaIn(203));

  transition_755_preds(0) <= place_1275_token;
  LambdaOut(206) <= transition_755_symbol_out;
  transition_755 : transition
    port map(
      preds      => transition_755_preds,
      symbol_out => transition_755_symbol_out,
      symbol_in  => true);

  transition_756_preds(0) <= place_759_token;
  transition_756 : transition
    port map(
      preds      => transition_756_preds,
      symbol_out => transition_756_symbol_out,
      symbol_in  => LambdaIn(204));

  transition_757_preds(0) <= place_760_token;
  LambdaOut(207) <= transition_757_symbol_out;
  transition_757 : transition
    port map(
      preds      => transition_757_preds,
      symbol_out => transition_757_symbol_out,
      symbol_in  => true);

  transition_758_preds(0) <= place_761_token;
  transition_758 : transition
    port map(
      preds      => transition_758_preds,
      symbol_out => transition_758_symbol_out,
      symbol_in  => LambdaIn(205));

  transition_762_preds(0) <= place_1272_token;
  transition_762_preds(1) <= place_1270_token;
  transition_762 : transition
    port map(
      preds      => transition_762_preds,
      symbol_out => transition_762_symbol_out,
      symbol_in  => true);

  transition_763_preds(0) <= place_1278_token;
  LambdaOut(208) <= transition_763_symbol_out;
  transition_763 : transition
    port map(
      preds      => transition_763_preds,
      symbol_out => transition_763_symbol_out,
      symbol_in  => true);

  transition_764_preds(0) <= place_767_token;
  transition_764 : transition
    port map(
      preds      => transition_764_preds,
      symbol_out => transition_764_symbol_out,
      symbol_in  => LambdaIn(206));

  transition_765_preds(0) <= place_768_token;
  LambdaOut(209) <= transition_765_symbol_out;
  transition_765 : transition
    port map(
      preds      => transition_765_preds,
      symbol_out => transition_765_symbol_out,
      symbol_in  => true);

  transition_766_preds(0) <= place_769_token;
  transition_766 : transition
    port map(
      preds      => transition_766_preds,
      symbol_out => transition_766_symbol_out,
      symbol_in  => LambdaIn(207));

  transition_770_preds(0) <= place_1279_token;
  LambdaOut(210) <= transition_770_symbol_out;
  transition_770 : transition
    port map(
      preds      => transition_770_preds,
      symbol_out => transition_770_symbol_out,
      symbol_in  => true);

  transition_771_preds(0) <= place_774_token;
  transition_771 : transition
    port map(
      preds      => transition_771_preds,
      symbol_out => transition_771_symbol_out,
      symbol_in  => LambdaIn(208));

  transition_772_preds(0) <= place_775_token;
  LambdaOut(211) <= transition_772_symbol_out;
  transition_772 : transition
    port map(
      preds      => transition_772_preds,
      symbol_out => transition_772_symbol_out,
      symbol_in  => true);

  transition_773_preds(0) <= place_776_token;
  transition_773 : transition
    port map(
      preds      => transition_773_preds,
      symbol_out => transition_773_symbol_out,
      symbol_in  => LambdaIn(209));

  transition_777_preds(0) <= place_1276_token;
  transition_777_preds(1) <= place_1277_token;
  transition_777 : transition
    port map(
      preds      => transition_777_preds,
      symbol_out => transition_777_symbol_out,
      symbol_in  => true);

  transition_778_preds(0) <= place_1280_token;
  LambdaOut(212) <= transition_778_symbol_out;
  transition_778 : transition
    port map(
      preds      => transition_778_preds,
      symbol_out => transition_778_symbol_out,
      symbol_in  => true);

  transition_779_preds(0) <= place_782_token;
  transition_779 : transition
    port map(
      preds      => transition_779_preds,
      symbol_out => transition_779_symbol_out,
      symbol_in  => LambdaIn(210));

  transition_780_preds(0) <= place_783_token;
  LambdaOut(213) <= transition_780_symbol_out;
  transition_780 : transition
    port map(
      preds      => transition_780_preds,
      symbol_out => transition_780_symbol_out,
      symbol_in  => true);

  transition_781_preds(0) <= place_784_token;
  transition_781 : transition
    port map(
      preds      => transition_781_preds,
      symbol_out => transition_781_symbol_out,
      symbol_in  => LambdaIn(211));

  transition_786_preds(0) <= place_785_token;
  transition_786 : transition
    port map(
      preds      => transition_786_preds,
      symbol_out => transition_786_symbol_out,
      symbol_in  => LambdaIn(212));

  transition_787_preds(0) <= place_1282_token;
  LambdaOut(214) <= transition_787_symbol_out;
  transition_787 : transition
    port map(
      preds      => transition_787_preds,
      symbol_out => transition_787_symbol_out,
      symbol_in  => true);

  transition_788_preds(0) <= place_1268_token;
  transition_788_preds(1) <= place_1281_token;
  transition_788 : transition
    port map(
      preds      => transition_788_preds,
      symbol_out => transition_788_symbol_out,
      symbol_in  => true);

  transition_789_preds(0) <= place_1285_token;
  LambdaOut(215) <= transition_789_symbol_out;
  transition_789 : transition
    port map(
      preds      => transition_789_preds,
      symbol_out => transition_789_symbol_out,
      symbol_in  => true);

  transition_790_preds(0) <= place_793_token;
  transition_790 : transition
    port map(
      preds      => transition_790_preds,
      symbol_out => transition_790_symbol_out,
      symbol_in  => LambdaIn(213));

  transition_791_preds(0) <= place_794_token;
  LambdaOut(216) <= transition_791_symbol_out;
  transition_791 : transition
    port map(
      preds      => transition_791_preds,
      symbol_out => transition_791_symbol_out,
      symbol_in  => true);

  transition_792_preds(0) <= place_795_token;
  transition_792 : transition
    port map(
      preds      => transition_792_preds,
      symbol_out => transition_792_symbol_out,
      symbol_in  => LambdaIn(214));

  transition_796_preds(0) <= place_1288_token;
  LambdaOut(217) <= transition_796_symbol_out;
  transition_796 : transition
    port map(
      preds      => transition_796_preds,
      symbol_out => transition_796_symbol_out,
      symbol_in  => true);

  transition_797_preds(0) <= place_800_token;
  transition_797 : transition
    port map(
      preds      => transition_797_preds,
      symbol_out => transition_797_symbol_out,
      symbol_in  => LambdaIn(215));

  transition_798_preds(0) <= place_801_token;
  LambdaOut(218) <= transition_798_symbol_out;
  transition_798 : transition
    port map(
      preds      => transition_798_preds,
      symbol_out => transition_798_symbol_out,
      symbol_in  => true);

  transition_799_preds(0) <= place_802_token;
  transition_799 : transition
    port map(
      preds      => transition_799_preds,
      symbol_out => transition_799_symbol_out,
      symbol_in  => LambdaIn(216));

  transition_803_preds(0) <= place_1289_token;
  LambdaOut(219) <= transition_803_symbol_out;
  transition_803 : transition
    port map(
      preds      => transition_803_preds,
      symbol_out => transition_803_symbol_out,
      symbol_in  => true);

  transition_804_preds(0) <= place_807_token;
  transition_804 : transition
    port map(
      preds      => transition_804_preds,
      symbol_out => transition_804_symbol_out,
      symbol_in  => LambdaIn(217));

  transition_805_preds(0) <= place_808_token;
  LambdaOut(220) <= transition_805_symbol_out;
  transition_805 : transition
    port map(
      preds      => transition_805_preds,
      symbol_out => transition_805_symbol_out,
      symbol_in  => true);

  transition_806_preds(0) <= place_809_token;
  transition_806 : transition
    port map(
      preds      => transition_806_preds,
      symbol_out => transition_806_symbol_out,
      symbol_in  => LambdaIn(218));

  transition_810_preds(0) <= place_1284_token;
  transition_810_preds(1) <= place_1287_token;
  transition_810 : transition
    port map(
      preds      => transition_810_preds,
      symbol_out => transition_810_symbol_out,
      symbol_in  => true);

  transition_811_preds(0) <= place_1292_token;
  LambdaOut(221) <= transition_811_symbol_out;
  transition_811 : transition
    port map(
      preds      => transition_811_preds,
      symbol_out => transition_811_symbol_out,
      symbol_in  => true);

  transition_812_preds(0) <= place_815_token;
  transition_812 : transition
    port map(
      preds      => transition_812_preds,
      symbol_out => transition_812_symbol_out,
      symbol_in  => LambdaIn(219));

  transition_813_preds(0) <= place_816_token;
  LambdaOut(222) <= transition_813_symbol_out;
  transition_813 : transition
    port map(
      preds      => transition_813_preds,
      symbol_out => transition_813_symbol_out,
      symbol_in  => true);

  transition_814_preds(0) <= place_817_token;
  transition_814 : transition
    port map(
      preds      => transition_814_preds,
      symbol_out => transition_814_symbol_out,
      symbol_in  => LambdaIn(220));

  transition_818_preds(0) <= place_1293_token;
  LambdaOut(223) <= transition_818_symbol_out;
  transition_818 : transition
    port map(
      preds      => transition_818_preds,
      symbol_out => transition_818_symbol_out,
      symbol_in  => true);

  transition_819_preds(0) <= place_822_token;
  transition_819 : transition
    port map(
      preds      => transition_819_preds,
      symbol_out => transition_819_symbol_out,
      symbol_in  => LambdaIn(221));

  transition_820_preds(0) <= place_823_token;
  LambdaOut(224) <= transition_820_symbol_out;
  transition_820 : transition
    port map(
      preds      => transition_820_preds,
      symbol_out => transition_820_symbol_out,
      symbol_in  => true);

  transition_821_preds(0) <= place_824_token;
  transition_821 : transition
    port map(
      preds      => transition_821_preds,
      symbol_out => transition_821_symbol_out,
      symbol_in  => LambdaIn(222));

  transition_825_preds(0) <= place_1290_token;
  transition_825_preds(1) <= place_1291_token;
  transition_825 : transition
    port map(
      preds      => transition_825_preds,
      symbol_out => transition_825_symbol_out,
      symbol_in  => true);

  transition_826_preds(0) <= place_1294_token;
  LambdaOut(225) <= transition_826_symbol_out;
  transition_826 : transition
    port map(
      preds      => transition_826_preds,
      symbol_out => transition_826_symbol_out,
      symbol_in  => true);

  transition_827_preds(0) <= place_830_token;
  transition_827 : transition
    port map(
      preds      => transition_827_preds,
      symbol_out => transition_827_symbol_out,
      symbol_in  => LambdaIn(223));

  transition_828_preds(0) <= place_831_token;
  LambdaOut(226) <= transition_828_symbol_out;
  transition_828 : transition
    port map(
      preds      => transition_828_preds,
      symbol_out => transition_828_symbol_out,
      symbol_in  => true);

  transition_829_preds(0) <= place_832_token;
  transition_829 : transition
    port map(
      preds      => transition_829_preds,
      symbol_out => transition_829_symbol_out,
      symbol_in  => LambdaIn(224));

  transition_834_preds(0) <= place_833_token;
  transition_834 : transition
    port map(
      preds      => transition_834_preds,
      symbol_out => transition_834_symbol_out,
      symbol_in  => LambdaIn(225));

  transition_835_preds(0) <= place_1296_token;
  LambdaOut(227) <= transition_835_symbol_out;
  transition_835 : transition
    port map(
      preds      => transition_835_preds,
      symbol_out => transition_835_symbol_out,
      symbol_in  => true);

  transition_836_preds(0) <= place_1283_token;
  transition_836_preds(1) <= place_1295_token;
  transition_836 : transition
    port map(
      preds      => transition_836_preds,
      symbol_out => transition_836_symbol_out,
      symbol_in  => true);

  transition_837_preds(0) <= place_1299_token;
  LambdaOut(228) <= transition_837_symbol_out;
  transition_837 : transition
    port map(
      preds      => transition_837_preds,
      symbol_out => transition_837_symbol_out,
      symbol_in  => true);

  transition_838_preds(0) <= place_841_token;
  transition_838 : transition
    port map(
      preds      => transition_838_preds,
      symbol_out => transition_838_symbol_out,
      symbol_in  => LambdaIn(226));

  transition_839_preds(0) <= place_842_token;
  LambdaOut(229) <= transition_839_symbol_out;
  transition_839 : transition
    port map(
      preds      => transition_839_preds,
      symbol_out => transition_839_symbol_out,
      symbol_in  => true);

  transition_840_preds(0) <= place_843_token;
  transition_840 : transition
    port map(
      preds      => transition_840_preds,
      symbol_out => transition_840_symbol_out,
      symbol_in  => LambdaIn(227));

  transition_844_preds(0) <= place_1302_token;
  LambdaOut(230) <= transition_844_symbol_out;
  transition_844 : transition
    port map(
      preds      => transition_844_preds,
      symbol_out => transition_844_symbol_out,
      symbol_in  => true);

  transition_845_preds(0) <= place_848_token;
  transition_845 : transition
    port map(
      preds      => transition_845_preds,
      symbol_out => transition_845_symbol_out,
      symbol_in  => LambdaIn(228));

  transition_846_preds(0) <= place_849_token;
  LambdaOut(231) <= transition_846_symbol_out;
  transition_846 : transition
    port map(
      preds      => transition_846_preds,
      symbol_out => transition_846_symbol_out,
      symbol_in  => true);

  transition_847_preds(0) <= place_850_token;
  transition_847 : transition
    port map(
      preds      => transition_847_preds,
      symbol_out => transition_847_symbol_out,
      symbol_in  => LambdaIn(229));

  transition_851_preds(0) <= place_1303_token;
  LambdaOut(232) <= transition_851_symbol_out;
  transition_851 : transition
    port map(
      preds      => transition_851_preds,
      symbol_out => transition_851_symbol_out,
      symbol_in  => true);

  transition_852_preds(0) <= place_855_token;
  transition_852 : transition
    port map(
      preds      => transition_852_preds,
      symbol_out => transition_852_symbol_out,
      symbol_in  => LambdaIn(230));

  transition_853_preds(0) <= place_856_token;
  LambdaOut(233) <= transition_853_symbol_out;
  transition_853 : transition
    port map(
      preds      => transition_853_preds,
      symbol_out => transition_853_symbol_out,
      symbol_in  => true);

  transition_854_preds(0) <= place_857_token;
  transition_854 : transition
    port map(
      preds      => transition_854_preds,
      symbol_out => transition_854_symbol_out,
      symbol_in  => LambdaIn(231));

  transition_858_preds(0) <= place_1298_token;
  transition_858_preds(1) <= place_1301_token;
  transition_858 : transition
    port map(
      preds      => transition_858_preds,
      symbol_out => transition_858_symbol_out,
      symbol_in  => true);

  transition_859_preds(0) <= place_1306_token;
  LambdaOut(234) <= transition_859_symbol_out;
  transition_859 : transition
    port map(
      preds      => transition_859_preds,
      symbol_out => transition_859_symbol_out,
      symbol_in  => true);

  transition_860_preds(0) <= place_863_token;
  transition_860 : transition
    port map(
      preds      => transition_860_preds,
      symbol_out => transition_860_symbol_out,
      symbol_in  => LambdaIn(232));

  transition_861_preds(0) <= place_864_token;
  LambdaOut(235) <= transition_861_symbol_out;
  transition_861 : transition
    port map(
      preds      => transition_861_preds,
      symbol_out => transition_861_symbol_out,
      symbol_in  => true);

  transition_862_preds(0) <= place_865_token;
  transition_862 : transition
    port map(
      preds      => transition_862_preds,
      symbol_out => transition_862_symbol_out,
      symbol_in  => LambdaIn(233));

  transition_866_preds(0) <= place_1307_token;
  LambdaOut(236) <= transition_866_symbol_out;
  transition_866 : transition
    port map(
      preds      => transition_866_preds,
      symbol_out => transition_866_symbol_out,
      symbol_in  => true);

  transition_867_preds(0) <= place_870_token;
  transition_867 : transition
    port map(
      preds      => transition_867_preds,
      symbol_out => transition_867_symbol_out,
      symbol_in  => LambdaIn(234));

  transition_868_preds(0) <= place_871_token;
  LambdaOut(237) <= transition_868_symbol_out;
  transition_868 : transition
    port map(
      preds      => transition_868_preds,
      symbol_out => transition_868_symbol_out,
      symbol_in  => true);

  transition_869_preds(0) <= place_872_token;
  transition_869 : transition
    port map(
      preds      => transition_869_preds,
      symbol_out => transition_869_symbol_out,
      symbol_in  => LambdaIn(235));

  transition_873_preds(0) <= place_1304_token;
  transition_873_preds(1) <= place_1305_token;
  transition_873 : transition
    port map(
      preds      => transition_873_preds,
      symbol_out => transition_873_symbol_out,
      symbol_in  => true);

  transition_874_preds(0) <= place_1308_token;
  LambdaOut(238) <= transition_874_symbol_out;
  transition_874 : transition
    port map(
      preds      => transition_874_preds,
      symbol_out => transition_874_symbol_out,
      symbol_in  => true);

  transition_875_preds(0) <= place_878_token;
  transition_875 : transition
    port map(
      preds      => transition_875_preds,
      symbol_out => transition_875_symbol_out,
      symbol_in  => LambdaIn(236));

  transition_876_preds(0) <= place_879_token;
  LambdaOut(239) <= transition_876_symbol_out;
  transition_876 : transition
    port map(
      preds      => transition_876_preds,
      symbol_out => transition_876_symbol_out,
      symbol_in  => true);

  transition_877_preds(0) <= place_880_token;
  transition_877 : transition
    port map(
      preds      => transition_877_preds,
      symbol_out => transition_877_symbol_out,
      symbol_in  => LambdaIn(237));

  transition_882_preds(0) <= place_881_token;
  transition_882 : transition
    port map(
      preds      => transition_882_preds,
      symbol_out => transition_882_symbol_out,
      symbol_in  => LambdaIn(238));

  transition_883_preds(0) <= place_1311_token;
  LambdaOut(240) <= transition_883_symbol_out;
  transition_883 : transition
    port map(
      preds      => transition_883_preds,
      symbol_out => transition_883_symbol_out,
      symbol_in  => true);

  transition_884_preds(0) <= place_1297_token;
  transition_884_preds(1) <= place_1309_token;
  transition_884 : transition
    port map(
      preds      => transition_884_preds,
      symbol_out => transition_884_symbol_out,
      symbol_in  => true);

  transition_885_preds(0) <= place_1314_token;
  LambdaOut(241) <= transition_885_symbol_out;
  transition_885 : transition
    port map(
      preds      => transition_885_preds,
      symbol_out => transition_885_symbol_out,
      symbol_in  => true);

  transition_886_preds(0) <= place_889_token;
  transition_886 : transition
    port map(
      preds      => transition_886_preds,
      symbol_out => transition_886_symbol_out,
      symbol_in  => LambdaIn(239));

  transition_887_preds(0) <= place_890_token;
  LambdaOut(242) <= transition_887_symbol_out;
  transition_887 : transition
    port map(
      preds      => transition_887_preds,
      symbol_out => transition_887_symbol_out,
      symbol_in  => true);

  transition_888_preds(0) <= place_891_token;
  transition_888 : transition
    port map(
      preds      => transition_888_preds,
      symbol_out => transition_888_symbol_out,
      symbol_in  => LambdaIn(240));

  transition_892_preds(0) <= place_1316_token;
  LambdaOut(243) <= transition_892_symbol_out;
  transition_892 : transition
    port map(
      preds      => transition_892_preds,
      symbol_out => transition_892_symbol_out,
      symbol_in  => true);

  transition_893_preds(0) <= place_896_token;
  transition_893 : transition
    port map(
      preds      => transition_893_preds,
      symbol_out => transition_893_symbol_out,
      symbol_in  => LambdaIn(241));

  transition_894_preds(0) <= place_897_token;
  LambdaOut(244) <= transition_894_symbol_out;
  transition_894 : transition
    port map(
      preds      => transition_894_preds,
      symbol_out => transition_894_symbol_out,
      symbol_in  => true);

  transition_895_preds(0) <= place_898_token;
  transition_895 : transition
    port map(
      preds      => transition_895_preds,
      symbol_out => transition_895_symbol_out,
      symbol_in  => LambdaIn(242));

  transition_899_preds(0) <= place_1317_token;
  LambdaOut(245) <= transition_899_symbol_out;
  transition_899 : transition
    port map(
      preds      => transition_899_preds,
      symbol_out => transition_899_symbol_out,
      symbol_in  => true);

  transition_900_preds(0) <= place_903_token;
  transition_900 : transition
    port map(
      preds      => transition_900_preds,
      symbol_out => transition_900_symbol_out,
      symbol_in  => LambdaIn(243));

  transition_901_preds(0) <= place_904_token;
  LambdaOut(246) <= transition_901_symbol_out;
  transition_901 : transition
    port map(
      preds      => transition_901_preds,
      symbol_out => transition_901_symbol_out,
      symbol_in  => true);

  transition_902_preds(0) <= place_905_token;
  transition_902 : transition
    port map(
      preds      => transition_902_preds,
      symbol_out => transition_902_symbol_out,
      symbol_in  => LambdaIn(244));

  transition_906_preds(0) <= place_1315_token;
  transition_906_preds(1) <= place_1313_token;
  transition_906 : transition
    port map(
      preds      => transition_906_preds,
      symbol_out => transition_906_symbol_out,
      symbol_in  => true);

  transition_907_preds(0) <= place_1321_token;
  LambdaOut(247) <= transition_907_symbol_out;
  transition_907 : transition
    port map(
      preds      => transition_907_preds,
      symbol_out => transition_907_symbol_out,
      symbol_in  => true);

  transition_908_preds(0) <= place_911_token;
  transition_908 : transition
    port map(
      preds      => transition_908_preds,
      symbol_out => transition_908_symbol_out,
      symbol_in  => LambdaIn(245));

  transition_909_preds(0) <= place_912_token;
  LambdaOut(248) <= transition_909_symbol_out;
  transition_909 : transition
    port map(
      preds      => transition_909_preds,
      symbol_out => transition_909_symbol_out,
      symbol_in  => true);

  transition_910_preds(0) <= place_913_token;
  transition_910 : transition
    port map(
      preds      => transition_910_preds,
      symbol_out => transition_910_symbol_out,
      symbol_in  => LambdaIn(246));

  transition_914_preds(0) <= place_1322_token;
  LambdaOut(249) <= transition_914_symbol_out;
  transition_914 : transition
    port map(
      preds      => transition_914_preds,
      symbol_out => transition_914_symbol_out,
      symbol_in  => true);

  transition_915_preds(0) <= place_918_token;
  transition_915 : transition
    port map(
      preds      => transition_915_preds,
      symbol_out => transition_915_symbol_out,
      symbol_in  => LambdaIn(247));

  transition_916_preds(0) <= place_919_token;
  LambdaOut(250) <= transition_916_symbol_out;
  transition_916 : transition
    port map(
      preds      => transition_916_preds,
      symbol_out => transition_916_symbol_out,
      symbol_in  => true);

  transition_917_preds(0) <= place_920_token;
  transition_917 : transition
    port map(
      preds      => transition_917_preds,
      symbol_out => transition_917_symbol_out,
      symbol_in  => LambdaIn(248));

  transition_921_preds(0) <= place_1320_token;
  transition_921_preds(1) <= place_1318_token;
  transition_921 : transition
    port map(
      preds      => transition_921_preds,
      symbol_out => transition_921_symbol_out,
      symbol_in  => true);

  transition_922_preds(0) <= place_1323_token;
  LambdaOut(251) <= transition_922_symbol_out;
  transition_922 : transition
    port map(
      preds      => transition_922_preds,
      symbol_out => transition_922_symbol_out,
      symbol_in  => true);

  transition_923_preds(0) <= place_926_token;
  transition_923 : transition
    port map(
      preds      => transition_923_preds,
      symbol_out => transition_923_symbol_out,
      symbol_in  => LambdaIn(249));

  transition_924_preds(0) <= place_927_token;
  LambdaOut(252) <= transition_924_symbol_out;
  transition_924 : transition
    port map(
      preds      => transition_924_preds,
      symbol_out => transition_924_symbol_out,
      symbol_in  => true);

  transition_925_preds(0) <= place_928_token;
  transition_925 : transition
    port map(
      preds      => transition_925_preds,
      symbol_out => transition_925_symbol_out,
      symbol_in  => LambdaIn(250));

  transition_930_preds(0) <= place_929_token;
  transition_930 : transition
    port map(
      preds      => transition_930_preds,
      symbol_out => transition_930_symbol_out,
      symbol_in  => LambdaIn(251));

  transition_931_preds(0) <= place_1326_token;
  LambdaOut(253) <= transition_931_symbol_out;
  transition_931 : transition
    port map(
      preds      => transition_931_preds,
      symbol_out => transition_931_symbol_out,
      symbol_in  => true);

  transition_932_preds(0) <= place_1312_token;
  transition_932_preds(1) <= place_1325_token;
  transition_932 : transition
    port map(
      preds      => transition_932_preds,
      symbol_out => transition_932_symbol_out,
      symbol_in  => true);

  transition_933_preds(0) <= place_1330_token;
  LambdaOut(254) <= transition_933_symbol_out;
  transition_933 : transition
    port map(
      preds      => transition_933_preds,
      symbol_out => transition_933_symbol_out,
      symbol_in  => true);

  transition_934_preds(0) <= place_937_token;
  transition_934 : transition
    port map(
      preds      => transition_934_preds,
      symbol_out => transition_934_symbol_out,
      symbol_in  => LambdaIn(252));

  transition_935_preds(0) <= place_938_token;
  LambdaOut(255) <= transition_935_symbol_out;
  transition_935 : transition
    port map(
      preds      => transition_935_preds,
      symbol_out => transition_935_symbol_out,
      symbol_in  => true);

  transition_936_preds(0) <= place_939_token;
  transition_936 : transition
    port map(
      preds      => transition_936_preds,
      symbol_out => transition_936_symbol_out,
      symbol_in  => LambdaIn(253));

  transition_940_preds(0) <= place_1332_token;
  LambdaOut(256) <= transition_940_symbol_out;
  transition_940 : transition
    port map(
      preds      => transition_940_preds,
      symbol_out => transition_940_symbol_out,
      symbol_in  => true);

  transition_941_preds(0) <= place_944_token;
  transition_941 : transition
    port map(
      preds      => transition_941_preds,
      symbol_out => transition_941_symbol_out,
      symbol_in  => LambdaIn(254));

  transition_942_preds(0) <= place_945_token;
  LambdaOut(257) <= transition_942_symbol_out;
  transition_942 : transition
    port map(
      preds      => transition_942_preds,
      symbol_out => transition_942_symbol_out,
      symbol_in  => true);

  transition_943_preds(0) <= place_946_token;
  transition_943 : transition
    port map(
      preds      => transition_943_preds,
      symbol_out => transition_943_symbol_out,
      symbol_in  => LambdaIn(255));

  transition_947_preds(0) <= place_1333_token;
  LambdaOut(258) <= transition_947_symbol_out;
  transition_947 : transition
    port map(
      preds      => transition_947_preds,
      symbol_out => transition_947_symbol_out,
      symbol_in  => true);

  transition_948_preds(0) <= place_951_token;
  transition_948 : transition
    port map(
      preds      => transition_948_preds,
      symbol_out => transition_948_symbol_out,
      symbol_in  => LambdaIn(256));

  transition_949_preds(0) <= place_952_token;
  LambdaOut(259) <= transition_949_symbol_out;
  transition_949 : transition
    port map(
      preds      => transition_949_preds,
      symbol_out => transition_949_symbol_out,
      symbol_in  => true);

  transition_950_preds(0) <= place_953_token;
  transition_950 : transition
    port map(
      preds      => transition_950_preds,
      symbol_out => transition_950_symbol_out,
      symbol_in  => LambdaIn(257));

  transition_954_preds(0) <= place_1328_token;
  transition_954_preds(1) <= place_1331_token;
  transition_954 : transition
    port map(
      preds      => transition_954_preds,
      symbol_out => transition_954_symbol_out,
      symbol_in  => true);

  transition_955_preds(0) <= place_1336_token;
  LambdaOut(260) <= transition_955_symbol_out;
  transition_955 : transition
    port map(
      preds      => transition_955_preds,
      symbol_out => transition_955_symbol_out,
      symbol_in  => true);

  transition_956_preds(0) <= place_959_token;
  transition_956 : transition
    port map(
      preds      => transition_956_preds,
      symbol_out => transition_956_symbol_out,
      symbol_in  => LambdaIn(258));

  transition_957_preds(0) <= place_960_token;
  LambdaOut(261) <= transition_957_symbol_out;
  transition_957 : transition
    port map(
      preds      => transition_957_preds,
      symbol_out => transition_957_symbol_out,
      symbol_in  => true);

  transition_958_preds(0) <= place_961_token;
  transition_958 : transition
    port map(
      preds      => transition_958_preds,
      symbol_out => transition_958_symbol_out,
      symbol_in  => LambdaIn(259));

  transition_962_preds(0) <= place_1337_token;
  LambdaOut(262) <= transition_962_symbol_out;
  transition_962 : transition
    port map(
      preds      => transition_962_preds,
      symbol_out => transition_962_symbol_out,
      symbol_in  => true);

  transition_963_preds(0) <= place_966_token;
  transition_963 : transition
    port map(
      preds      => transition_963_preds,
      symbol_out => transition_963_symbol_out,
      symbol_in  => LambdaIn(260));

  transition_964_preds(0) <= place_967_token;
  LambdaOut(263) <= transition_964_symbol_out;
  transition_964 : transition
    port map(
      preds      => transition_964_preds,
      symbol_out => transition_964_symbol_out,
      symbol_in  => true);

  transition_965_preds(0) <= place_968_token;
  transition_965 : transition
    port map(
      preds      => transition_965_preds,
      symbol_out => transition_965_symbol_out,
      symbol_in  => LambdaIn(261));

  transition_969_preds(0) <= place_1334_token;
  transition_969_preds(1) <= place_1335_token;
  transition_969 : transition
    port map(
      preds      => transition_969_preds,
      symbol_out => transition_969_symbol_out,
      symbol_in  => true);

  transition_970_preds(0) <= place_1338_token;
  LambdaOut(264) <= transition_970_symbol_out;
  transition_970 : transition
    port map(
      preds      => transition_970_preds,
      symbol_out => transition_970_symbol_out,
      symbol_in  => true);

  transition_971_preds(0) <= place_974_token;
  transition_971 : transition
    port map(
      preds      => transition_971_preds,
      symbol_out => transition_971_symbol_out,
      symbol_in  => LambdaIn(262));

  transition_972_preds(0) <= place_975_token;
  LambdaOut(265) <= transition_972_symbol_out;
  transition_972 : transition
    port map(
      preds      => transition_972_preds,
      symbol_out => transition_972_symbol_out,
      symbol_in  => true);

  transition_973_preds(0) <= place_976_token;
  transition_973 : transition
    port map(
      preds      => transition_973_preds,
      symbol_out => transition_973_symbol_out,
      symbol_in  => LambdaIn(263));

  transition_978_preds(0) <= place_977_token;
  transition_978 : transition
    port map(
      preds      => transition_978_preds,
      symbol_out => transition_978_symbol_out,
      symbol_in  => LambdaIn(264));

  transition_979_preds(0) <= place_1340_token;
  LambdaOut(266) <= transition_979_symbol_out;
  transition_979 : transition
    port map(
      preds      => transition_979_preds,
      symbol_out => transition_979_symbol_out,
      symbol_in  => true);

  transition_980_preds(0) <= place_1327_token;
  transition_980_preds(1) <= place_1339_token;
  transition_980 : transition
    port map(
      preds      => transition_980_preds,
      symbol_out => transition_980_symbol_out,
      symbol_in  => true);

  transition_981_preds(0) <= place_1343_token;
  LambdaOut(267) <= transition_981_symbol_out;
  transition_981 : transition
    port map(
      preds      => transition_981_preds,
      symbol_out => transition_981_symbol_out,
      symbol_in  => true);

  transition_982_preds(0) <= place_985_token;
  transition_982 : transition
    port map(
      preds      => transition_982_preds,
      symbol_out => transition_982_symbol_out,
      symbol_in  => LambdaIn(265));

  transition_983_preds(0) <= place_986_token;
  LambdaOut(268) <= transition_983_symbol_out;
  transition_983 : transition
    port map(
      preds      => transition_983_preds,
      symbol_out => transition_983_symbol_out,
      symbol_in  => true);

  transition_984_preds(0) <= place_987_token;
  transition_984 : transition
    port map(
      preds      => transition_984_preds,
      symbol_out => transition_984_symbol_out,
      symbol_in  => LambdaIn(266));

  transition_988_preds(0) <= place_1345_token;
  LambdaOut(269) <= transition_988_symbol_out;
  transition_988 : transition
    port map(
      preds      => transition_988_preds,
      symbol_out => transition_988_symbol_out,
      symbol_in  => true);

  transition_989_preds(0) <= place_992_token;
  transition_989 : transition
    port map(
      preds      => transition_989_preds,
      symbol_out => transition_989_symbol_out,
      symbol_in  => LambdaIn(267));

  transition_990_preds(0) <= place_993_token;
  LambdaOut(270) <= transition_990_symbol_out;
  transition_990 : transition
    port map(
      preds      => transition_990_preds,
      symbol_out => transition_990_symbol_out,
      symbol_in  => true);

  transition_991_preds(0) <= place_994_token;
  transition_991 : transition
    port map(
      preds      => transition_991_preds,
      symbol_out => transition_991_symbol_out,
      symbol_in  => LambdaIn(268));

  transition_995_preds(0) <= place_1346_token;
  LambdaOut(271) <= transition_995_symbol_out;
  transition_995 : transition
    port map(
      preds      => transition_995_preds,
      symbol_out => transition_995_symbol_out,
      symbol_in  => true);

  transition_996_preds(0) <= place_999_token;
  transition_996 : transition
    port map(
      preds      => transition_996_preds,
      symbol_out => transition_996_symbol_out,
      symbol_in  => LambdaIn(269));

  transition_997_preds(0) <= place_1000_token;
  LambdaOut(272) <= transition_997_symbol_out;
  transition_997 : transition
    port map(
      preds      => transition_997_preds,
      symbol_out => transition_997_symbol_out,
      symbol_in  => true);

  transition_998_preds(0) <= place_1001_token;
  transition_998 : transition
    port map(
      preds      => transition_998_preds,
      symbol_out => transition_998_symbol_out,
      symbol_in  => LambdaIn(270));

  transition_1002_preds(0) <= place_1344_token;
  transition_1002_preds(1) <= place_1342_token;
  transition_1002 : transition
    port map(
      preds      => transition_1002_preds,
      symbol_out => transition_1002_symbol_out,
      symbol_in  => true);

  transition_1003_preds(0) <= place_1349_token;
  LambdaOut(273) <= transition_1003_symbol_out;
  transition_1003 : transition
    port map(
      preds      => transition_1003_preds,
      symbol_out => transition_1003_symbol_out,
      symbol_in  => true);

  transition_1004_preds(0) <= place_1007_token;
  transition_1004 : transition
    port map(
      preds      => transition_1004_preds,
      symbol_out => transition_1004_symbol_out,
      symbol_in  => LambdaIn(271));

  transition_1005_preds(0) <= place_1008_token;
  LambdaOut(274) <= transition_1005_symbol_out;
  transition_1005 : transition
    port map(
      preds      => transition_1005_preds,
      symbol_out => transition_1005_symbol_out,
      symbol_in  => true);

  transition_1006_preds(0) <= place_1009_token;
  transition_1006 : transition
    port map(
      preds      => transition_1006_preds,
      symbol_out => transition_1006_symbol_out,
      symbol_in  => LambdaIn(272));

  transition_1010_preds(0) <= place_1350_token;
  LambdaOut(275) <= transition_1010_symbol_out;
  transition_1010 : transition
    port map(
      preds      => transition_1010_preds,
      symbol_out => transition_1010_symbol_out,
      symbol_in  => true);

  transition_1011_preds(0) <= place_1014_token;
  transition_1011 : transition
    port map(
      preds      => transition_1011_preds,
      symbol_out => transition_1011_symbol_out,
      symbol_in  => LambdaIn(273));

  transition_1012_preds(0) <= place_1015_token;
  LambdaOut(276) <= transition_1012_symbol_out;
  transition_1012 : transition
    port map(
      preds      => transition_1012_preds,
      symbol_out => transition_1012_symbol_out,
      symbol_in  => true);

  transition_1013_preds(0) <= place_1016_token;
  transition_1013 : transition
    port map(
      preds      => transition_1013_preds,
      symbol_out => transition_1013_symbol_out,
      symbol_in  => LambdaIn(274));

  transition_1017_preds(0) <= place_1347_token;
  transition_1017_preds(1) <= place_1348_token;
  transition_1017 : transition
    port map(
      preds      => transition_1017_preds,
      symbol_out => transition_1017_symbol_out,
      symbol_in  => true);

  transition_1018_preds(0) <= place_1351_token;
  LambdaOut(277) <= transition_1018_symbol_out;
  transition_1018 : transition
    port map(
      preds      => transition_1018_preds,
      symbol_out => transition_1018_symbol_out,
      symbol_in  => true);

  transition_1019_preds(0) <= place_1022_token;
  transition_1019 : transition
    port map(
      preds      => transition_1019_preds,
      symbol_out => transition_1019_symbol_out,
      symbol_in  => LambdaIn(275));

  transition_1020_preds(0) <= place_1023_token;
  LambdaOut(278) <= transition_1020_symbol_out;
  transition_1020 : transition
    port map(
      preds      => transition_1020_preds,
      symbol_out => transition_1020_symbol_out,
      symbol_in  => true);

  transition_1021_preds(0) <= place_1024_token;
  transition_1021 : transition
    port map(
      preds      => transition_1021_preds,
      symbol_out => transition_1021_symbol_out,
      symbol_in  => LambdaIn(276));

  transition_1026_preds(0) <= place_1025_token;
  transition_1026 : transition
    port map(
      preds      => transition_1026_preds,
      symbol_out => transition_1026_symbol_out,
      symbol_in  => LambdaIn(277));

  transition_1027_preds(0) <= place_1354_token;
  LambdaOut(279) <= transition_1027_symbol_out;
  transition_1027 : transition
    port map(
      preds      => transition_1027_preds,
      symbol_out => transition_1027_symbol_out,
      symbol_in  => true);

  transition_1028_preds(0) <= place_1341_token;
  transition_1028_preds(1) <= place_1353_token;
  transition_1028 : transition
    port map(
      preds      => transition_1028_preds,
      symbol_out => transition_1028_symbol_out,
      symbol_in  => true);

  transition_1030_preds(0) <= place_1029_token;
  transition_1030 : transition
    port map(
      preds      => transition_1030_preds,
      symbol_out => transition_1030_symbol_out,
      symbol_in  => LambdaIn(278));

  transition_1031_preds(0) <= place_1355_token;
  LambdaOut(280) <= transition_1031_symbol_out;
  transition_1031 : transition
    port map(
      preds      => transition_1031_preds,
      symbol_out => transition_1031_symbol_out,
      symbol_in  => true);

  transition_1033_preds(0) <= place_1032_token;
  transition_1033 : transition
    port map(
      preds      => transition_1033_preds,
      symbol_out => transition_1033_symbol_out,
      symbol_in  => LambdaIn(279));

  transition_1034_preds(0) <= place_1356_token;
  LambdaOut(281) <= transition_1034_symbol_out;
  transition_1034 : transition
    port map(
      preds      => transition_1034_preds,
      symbol_out => transition_1034_symbol_out,
      symbol_in  => true);

  transition_1035_preds(0) <= place_1357_token;
  transition_1035 : transition
    port map(
      preds      => transition_1035_preds,
      symbol_out => transition_1035_symbol_out,
      symbol_in  => true);

  transition_1037_preds(0) <= place_1036_token;
  transition_1037 : transition
    port map(
      preds      => transition_1037_preds,
      symbol_out => transition_1037_symbol_out,
      symbol_in  => LambdaIn(280));

  transition_1038_preds(0) <= place_1361_token;
  LambdaOut(282) <= transition_1038_symbol_out;
  transition_1038 : transition
    port map(
      preds      => transition_1038_preds,
      symbol_out => transition_1038_symbol_out,
      symbol_in  => true);

  transition_1040_preds(0) <= place_1039_token;
  transition_1040 : transition
    port map(
      preds      => transition_1040_preds,
      symbol_out => transition_1040_symbol_out,
      symbol_in  => LambdaIn(281));

  transition_1041_preds(0) <= place_1358_token;
  LambdaOut(283) <= transition_1041_symbol_out;
  transition_1041 : transition
    port map(
      preds      => transition_1041_preds,
      symbol_out => transition_1041_symbol_out,
      symbol_in  => true);

  transition_1042_preds(0) <= place_1360_token;
  transition_1042 : transition
    port map(
      preds      => transition_1042_preds,
      symbol_out => transition_1042_symbol_out,
      symbol_in  => true);

  transition_1043_preds(0) <= place_1363_token;
  LambdaOut(284) <= transition_1043_symbol_out;
  transition_1043 : transition
    port map(
      preds      => transition_1043_preds,
      symbol_out => transition_1043_symbol_out,
      symbol_in  => true);

  transition_1044_preds(0) <= place_1047_token;
  transition_1044 : transition
    port map(
      preds      => transition_1044_preds,
      symbol_out => transition_1044_symbol_out,
      symbol_in  => LambdaIn(282));

  transition_1045_preds(0) <= place_1048_token;
  LambdaOut(285) <= transition_1045_symbol_out;
  transition_1045 : transition
    port map(
      preds      => transition_1045_preds,
      symbol_out => transition_1045_symbol_out,
      symbol_in  => true);

  transition_1046_preds(0) <= place_1049_token;
  transition_1046 : transition
    port map(
      preds      => transition_1046_preds,
      symbol_out => transition_1046_symbol_out,
      symbol_in  => LambdaIn(283));

  transition_1051_preds(0) <= place_1050_token;
  transition_1051 : transition
    port map(
      preds      => transition_1051_preds,
      symbol_out => transition_1051_symbol_out,
      symbol_in  => LambdaIn(284));

  transition_1052_preds(0) <= place_1368_token;
  LambdaOut(286) <= transition_1052_symbol_out;
  transition_1052 : transition
    port map(
      preds      => transition_1052_preds,
      symbol_out => transition_1052_symbol_out,
      symbol_in  => true);

  transition_1054_preds(0) <= place_1053_token;
  transition_1054 : transition
    port map(
      preds      => transition_1054_preds,
      symbol_out => transition_1054_symbol_out,
      symbol_in  => LambdaIn(285));

  transition_1055_preds(0) <= place_1364_token;
  LambdaOut(287) <= transition_1055_symbol_out;
  transition_1055 : transition
    port map(
      preds      => transition_1055_preds,
      symbol_out => transition_1055_symbol_out,
      symbol_in  => true);

  transition_1056_preds(0) <= place_1367_token;
  LambdaOut(288) <= transition_1056_symbol_out;
  transition_1056 : transition
    port map(
      preds      => transition_1056_preds,
      symbol_out => transition_1056_symbol_out,
      symbol_in  => true);

  transition_1057_preds(0) <= place_1060_token;
  transition_1057 : transition
    port map(
      preds      => transition_1057_preds,
      symbol_out => transition_1057_symbol_out,
      symbol_in  => LambdaIn(286));

  transition_1058_preds(0) <= place_1061_token;
  LambdaOut(289) <= transition_1058_symbol_out;
  transition_1058 : transition
    port map(
      preds      => transition_1058_preds,
      symbol_out => transition_1058_symbol_out,
      symbol_in  => true);

  transition_1059_preds(0) <= place_1062_token;
  transition_1059 : transition
    port map(
      preds      => transition_1059_preds,
      symbol_out => transition_1059_symbol_out,
      symbol_in  => LambdaIn(287));

  transition_1063_preds(0) <= place_1370_token;
  LambdaOut(290) <= transition_1063_symbol_out;
  transition_1063 : transition
    port map(
      preds      => transition_1063_preds,
      symbol_out => transition_1063_symbol_out,
      symbol_in  => true);

  transition_1064_preds(0) <= place_1067_token;
  transition_1064 : transition
    port map(
      preds      => transition_1064_preds,
      symbol_out => transition_1064_symbol_out,
      symbol_in  => LambdaIn(288));

  transition_1065_preds(0) <= place_1068_token;
  LambdaOut(291) <= transition_1065_symbol_out;
  transition_1065 : transition
    port map(
      preds      => transition_1065_preds,
      symbol_out => transition_1065_symbol_out,
      symbol_in  => true);

  transition_1066_preds(0) <= place_1069_token;
  transition_1066 : transition
    port map(
      preds      => transition_1066_preds,
      symbol_out => transition_1066_symbol_out,
      symbol_in  => LambdaIn(289));

  transition_1070_preds(0) <= place_1362_token;
  transition_1070_preds(1) <= place_1373_token;
  transition_1070 : transition
    port map(
      preds      => transition_1070_preds,
      symbol_out => transition_1070_symbol_out,
      symbol_in  => true);

  transition_1071_preds(0) <= place_1374_token;
  LambdaOut(292) <= transition_1071_symbol_out;
  transition_1071 : transition
    port map(
      preds      => transition_1071_preds,
      symbol_out => transition_1071_symbol_out,
      symbol_in  => true);

  transition_1072_preds(0) <= place_1075_token;
  transition_1072 : transition
    port map(
      preds      => transition_1072_preds,
      symbol_out => transition_1072_symbol_out,
      symbol_in  => LambdaIn(290));

  transition_1073_preds(0) <= place_1076_token;
  LambdaOut(293) <= transition_1073_symbol_out;
  transition_1073 : transition
    port map(
      preds      => transition_1073_preds,
      symbol_out => transition_1073_symbol_out,
      symbol_in  => true);

  transition_1074_preds(0) <= place_1077_token;
  transition_1074 : transition
    port map(
      preds      => transition_1074_preds,
      symbol_out => transition_1074_symbol_out,
      symbol_in  => LambdaIn(291));

  transition_1078_preds(0) <= place_1369_token;
  transition_1078_preds(1) <= place_1372_token;
  transition_1078 : transition
    port map(
      preds      => transition_1078_preds,
      symbol_out => transition_1078_symbol_out,
      symbol_in  => true);

  transition_1080_preds(0) <= place_1079_token;
  transition_1080 : transition
    port map(
      preds      => transition_1080_preds,
      symbol_out => transition_1080_symbol_out,
      symbol_in  => LambdaIn(292));

  transition_1081_preds(0) <= place_1375_token;
  LambdaOut(294) <= transition_1081_symbol_out;
  transition_1081 : transition
    port map(
      preds      => transition_1081_preds,
      symbol_out => transition_1081_symbol_out,
      symbol_in  => true);

end architecture default_arch;