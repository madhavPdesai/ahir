-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant foo_base_address : std_logic_vector(3 downto 0) := "0000";
  constant free_queue_base_address : std_logic_vector(2 downto 0) := "000";
  constant free_queue_ram_base_address : std_logic_vector(10 downto 0) := "00000000000";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  constant xx_xstr10_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr11_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr12_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr1_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr2_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr3_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr4_base_address : std_logic_vector(4 downto 0) := "00000";
  constant xx_xstr5_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr6_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr7_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr8_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr9_base_address : std_logic_vector(3 downto 0) := "0000";
  constant xx_xstr_base_address : std_logic_vector(3 downto 0) := "0000";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_manager is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
    free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity free_queue_manager;
architecture Default of free_queue_manager is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal free_queue_manager_CP_3612_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_879_offset_inst_ack_0 : boolean;
  signal ptr_deref_805_store_0_req_1 : boolean;
  signal switch_stmt_842_select_expr_1_req_0 : boolean;
  signal ptr_deref_794_gather_scatter_req_0 : boolean;
  signal ptr_deref_805_store_0_ack_1 : boolean;
  signal ptr_deref_794_gather_scatter_ack_0 : boolean;
  signal ptr_deref_794_store_0_req_0 : boolean;
  signal ptr_deref_805_gather_scatter_ack_0 : boolean;
  signal ptr_deref_805_store_0_ack_0 : boolean;
  signal ptr_deref_805_gather_scatter_req_0 : boolean;
  signal ptr_deref_827_store_0_req_0 : boolean;
  signal switch_stmt_842_branch_0_ack_1 : boolean;
  signal ptr_deref_805_store_0_req_0 : boolean;
  signal ptr_deref_816_gather_scatter_ack_0 : boolean;
  signal ptr_deref_827_store_0_req_1 : boolean;
  signal ptr_deref_827_store_0_ack_1 : boolean;
  signal switch_stmt_842_select_expr_1_ack_1 : boolean;
  signal switch_stmt_842_select_expr_1_req_1 : boolean;
  signal ptr_deref_827_store_0_ack_0 : boolean;
  signal simple_obj_ref_840_inst_req_0 : boolean;
  signal simple_obj_ref_840_inst_ack_0 : boolean;
  signal if_stmt_870_branch_ack_1 : boolean;
  signal ptr_deref_816_store_0_ack_0 : boolean;
  signal switch_stmt_842_select_expr_0_req_0 : boolean;
  signal ptr_deref_794_store_0_ack_0 : boolean;
  signal switch_stmt_842_select_expr_0_ack_0 : boolean;
  signal ptr_deref_816_store_0_req_1 : boolean;
  signal ptr_deref_816_gather_scatter_req_0 : boolean;
  signal ptr_deref_816_store_0_req_0 : boolean;
  signal array_obj_ref_879_index_0_rename_ack_0 : boolean;
  signal ptr_deref_816_store_0_ack_1 : boolean;
  signal binary_868_inst_ack_1 : boolean;
  signal ptr_deref_884_addr_0_req_0 : boolean;
  signal ptr_deref_884_gather_scatter_ack_0 : boolean;
  signal switch_stmt_842_branch_1_req_0 : boolean;
  signal binary_868_inst_req_1 : boolean;
  signal ptr_deref_794_store_0_ack_1 : boolean;
  signal ptr_deref_794_store_0_req_1 : boolean;
  signal switch_stmt_842_branch_default_req_0 : boolean;
  signal ptr_deref_884_root_address_inst_ack_0 : boolean;
  signal switch_stmt_842_select_expr_1_ack_0 : boolean;
  signal binary_868_inst_ack_0 : boolean;
  signal array_obj_ref_879_root_address_inst_ack_0 : boolean;
  signal ptr_deref_884_load_0_req_0 : boolean;
  signal ptr_deref_884_load_0_ack_1 : boolean;
  signal ptr_deref_884_root_address_inst_req_0 : boolean;
  signal switch_stmt_842_select_expr_0_req_1 : boolean;
  signal binary_890_inst_ack_0 : boolean;
  signal ptr_deref_884_load_0_ack_0 : boolean;
  signal if_stmt_870_branch_ack_0 : boolean;
  signal array_obj_ref_879_index_0_resize_req_0 : boolean;
  signal ptr_deref_884_addr_0_ack_0 : boolean;
  signal ptr_deref_884_base_resize_req_0 : boolean;
  signal array_obj_ref_879_index_0_resize_ack_0 : boolean;
  signal switch_stmt_842_branch_1_ack_1 : boolean;
  signal ptr_deref_884_base_resize_ack_0 : boolean;
  signal array_obj_ref_879_offset_inst_req_0 : boolean;
  signal array_obj_ref_879_index_0_rename_req_0 : boolean;
  signal if_stmt_892_branch_req_0 : boolean;
  signal ptr_deref_884_gather_scatter_req_0 : boolean;
  signal if_stmt_892_branch_ack_1 : boolean;
  signal binary_911_inst_ack_0 : boolean;
  signal binary_911_inst_req_1 : boolean;
  signal binary_911_inst_ack_1 : boolean;
  signal ptr_deref_884_load_0_req_1 : boolean;
  signal ptr_deref_827_gather_scatter_req_0 : boolean;
  signal addr_of_916_final_reg_req_0 : boolean;
  signal addr_of_916_final_reg_ack_0 : boolean;
  signal if_stmt_892_branch_ack_0 : boolean;
  signal ptr_deref_827_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_915_root_address_inst_ack_0 : boolean;
  signal binary_911_inst_req_0 : boolean;
  signal array_obj_ref_879_root_address_inst_req_0 : boolean;
  signal binary_890_inst_req_0 : boolean;
  signal if_stmt_870_branch_req_0 : boolean;
  signal binary_890_inst_req_1 : boolean;
  signal binary_890_inst_ack_1 : boolean;
  signal array_obj_ref_915_offset_inst_req_0 : boolean;
  signal array_obj_ref_915_offset_inst_ack_0 : boolean;
  signal ptr_deref_923_root_address_inst_req_0 : boolean;
  signal ptr_deref_923_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_915_index_0_resize_ack_0 : boolean;
  signal ptr_deref_923_base_resize_req_0 : boolean;
  signal ptr_deref_923_base_resize_ack_0 : boolean;
  signal binary_903_inst_req_1 : boolean;
  signal binary_903_inst_ack_1 : boolean;
  signal array_obj_ref_915_index_0_resize_req_0 : boolean;
  signal binary_903_inst_req_0 : boolean;
  signal binary_903_inst_ack_0 : boolean;
  signal type_cast_920_inst_ack_0 : boolean;
  signal type_cast_920_inst_req_0 : boolean;
  signal ptr_deref_923_addr_0_req_0 : boolean;
  signal ptr_deref_923_addr_0_ack_0 : boolean;
  signal array_obj_ref_915_index_0_rename_req_0 : boolean;
  signal array_obj_ref_915_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_915_root_address_inst_req_0 : boolean;
  signal binary_868_inst_req_0 : boolean;
  signal switch_stmt_842_branch_default_ack_0 : boolean;
  signal switch_stmt_842_branch_0_req_0 : boolean;
  signal type_cast_864_inst_ack_0 : boolean;
  signal type_cast_864_inst_req_0 : boolean;
  signal addr_of_880_final_reg_ack_0 : boolean;
  signal switch_stmt_842_select_expr_0_ack_1 : boolean;
  signal addr_of_880_final_reg_req_0 : boolean;
  signal ptr_deref_923_gather_scatter_req_0 : boolean;
  signal ptr_deref_923_gather_scatter_ack_0 : boolean;
  signal ptr_deref_923_store_0_req_0 : boolean;
  signal ptr_deref_923_store_0_ack_0 : boolean;
  signal ptr_deref_923_store_0_req_1 : boolean;
  signal ptr_deref_923_store_0_ack_1 : boolean;
  signal simple_obj_ref_933_inst_req_0 : boolean;
  signal simple_obj_ref_933_inst_ack_0 : boolean;
  signal simple_obj_ref_943_inst_req_0 : boolean;
  signal simple_obj_ref_943_inst_ack_0 : boolean;
  signal simple_obj_ref_954_inst_req_0 : boolean;
  signal simple_obj_ref_954_inst_ack_0 : boolean;
  signal simple_obj_ref_967_inst_req_0 : boolean;
  signal simple_obj_ref_967_inst_ack_0 : boolean;
  signal binary_973_inst_req_0 : boolean;
  signal binary_973_inst_ack_0 : boolean;
  signal binary_973_inst_req_1 : boolean;
  signal binary_973_inst_ack_1 : boolean;
  signal if_stmt_975_branch_req_0 : boolean;
  signal if_stmt_975_branch_ack_1 : boolean;
  signal if_stmt_975_branch_ack_0 : boolean;
  signal binary_994_inst_req_0 : boolean;
  signal binary_994_inst_ack_0 : boolean;
  signal binary_994_inst_req_1 : boolean;
  signal binary_994_inst_ack_1 : boolean;
  signal binary_1000_inst_req_0 : boolean;
  signal binary_1000_inst_ack_0 : boolean;
  signal binary_1000_inst_req_1 : boolean;
  signal binary_1000_inst_ack_1 : boolean;
  signal binary_1006_inst_req_0 : boolean;
  signal binary_1006_inst_ack_0 : boolean;
  signal binary_1006_inst_req_1 : boolean;
  signal binary_1006_inst_ack_1 : boolean;
  signal binary_1011_inst_req_0 : boolean;
  signal binary_1011_inst_ack_0 : boolean;
  signal binary_1011_inst_req_1 : boolean;
  signal binary_1011_inst_ack_1 : boolean;
  signal if_stmt_1013_branch_req_0 : boolean;
  signal if_stmt_1013_branch_ack_1 : boolean;
  signal if_stmt_1013_branch_ack_0 : boolean;
  signal type_cast_1022_inst_req_0 : boolean;
  signal type_cast_1022_inst_ack_0 : boolean;
  signal binary_1026_inst_req_0 : boolean;
  signal binary_1026_inst_ack_0 : boolean;
  signal binary_1026_inst_req_1 : boolean;
  signal binary_1026_inst_ack_1 : boolean;
  signal if_stmt_1028_branch_req_0 : boolean;
  signal if_stmt_1028_branch_ack_1 : boolean;
  signal if_stmt_1028_branch_ack_0 : boolean;
  signal array_obj_ref_1045_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1045_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1045_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1045_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1045_offset_inst_req_0 : boolean;
  signal array_obj_ref_1045_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1045_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1045_root_address_inst_ack_0 : boolean;
  signal addr_of_1046_final_reg_req_0 : boolean;
  signal addr_of_1046_final_reg_ack_0 : boolean;
  signal ptr_deref_1049_base_resize_req_0 : boolean;
  signal ptr_deref_1049_base_resize_ack_0 : boolean;
  signal ptr_deref_1049_root_address_inst_req_0 : boolean;
  signal ptr_deref_1049_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1049_addr_0_req_0 : boolean;
  signal ptr_deref_1049_addr_0_ack_0 : boolean;
  signal ptr_deref_1049_gather_scatter_req_0 : boolean;
  signal ptr_deref_1049_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1049_store_0_req_0 : boolean;
  signal ptr_deref_1049_store_0_ack_0 : boolean;
  signal ptr_deref_1049_store_0_req_1 : boolean;
  signal ptr_deref_1049_store_0_ack_1 : boolean;
  signal type_cast_856_inst_req_0 : boolean;
  signal type_cast_856_inst_ack_0 : boolean;
  signal phi_stmt_853_req_0 : boolean;
  signal phi_stmt_853_req_1 : boolean;
  signal phi_stmt_853_ack_0 : boolean;
  signal phi_stmt_982_req_1 : boolean;
  signal type_cast_985_inst_req_0 : boolean;
  signal type_cast_985_inst_ack_0 : boolean;
  signal phi_stmt_982_req_0 : boolean;
  signal phi_stmt_982_ack_0 : boolean;
  signal phi_stmt_1035_req_1 : boolean;
  signal type_cast_1038_inst_req_0 : boolean;
  signal type_cast_1038_inst_ack_0 : boolean;
  signal phi_stmt_1035_req_0 : boolean;
  signal phi_stmt_1035_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  free_queue_manager_CP_3612: Block -- control-path 
    signal cp_elements: BooleanArray(255 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(43);
    cp_elements(3) <= OrReduce(cp_elements(233) & cp_elements(237));
    cp_elements(4) <= OrReduce(cp_elements(239) & cp_elements(79));
    cp_elements(5) <= OrReduce(cp_elements(241) & cp_elements(111));
    cp_elements(6) <= cp_elements(144);
    simple_obj_ref_933_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= OrReduce(cp_elements(243) & cp_elements(247));
    cp_elements(8) <= cp_elements(184);
    cp_elements(9) <= OrReduce(cp_elements(249) & cp_elements(193));
    cp_elements(10) <= OrReduce(cp_elements(251) & cp_elements(255));
    cp_elements(11) <= cp_elements(0);
    cp_elements(12) <= cp_elements(11);
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(15));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_794_gather_scatter_req_0 <= cp_elements(13);
    cp_elements(14) <= cp_elements(11);
    cp_elements(15) <= cp_elements(11);
    cp_elements(16) <= ptr_deref_794_gather_scatter_ack_0;
    ptr_deref_794_store_0_req_0 <= cp_elements(16);
    cp_elements(17) <= ptr_deref_794_store_0_ack_0;
    cp_elements(18) <= cp_elements(17);
    ptr_deref_794_store_0_req_1 <= cp_elements(18);
    cp_elements(19) <= ptr_deref_794_store_0_ack_1;
    cp_elements(20) <= cp_elements(11);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(23) & cp_elements(17) & cp_elements(20));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_805_gather_scatter_req_0 <= cp_elements(21);
    cp_elements(22) <= cp_elements(11);
    cp_elements(23) <= cp_elements(11);
    cp_elements(24) <= ptr_deref_805_gather_scatter_ack_0;
    ptr_deref_805_store_0_req_0 <= cp_elements(24);
    cp_elements(25) <= ptr_deref_805_store_0_ack_0;
    cp_elements(26) <= cp_elements(25);
    ptr_deref_805_store_0_req_1 <= cp_elements(26);
    cp_elements(27) <= ptr_deref_805_store_0_ack_1;
    cp_elements(28) <= cp_elements(11);
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(25) & cp_elements(28) & cp_elements(31));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_816_gather_scatter_req_0 <= cp_elements(29);
    cp_elements(30) <= cp_elements(11);
    cp_elements(31) <= cp_elements(11);
    cp_elements(32) <= ptr_deref_816_gather_scatter_ack_0;
    ptr_deref_816_store_0_req_0 <= cp_elements(32);
    cp_elements(33) <= ptr_deref_816_store_0_ack_0;
    cp_elements(34) <= cp_elements(33);
    ptr_deref_816_store_0_req_1 <= cp_elements(34);
    cp_elements(35) <= ptr_deref_816_store_0_ack_1;
    cp_elements(36) <= cp_elements(11);
    cpelement_group_37 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(36) & cp_elements(39) & cp_elements(33));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(37),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_827_gather_scatter_req_0 <= cp_elements(37);
    cp_elements(38) <= cp_elements(11);
    cp_elements(39) <= cp_elements(11);
    cp_elements(40) <= ptr_deref_827_gather_scatter_ack_0;
    ptr_deref_827_store_0_req_0 <= cp_elements(40);
    cp_elements(41) <= ptr_deref_827_store_0_ack_0;
    ptr_deref_827_store_0_req_1 <= cp_elements(41);
    cp_elements(42) <= ptr_deref_827_store_0_ack_1;
    cpelement_group_43 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(35) & cp_elements(14) & cp_elements(19) & cp_elements(38) & cp_elements(27) & cp_elements(42) & cp_elements(30));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(43),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(44) <= simple_obj_ref_840_inst_ack_0;
    cp_elements(45) <= cp_elements(44);
    cp_elements(46) <= false;
    cp_elements(47) <= cp_elements(46);
    cp_elements(48) <= cp_elements(44);
    cp_elements(49) <= cp_elements(48);
    cp_elements(50) <= cp_elements(49);
    switch_stmt_842_select_expr_0_req_0 <= cp_elements(50);
    cp_elements(51) <= switch_stmt_842_select_expr_0_ack_0;
    switch_stmt_842_select_expr_0_req_1 <= cp_elements(51);
    cp_elements(52) <= switch_stmt_842_select_expr_0_ack_1;
    switch_stmt_842_branch_0_req_0 <= cp_elements(52);
    cp_elements(53) <= cp_elements(49);
    switch_stmt_842_select_expr_1_req_0 <= cp_elements(53);
    cp_elements(54) <= switch_stmt_842_select_expr_1_ack_0;
    switch_stmt_842_select_expr_1_req_1 <= cp_elements(54);
    cp_elements(55) <= switch_stmt_842_select_expr_1_ack_1;
    switch_stmt_842_branch_1_req_0 <= cp_elements(55);
    cpelement_group_56 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(55) & cp_elements(52));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(56),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_842_branch_default_req_0 <= cp_elements(56);
    cp_elements(57) <= cp_elements(56);
    cp_elements(58) <= cp_elements(57);
    cp_elements(59) <= switch_stmt_842_branch_0_ack_1;
    phi_stmt_853_req_1 <= cp_elements(59);
    cp_elements(60) <= cp_elements(57);
    cp_elements(61) <= switch_stmt_842_branch_1_ack_1;
    simple_obj_ref_967_inst_req_0 <= cp_elements(61);
    cp_elements(62) <= cp_elements(57);
    cp_elements(63) <= switch_stmt_842_branch_default_ack_0;
    cp_elements(64) <= cp_elements(3);
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(66));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_868_inst_req_0 <= cp_elements(65);
    cp_elements(66) <= cp_elements(64);
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(69));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_864_inst_req_0 <= cp_elements(67);
    cp_elements(68) <= cp_elements(64);
    cp_elements(69) <= cp_elements(64);
    cp_elements(70) <= type_cast_864_inst_ack_0;
    cp_elements(71) <= binary_868_inst_ack_0;
    binary_868_inst_req_1 <= cp_elements(71);
    cp_elements(72) <= binary_868_inst_ack_1;
    cp_elements(73) <= cp_elements(72);
    cp_elements(74) <= false;
    cp_elements(75) <= cp_elements(74);
    cp_elements(76) <= cp_elements(72);
    if_stmt_870_branch_req_0 <= cp_elements(76);
    cp_elements(77) <= cp_elements(76);
    cp_elements(78) <= cp_elements(77);
    cp_elements(79) <= if_stmt_870_branch_ack_1;
    cp_elements(80) <= cp_elements(77);
    cp_elements(81) <= if_stmt_870_branch_ack_0;
    simple_obj_ref_954_inst_req_0 <= cp_elements(81);
    cp_elements(82) <= cp_elements(4);
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(84));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_880_final_reg_req_0 <= cp_elements(83);
    cp_elements(84) <= cp_elements(82);
    cp_elements(85) <= cp_elements(82);
    array_obj_ref_879_index_0_resize_req_0 <= cp_elements(85);
    cp_elements(86) <= array_obj_ref_879_index_0_resize_ack_0;
    array_obj_ref_879_index_0_rename_req_0 <= cp_elements(86);
    cp_elements(87) <= array_obj_ref_879_index_0_rename_ack_0;
    array_obj_ref_879_offset_inst_req_0 <= cp_elements(87);
    cp_elements(88) <= array_obj_ref_879_offset_inst_ack_0;
    array_obj_ref_879_root_address_inst_req_0 <= cp_elements(88);
    cp_elements(89) <= array_obj_ref_879_root_address_inst_ack_0;
    cp_elements(90) <= addr_of_880_final_reg_ack_0;
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_884_load_0_req_0 <= cp_elements(91);
    cp_elements(92) <= cp_elements(90);
    ptr_deref_884_base_resize_req_0 <= cp_elements(92);
    cp_elements(93) <= ptr_deref_884_base_resize_ack_0;
    ptr_deref_884_root_address_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= ptr_deref_884_root_address_inst_ack_0;
    ptr_deref_884_addr_0_req_0 <= cp_elements(94);
    cp_elements(95) <= ptr_deref_884_addr_0_ack_0;
    cp_elements(96) <= ptr_deref_884_load_0_ack_0;
    ptr_deref_884_load_0_req_1 <= cp_elements(96);
    cp_elements(97) <= ptr_deref_884_load_0_ack_1;
    ptr_deref_884_gather_scatter_req_0 <= cp_elements(97);
    cp_elements(98) <= ptr_deref_884_gather_scatter_ack_0;
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(98) & cp_elements(100));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_890_inst_req_0 <= cp_elements(99);
    cp_elements(100) <= cp_elements(82);
    cp_elements(101) <= binary_890_inst_ack_0;
    binary_890_inst_req_1 <= cp_elements(101);
    cp_elements(102) <= binary_890_inst_ack_1;
    cp_elements(103) <= cp_elements(102);
    cp_elements(104) <= false;
    cp_elements(105) <= cp_elements(104);
    cp_elements(106) <= cp_elements(102);
    if_stmt_892_branch_req_0 <= cp_elements(106);
    cp_elements(107) <= cp_elements(106);
    cp_elements(108) <= cp_elements(107);
    cp_elements(109) <= if_stmt_892_branch_ack_1;
    cp_elements(110) <= cp_elements(107);
    cp_elements(111) <= if_stmt_892_branch_ack_0;
    cp_elements(112) <= cp_elements(5);
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(115));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_903_inst_req_0 <= cp_elements(113);
    cp_elements(114) <= cp_elements(112);
    cp_elements(115) <= cp_elements(112);
    cp_elements(116) <= binary_903_inst_ack_0;
    binary_903_inst_req_1 <= cp_elements(116);
    cp_elements(117) <= binary_903_inst_ack_1;
    type_cast_856_inst_req_0 <= cp_elements(117);
    cp_elements(118) <= cp_elements(109);
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(121) & cp_elements(120));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_911_inst_req_0 <= cp_elements(119);
    cp_elements(120) <= cp_elements(118);
    cp_elements(121) <= cp_elements(118);
    cp_elements(122) <= binary_911_inst_ack_0;
    binary_911_inst_req_1 <= cp_elements(122);
    cp_elements(123) <= binary_911_inst_ack_1;
    array_obj_ref_915_index_0_resize_req_0 <= cp_elements(123);
    cpelement_group_124 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(129));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_916_final_reg_req_0 <= cp_elements(124);
    cp_elements(125) <= cp_elements(118);
    cp_elements(126) <= array_obj_ref_915_index_0_resize_ack_0;
    array_obj_ref_915_index_0_rename_req_0 <= cp_elements(126);
    cp_elements(127) <= array_obj_ref_915_index_0_rename_ack_0;
    array_obj_ref_915_offset_inst_req_0 <= cp_elements(127);
    cp_elements(128) <= array_obj_ref_915_offset_inst_ack_0;
    array_obj_ref_915_root_address_inst_req_0 <= cp_elements(128);
    cp_elements(129) <= array_obj_ref_915_root_address_inst_ack_0;
    cp_elements(130) <= addr_of_916_final_reg_ack_0;
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(130));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_920_inst_req_0 <= cp_elements(131);
    cp_elements(132) <= cp_elements(118);
    cp_elements(133) <= type_cast_920_inst_ack_0;
    cp_elements(134) <= cp_elements(118);
    cpelement_group_135 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(140) & cp_elements(136) & cp_elements(134));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(135),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_923_gather_scatter_req_0 <= cp_elements(135);
    cp_elements(136) <= cp_elements(118);
    cp_elements(137) <= cp_elements(136);
    ptr_deref_923_base_resize_req_0 <= cp_elements(137);
    cp_elements(138) <= ptr_deref_923_base_resize_ack_0;
    ptr_deref_923_root_address_inst_req_0 <= cp_elements(138);
    cp_elements(139) <= ptr_deref_923_root_address_inst_ack_0;
    ptr_deref_923_addr_0_req_0 <= cp_elements(139);
    cp_elements(140) <= ptr_deref_923_addr_0_ack_0;
    cp_elements(141) <= ptr_deref_923_gather_scatter_ack_0;
    ptr_deref_923_store_0_req_0 <= cp_elements(141);
    cp_elements(142) <= ptr_deref_923_store_0_ack_0;
    ptr_deref_923_store_0_req_1 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_923_store_0_ack_1;
    cpelement_group_144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(133));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(145) <= simple_obj_ref_933_inst_ack_0;
    simple_obj_ref_943_inst_req_0 <= cp_elements(145);
    cp_elements(146) <= simple_obj_ref_943_inst_ack_0;
    cp_elements(147) <= simple_obj_ref_954_inst_ack_0;
    cp_elements(148) <= simple_obj_ref_967_inst_ack_0;
    cp_elements(149) <= cp_elements(148);
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(151) & cp_elements(152));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_973_inst_req_0 <= cp_elements(150);
    cp_elements(151) <= cp_elements(149);
    cp_elements(152) <= cp_elements(149);
    cp_elements(153) <= binary_973_inst_ack_0;
    binary_973_inst_req_1 <= cp_elements(153);
    cp_elements(154) <= binary_973_inst_ack_1;
    cp_elements(155) <= cp_elements(154);
    cp_elements(156) <= false;
    cp_elements(157) <= cp_elements(156);
    cp_elements(158) <= cp_elements(154);
    if_stmt_975_branch_req_0 <= cp_elements(158);
    cp_elements(159) <= cp_elements(158);
    cp_elements(160) <= cp_elements(159);
    cp_elements(161) <= if_stmt_975_branch_ack_1;
    phi_stmt_982_req_1 <= cp_elements(161);
    cp_elements(162) <= cp_elements(159);
    cp_elements(163) <= if_stmt_975_branch_ack_0;
    phi_stmt_1035_req_1 <= cp_elements(163);
    cp_elements(164) <= cp_elements(7);
    cpelement_group_165 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(166) & cp_elements(167));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(165),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_994_inst_req_0 <= cp_elements(165);
    cp_elements(166) <= cp_elements(164);
    cp_elements(167) <= cp_elements(164);
    cp_elements(168) <= binary_994_inst_ack_0;
    binary_994_inst_req_1 <= cp_elements(168);
    cp_elements(169) <= binary_994_inst_ack_1;
    cpelement_group_170 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(172));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(170),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1000_inst_req_0 <= cp_elements(170);
    cp_elements(171) <= cp_elements(164);
    cp_elements(172) <= cp_elements(164);
    cp_elements(173) <= binary_1000_inst_ack_0;
    binary_1000_inst_req_1 <= cp_elements(173);
    cp_elements(174) <= binary_1000_inst_ack_1;
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(176));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1006_inst_req_0 <= cp_elements(175);
    cp_elements(176) <= cp_elements(164);
    cp_elements(177) <= binary_1006_inst_ack_0;
    binary_1006_inst_req_1 <= cp_elements(177);
    cp_elements(178) <= binary_1006_inst_ack_1;
    cpelement_group_179 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(180) & cp_elements(181));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(179),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1011_inst_req_0 <= cp_elements(179);
    cp_elements(180) <= cp_elements(164);
    cp_elements(181) <= cp_elements(164);
    cp_elements(182) <= binary_1011_inst_ack_0;
    binary_1011_inst_req_1 <= cp_elements(182);
    cp_elements(183) <= binary_1011_inst_ack_1;
    cpelement_group_184 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(174) & cp_elements(183));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(185) <= cp_elements(8);
    cp_elements(186) <= false;
    cp_elements(187) <= cp_elements(186);
    cp_elements(188) <= cp_elements(8);
    if_stmt_1013_branch_req_0 <= cp_elements(188);
    cp_elements(189) <= cp_elements(188);
    cp_elements(190) <= cp_elements(189);
    cp_elements(191) <= if_stmt_1013_branch_ack_1;
    type_cast_985_inst_req_0 <= cp_elements(191);
    cp_elements(192) <= cp_elements(189);
    cp_elements(193) <= if_stmt_1013_branch_ack_0;
    cp_elements(194) <= cp_elements(9);
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(196));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1026_inst_req_0 <= cp_elements(195);
    cp_elements(196) <= cp_elements(194);
    cpelement_group_197 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(198) & cp_elements(199));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(197),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1022_inst_req_0 <= cp_elements(197);
    cp_elements(198) <= cp_elements(194);
    cp_elements(199) <= cp_elements(194);
    cp_elements(200) <= type_cast_1022_inst_ack_0;
    cp_elements(201) <= binary_1026_inst_ack_0;
    binary_1026_inst_req_1 <= cp_elements(201);
    cp_elements(202) <= binary_1026_inst_ack_1;
    cp_elements(203) <= cp_elements(202);
    cp_elements(204) <= false;
    cp_elements(205) <= cp_elements(204);
    cp_elements(206) <= cp_elements(202);
    if_stmt_1028_branch_req_0 <= cp_elements(206);
    cp_elements(207) <= cp_elements(206);
    cp_elements(208) <= cp_elements(207);
    cp_elements(209) <= if_stmt_1028_branch_ack_1;
    type_cast_1038_inst_req_0 <= cp_elements(209);
    cp_elements(210) <= cp_elements(207);
    cp_elements(211) <= if_stmt_1028_branch_ack_0;
    cp_elements(212) <= cp_elements(10);
    cpelement_group_213 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(214) & cp_elements(219));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(213),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    addr_of_1046_final_reg_req_0 <= cp_elements(213);
    cp_elements(214) <= cp_elements(212);
    cp_elements(215) <= cp_elements(212);
    array_obj_ref_1045_index_0_resize_req_0 <= cp_elements(215);
    cp_elements(216) <= array_obj_ref_1045_index_0_resize_ack_0;
    array_obj_ref_1045_index_0_rename_req_0 <= cp_elements(216);
    cp_elements(217) <= array_obj_ref_1045_index_0_rename_ack_0;
    array_obj_ref_1045_offset_inst_req_0 <= cp_elements(217);
    cp_elements(218) <= array_obj_ref_1045_offset_inst_ack_0;
    array_obj_ref_1045_root_address_inst_req_0 <= cp_elements(218);
    cp_elements(219) <= array_obj_ref_1045_root_address_inst_ack_0;
    cp_elements(220) <= addr_of_1046_final_reg_ack_0;
    cp_elements(221) <= cp_elements(212);
    cpelement_group_222 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(220) & cp_elements(221) & cp_elements(226));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(222),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1049_gather_scatter_req_0 <= cp_elements(222);
    cp_elements(223) <= cp_elements(220);
    ptr_deref_1049_base_resize_req_0 <= cp_elements(223);
    cp_elements(224) <= ptr_deref_1049_base_resize_ack_0;
    ptr_deref_1049_root_address_inst_req_0 <= cp_elements(224);
    cp_elements(225) <= ptr_deref_1049_root_address_inst_ack_0;
    ptr_deref_1049_addr_0_req_0 <= cp_elements(225);
    cp_elements(226) <= ptr_deref_1049_addr_0_ack_0;
    cp_elements(227) <= ptr_deref_1049_gather_scatter_ack_0;
    ptr_deref_1049_store_0_req_0 <= cp_elements(227);
    cp_elements(228) <= ptr_deref_1049_store_0_ack_0;
    ptr_deref_1049_store_0_req_1 <= cp_elements(228);
    cp_elements(229) <= ptr_deref_1049_store_0_ack_1;
    cp_elements(230) <= OrReduce(cp_elements(211) & cp_elements(229) & cp_elements(2) & cp_elements(63) & cp_elements(146) & cp_elements(147));
    cp_elements(231) <= cp_elements(230);
    simple_obj_ref_840_inst_req_0 <= cp_elements(231);
    cp_elements(232) <= false;
    cp_elements(233) <= cp_elements(232);
    cp_elements(234) <= type_cast_856_inst_ack_0;
    phi_stmt_853_req_0 <= cp_elements(234);
    cp_elements(235) <= OrReduce(cp_elements(234) & cp_elements(59));
    cp_elements(236) <= cp_elements(235);
    cp_elements(237) <= phi_stmt_853_ack_0;
    cp_elements(238) <= false;
    cp_elements(239) <= cp_elements(238);
    cp_elements(240) <= false;
    cp_elements(241) <= cp_elements(240);
    cp_elements(242) <= false;
    cp_elements(243) <= cp_elements(242);
    cp_elements(244) <= type_cast_985_inst_ack_0;
    phi_stmt_982_req_0 <= cp_elements(244);
    cp_elements(245) <= OrReduce(cp_elements(161) & cp_elements(244));
    cp_elements(246) <= cp_elements(245);
    cp_elements(247) <= phi_stmt_982_ack_0;
    cp_elements(248) <= false;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= false;
    cp_elements(251) <= cp_elements(250);
    cp_elements(252) <= type_cast_1038_inst_ack_0;
    phi_stmt_1035_req_0 <= cp_elements(252);
    cp_elements(253) <= OrReduce(cp_elements(163) & cp_elements(252));
    cp_elements(254) <= cp_elements(253);
    cp_elements(255) <= phi_stmt_1035_ack_0;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1045_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_1045_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_1045_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_1045_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_879_final_offset : std_logic_vector(2 downto 0);
    signal array_obj_ref_879_offset_scale_factor_0 : std_logic_vector(2 downto 0);
    signal array_obj_ref_879_resized_base_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_879_root_address : std_logic_vector(2 downto 0);
    signal array_obj_ref_915_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_915_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_915_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_915_root_address : std_logic_vector(10 downto 0);
    signal expr_844_wire_constant : std_logic_vector(7 downto 0);
    signal expr_844_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_847_wire_constant : std_logic_vector(7 downto 0);
    signal expr_847_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal i3x_x044_982 : std_logic_vector(31 downto 0);
    signal i3x_x0x_xlcssa53_1035 : std_logic_vector(31 downto 0);
    signal iNsTr_0_792 : std_logic_vector(31 downto 0);
    signal iNsTr_11_853 : std_logic_vector(31 downto 0);
    signal iNsTr_13_965 : std_logic_vector(31 downto 0);
    signal iNsTr_16_953 : std_logic_vector(31 downto 0);
    signal iNsTr_19_1001 : std_logic_vector(31 downto 0);
    signal iNsTr_24_932 : std_logic_vector(31 downto 0);
    signal iNsTr_26_942 : std_logic_vector(31 downto 0);
    signal iNsTr_2_803 : std_logic_vector(31 downto 0);
    signal iNsTr_4_814 : std_logic_vector(31 downto 0);
    signal iNsTr_6_825 : std_logic_vector(31 downto 0);
    signal iNsTr_9_838 : std_logic_vector(31 downto 0);
    signal ptr_deref_1049_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1049_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1049_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_1049_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1049_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_1049_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_794_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_794_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_794_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_805_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_805_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_805_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_816_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_816_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_816_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_827_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_827_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_827_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_884_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_884_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_884_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_884_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_884_word_offset_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_923_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_923_resized_base_address : std_logic_vector(2 downto 0);
    signal ptr_deref_923_root_address : std_logic_vector(2 downto 0);
    signal ptr_deref_923_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_923_word_address_0 : std_logic_vector(2 downto 0);
    signal ptr_deref_923_word_offset_0 : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1044_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_1044_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_878_resized : std_logic_vector(2 downto 0);
    signal simple_obj_ref_878_scaled : std_logic_vector(2 downto 0);
    signal simple_obj_ref_914_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_914_scaled : std_logic_vector(10 downto 0);
    signal tmp10_869 : std_logic_vector(0 downto 0);
    signal tmp12_881 : std_logic_vector(31 downto 0);
    signal tmp13_885 : std_logic_vector(7 downto 0);
    signal tmp14_891 : std_logic_vector(0 downto 0);
    signal tmp16_912 : std_logic_vector(31 downto 0);
    signal tmp17_917 : std_logic_vector(31 downto 0);
    signal tmp18_921 : std_logic_vector(31 downto 0);
    signal tmp21_904 : std_logic_vector(31 downto 0);
    signal tmp28_968 : std_logic_vector(31 downto 0);
    signal tmp31_1007 : std_logic_vector(31 downto 0);
    signal tmp3243_974 : std_logic_vector(0 downto 0);
    signal tmp32_1012 : std_logic_vector(0 downto 0);
    signal tmp36_1027 : std_logic_vector(0 downto 0);
    signal tmp38_1047 : std_logic_vector(31 downto 0);
    signal tmp50_995 : std_logic_vector(31 downto 0);
    signal tmp6_841 : std_logic_vector(7 downto 0);
    signal type_cast_1005_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1022_wire : std_logic_vector(31 downto 0);
    signal type_cast_1025_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1038_wire : std_logic_vector(31 downto 0);
    signal type_cast_1041_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1051_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_796_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_807_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_818_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_829_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_856_wire : std_logic_vector(31 downto 0);
    signal type_cast_859_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_864_wire : std_logic_vector(31 downto 0);
    signal type_cast_867_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_889_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_902_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_910_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_925_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_935_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_956_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_972_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_985_wire : std_logic_vector(31 downto 0);
    signal type_cast_988_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_993_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_999_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1045_offset_scale_factor_0 <= "001";
    array_obj_ref_1045_resized_base_address <= "000";
    array_obj_ref_879_offset_scale_factor_0 <= "001";
    array_obj_ref_879_resized_base_address <= "000";
    array_obj_ref_915_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_915_resized_base_address <= "00000000000";
    expr_844_wire_constant <= "00000010";
    expr_847_wire_constant <= "00000001";
    iNsTr_0_792 <= "00000000000000000000000000000000";
    iNsTr_13_965 <= "00000000000000000000000000000000";
    iNsTr_16_953 <= "00000000000000000000000000000000";
    iNsTr_24_932 <= "00000000000000000000000000000000";
    iNsTr_26_942 <= "00000000000000000000000000000000";
    iNsTr_2_803 <= "00000000000000000000000000000001";
    iNsTr_4_814 <= "00000000000000000000000000000010";
    iNsTr_6_825 <= "00000000000000000000000000000011";
    iNsTr_9_838 <= "00000000000000000000000000000000";
    ptr_deref_1049_word_offset_0 <= "000";
    ptr_deref_794_word_address_0 <= "000";
    ptr_deref_805_word_address_0 <= "001";
    ptr_deref_816_word_address_0 <= "010";
    ptr_deref_827_word_address_0 <= "011";
    ptr_deref_884_word_offset_0 <= "000";
    ptr_deref_923_word_offset_0 <= "000";
    type_cast_1005_wire_constant <= "00000000000000000000001000000000";
    type_cast_1025_wire_constant <= "00000000000000000000000000000100";
    type_cast_1041_wire_constant <= "00000000000000000000000000000000";
    type_cast_1051_wire_constant <= "00000001";
    type_cast_796_wire_constant <= "00000001";
    type_cast_807_wire_constant <= "00000001";
    type_cast_818_wire_constant <= "00000001";
    type_cast_829_wire_constant <= "00000001";
    type_cast_859_wire_constant <= "00000000000000000000000000000000";
    type_cast_867_wire_constant <= "00000000000000000000000000000100";
    type_cast_889_wire_constant <= "00000001";
    type_cast_902_wire_constant <= "00000000000000000000000000000001";
    type_cast_910_wire_constant <= "00000000000000000000000000001000";
    type_cast_925_wire_constant <= "00000000";
    type_cast_935_wire_constant <= "00000011";
    type_cast_956_wire_constant <= "00000100";
    type_cast_972_wire_constant <= "00000000000000000000000100000000";
    type_cast_988_wire_constant <= "00000000000000000000000000000000";
    type_cast_993_wire_constant <= "00000000000000000000000000001000";
    type_cast_999_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1035: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1038_wire & type_cast_1041_wire_constant;
      req <= phi_stmt_1035_req_0 & phi_stmt_1035_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1035_ack_0,
          idata => idata,
          odata => i3x_x0x_xlcssa53_1035,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1035
    phi_stmt_853: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_856_wire & type_cast_859_wire_constant;
      req <= phi_stmt_853_req_0 & phi_stmt_853_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_853_ack_0,
          idata => idata,
          odata => iNsTr_11_853,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_853
    phi_stmt_982: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_985_wire & type_cast_988_wire_constant;
      req <= phi_stmt_982_req_0 & phi_stmt_982_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_982_ack_0,
          idata => idata,
          odata => i3x_x044_982,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_982
    addr_of_1046_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1045_root_address, dout => tmp38_1047, req => addr_of_1046_final_reg_req_0, ack => addr_of_1046_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_880_final_reg: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_879_root_address, dout => tmp12_881, req => addr_of_880_final_reg_req_0, ack => addr_of_880_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_916_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_915_root_address, dout => tmp17_917, req => addr_of_916_final_reg_req_0, ack => addr_of_916_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1045_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => i3x_x0x_xlcssa53_1035, dout => simple_obj_ref_1044_resized, req => array_obj_ref_1045_index_0_resize_req_0, ack => array_obj_ref_1045_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1045_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_1044_scaled, dout => array_obj_ref_1045_final_offset, req => array_obj_ref_1045_offset_inst_req_0, ack => array_obj_ref_1045_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_879_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => iNsTr_11_853, dout => simple_obj_ref_878_resized, req => array_obj_ref_879_index_0_resize_req_0, ack => array_obj_ref_879_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_879_offset_inst: RegisterBase --
      generic map(in_data_width => 3,out_data_width => 3, flow_through => true ) 
      port map( din => simple_obj_ref_878_scaled, dout => array_obj_ref_879_final_offset, req => array_obj_ref_879_offset_inst_req_0, ack => array_obj_ref_879_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_915_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp16_912, dout => simple_obj_ref_914_resized, req => array_obj_ref_915_index_0_resize_req_0, ack => array_obj_ref_915_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_915_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_914_scaled, dout => array_obj_ref_915_final_offset, req => array_obj_ref_915_offset_inst_req_0, ack => array_obj_ref_915_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1049_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp38_1047, dout => ptr_deref_1049_resized_base_address, req => ptr_deref_1049_base_resize_req_0, ack => ptr_deref_1049_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_884_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_881, dout => ptr_deref_884_resized_base_address, req => ptr_deref_884_base_resize_req_0, ack => ptr_deref_884_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_923_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 3, flow_through => true ) 
      port map( din => tmp12_881, dout => ptr_deref_923_resized_base_address, req => ptr_deref_923_base_resize_req_0, ack => ptr_deref_923_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1022_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_19_1001, dout => type_cast_1022_wire, req => type_cast_1022_inst_req_0, ack => type_cast_1022_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1038_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_19_1001, dout => type_cast_1038_wire, req => type_cast_1038_inst_req_0, ack => type_cast_1038_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_856_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp21_904, dout => type_cast_856_wire, req => type_cast_856_inst_req_0, ack => type_cast_856_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_864_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_11_853, dout => type_cast_864_wire, req => type_cast_864_inst_req_0, ack => type_cast_864_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_920_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_917, dout => tmp18_921, req => type_cast_920_inst_req_0, ack => type_cast_920_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_985_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_19_1001, dout => type_cast_985_wire, req => type_cast_985_inst_req_0, ack => type_cast_985_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1045_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1045_index_0_rename_ack_0 <= array_obj_ref_1045_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1044_resized;
      simple_obj_ref_1044_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_1045_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_1045_root_address_inst_ack_0 <= array_obj_ref_1045_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1045_final_offset;
      array_obj_ref_1045_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_879_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_879_index_0_rename_ack_0 <= array_obj_ref_879_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_878_resized;
      simple_obj_ref_878_scaled <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_879_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      array_obj_ref_879_root_address_inst_ack_0 <= array_obj_ref_879_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_879_final_offset;
      array_obj_ref_879_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    array_obj_ref_915_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_915_index_0_rename_ack_0 <= array_obj_ref_915_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_914_resized;
      simple_obj_ref_914_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_915_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_915_root_address_inst_ack_0 <= array_obj_ref_915_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_915_final_offset;
      array_obj_ref_915_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1049_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1049_addr_0_ack_0 <= ptr_deref_1049_addr_0_req_0;
      aggregated_sig <= ptr_deref_1049_root_address;
      ptr_deref_1049_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_1049_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1049_gather_scatter_ack_0 <= ptr_deref_1049_gather_scatter_req_0;
      aggregated_sig <= type_cast_1051_wire_constant;
      ptr_deref_1049_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1049_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_1049_root_address_inst_ack_0 <= ptr_deref_1049_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1049_resized_base_address;
      ptr_deref_1049_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_794_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_794_gather_scatter_ack_0 <= ptr_deref_794_gather_scatter_req_0;
      aggregated_sig <= type_cast_796_wire_constant;
      ptr_deref_794_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_805_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_805_gather_scatter_ack_0 <= ptr_deref_805_gather_scatter_req_0;
      aggregated_sig <= type_cast_807_wire_constant;
      ptr_deref_805_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_816_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_816_gather_scatter_ack_0 <= ptr_deref_816_gather_scatter_req_0;
      aggregated_sig <= type_cast_818_wire_constant;
      ptr_deref_816_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_827_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_827_gather_scatter_ack_0 <= ptr_deref_827_gather_scatter_req_0;
      aggregated_sig <= type_cast_829_wire_constant;
      ptr_deref_827_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_884_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_884_addr_0_ack_0 <= ptr_deref_884_addr_0_req_0;
      aggregated_sig <= ptr_deref_884_root_address;
      ptr_deref_884_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_884_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_884_gather_scatter_ack_0 <= ptr_deref_884_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_884_data_0;
      tmp13_885 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_884_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_884_root_address_inst_ack_0 <= ptr_deref_884_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_884_resized_base_address;
      ptr_deref_884_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_923_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_923_addr_0_ack_0 <= ptr_deref_923_addr_0_req_0;
      aggregated_sig <= ptr_deref_923_root_address;
      ptr_deref_923_word_address_0 <= aggregated_sig(2 downto 0);
      --
    end Block;
    ptr_deref_923_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_923_gather_scatter_ack_0 <= ptr_deref_923_gather_scatter_req_0;
      aggregated_sig <= type_cast_925_wire_constant;
      ptr_deref_923_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_923_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(2 downto 0); --
    begin -- 
      ptr_deref_923_root_address_inst_ack_0 <= ptr_deref_923_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_923_resized_base_address;
      ptr_deref_923_root_address <= aggregated_sig(2 downto 0);
      --
    end Block;
    if_stmt_1013_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp32_1012;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1013_branch_req_0,
          ack0 => if_stmt_1013_branch_ack_0,
          ack1 => if_stmt_1013_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1028_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_1027;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1028_branch_req_0,
          ack0 => if_stmt_1028_branch_ack_0,
          ack1 => if_stmt_1028_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_870_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp10_869;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_870_branch_req_0,
          ack0 => if_stmt_870_branch_ack_0,
          ack1 => if_stmt_870_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_892_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp14_891;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_892_branch_req_0,
          ack0 => if_stmt_892_branch_ack_0,
          ack1 => if_stmt_892_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_975_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp3243_974;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_975_branch_req_0,
          ack0 => if_stmt_975_branch_ack_0,
          ack1 => if_stmt_975_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_842_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_844_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_842_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_842_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_842_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_847_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_842_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_842_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_842_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_844_wire_constant_cmp & expr_847_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_842_branch_default_req_0,
          ack0 => switch_stmt_842_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1000_inst binary_903_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= i3x_x044_982 & iNsTr_11_853;
      iNsTr_19_1001 <= data_out(63 downto 32);
      tmp21_904 <= data_out(31 downto 0);
      reqL(1) <= binary_1000_inst_req_0;
      reqL(0) <= binary_903_inst_req_0;
      binary_1000_inst_ack_0 <= ackL(1);
      binary_903_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1000_inst_req_1;
      reqR(0) <= binary_903_inst_req_1;
      binary_1000_inst_ack_1 <= ackR(1);
      binary_903_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1006_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_995;
      tmp31_1007 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000001000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1006_inst_req_0,
          ackL => binary_1006_inst_ack_0,
          reqR => binary_1006_inst_req_1,
          ackR => binary_1006_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1011_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_968 & tmp31_1007;
      tmp32_1012 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1011_inst_req_0,
          ackL => binary_1011_inst_ack_0,
          reqR => binary_1011_inst_req_1,
          ackR => binary_1011_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1026_inst binary_868_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1022_wire & type_cast_864_wire;
      tmp36_1027 <= data_out(1 downto 1);
      tmp10_869 <= data_out(0 downto 0);
      reqL(1) <= binary_1026_inst_req_0;
      reqL(0) <= binary_868_inst_req_0;
      binary_1026_inst_ack_0 <= ackL(1);
      binary_868_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1026_inst_req_1;
      reqR(0) <= binary_868_inst_req_1;
      binary_1026_inst_ack_1 <= ackR(1);
      binary_868_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : switch_stmt_842_select_expr_1 binary_890_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_841 & tmp13_885;
      expr_847_wire_constant_cmp <= data_out(1 downto 1);
      tmp14_891 <= data_out(0 downto 0);
      reqL(1) <= switch_stmt_842_select_expr_1_req_0;
      reqL(0) <= binary_890_inst_req_0;
      switch_stmt_842_select_expr_1_ack_0 <= ackL(1);
      binary_890_inst_ack_0 <= ackL(0);
      reqR(1) <= switch_stmt_842_select_expr_1_req_1;
      reqR(0) <= binary_890_inst_req_1;
      switch_stmt_842_select_expr_1_ack_1 <= ackR(1);
      binary_890_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_911_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_11_853;
      tmp16_912 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_911_inst_req_0,
          ackL => binary_911_inst_ack_0,
          reqR => binary_911_inst_req_1,
          ackR => binary_911_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_973_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp28_968;
      tmp3243_974 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000100000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_973_inst_req_0,
          ackL => binary_973_inst_ack_0,
          reqR => binary_973_inst_req_1,
          ackR => binary_973_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_994_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i3x_x044_982;
      tmp50_995 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_994_inst_req_0,
          ackL => binary_994_inst_ack_0,
          reqR => binary_994_inst_req_1,
          ackR => binary_994_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : switch_stmt_842_select_expr_0 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_841;
      expr_844_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_842_select_expr_0_req_0,
          ackL => switch_stmt_842_select_expr_0_ack_0,
          reqR => switch_stmt_842_select_expr_0_req_1,
          ackR => switch_stmt_842_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared load operator group (0) : ptr_deref_884_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_884_load_0_req_0;
      ptr_deref_884_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_884_load_0_req_1;
      ptr_deref_884_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_884_word_address_0;
      ptr_deref_884_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 3,  num_reqs => 1,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(2 downto 0),
          mtag => memory_space_2_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 1,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(7 downto 0),
          mtag => memory_space_2_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : ptr_deref_794_store_0 ptr_deref_923_store_0 ptr_deref_1049_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(8 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_794_store_0_req_0;
      reqL(1) <= ptr_deref_923_store_0_req_0;
      reqL(0) <= ptr_deref_1049_store_0_req_0;
      ptr_deref_794_store_0_ack_0 <= ackL(2);
      ptr_deref_923_store_0_ack_0 <= ackL(1);
      ptr_deref_1049_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_794_store_0_req_1;
      reqR(1) <= ptr_deref_923_store_0_req_1;
      reqR(0) <= ptr_deref_1049_store_0_req_1;
      ptr_deref_794_store_0_ack_1 <= ackR(2);
      ptr_deref_923_store_0_ack_1 <= ackR(1);
      ptr_deref_1049_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_794_word_address_0 & ptr_deref_923_word_address_0 & ptr_deref_1049_word_address_0;
      data_in <= ptr_deref_794_data_0 & ptr_deref_923_data_0 & ptr_deref_1049_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(3),
          mack => memory_space_2_sr_ack(3),
          maddr => memory_space_2_sr_addr(11 downto 9),
          mdata => memory_space_2_sr_data(31 downto 24),
          mtag => memory_space_2_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(3),
          mack => memory_space_2_sc_ack(3),
          mtag => memory_space_2_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_805_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_805_store_0_req_0;
      ptr_deref_805_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_805_store_0_req_1;
      ptr_deref_805_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_805_word_address_0;
      data_in <= ptr_deref_805_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(2),
          mack => memory_space_2_sr_ack(2),
          maddr => memory_space_2_sr_addr(8 downto 6),
          mdata => memory_space_2_sr_data(23 downto 16),
          mtag => memory_space_2_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(2),
          mack => memory_space_2_sc_ack(2),
          mtag => memory_space_2_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_816_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_816_store_0_req_0;
      ptr_deref_816_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_816_store_0_req_1;
      ptr_deref_816_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_816_word_address_0;
      data_in <= ptr_deref_816_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(1),
          mack => memory_space_2_sr_ack(1),
          maddr => memory_space_2_sr_addr(5 downto 3),
          mdata => memory_space_2_sr_data(15 downto 8),
          mtag => memory_space_2_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(1),
          mack => memory_space_2_sc_ack(1),
          mtag => memory_space_2_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_827_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(2 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_827_store_0_req_0;
      ptr_deref_827_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_827_store_0_req_1;
      ptr_deref_827_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_827_word_address_0;
      data_in <= ptr_deref_827_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 3,
        data_width => 8,
        num_reqs => 1,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(2 downto 0),
          mdata => memory_space_2_sr_data(7 downto 0),
          mtag => memory_space_2_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared inport operator group (0) : simple_obj_ref_840_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_840_inst_req_0;
      simple_obj_ref_840_inst_ack_0 <= ack(0);
      tmp6_841 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_request_pipe_read_req(0),
          oack => free_queue_request_pipe_read_ack(0),
          odata => free_queue_request_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_967_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_967_inst_req_0;
      simple_obj_ref_967_inst_ack_0 <= ack(0);
      tmp28_968 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_put_pipe_read_req(0),
          oack => free_queue_put_pipe_read_ack(0),
          odata => free_queue_put_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_933_inst simple_obj_ref_954_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_933_inst_req_0;
      req(0) <= simple_obj_ref_954_inst_req_0;
      simple_obj_ref_933_inst_ack_0 <= ack(1);
      simple_obj_ref_954_inst_ack_0 <= ack(0);
      data_in <= type_cast_935_wire_constant & type_cast_956_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 2,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_ack_pipe_write_req(0),
          oack => free_queue_ack_pipe_write_ack(0),
          odata => free_queue_ack_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_943_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_943_inst_req_0;
      simple_obj_ref_943_inst_ack_0 <= ack(0);
      data_in <= tmp18_921;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_get_pipe_write_req(0),
          oack => free_queue_get_pipe_write_ack(0),
          odata => free_queue_get_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity output_port_lookup is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    op_lut_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    op_lut_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    op_lut_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    op_lut_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity output_port_lookup;
architecture Default of output_port_lookup is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal output_port_lookup_CP_5084_start: Boolean;
  -- links between control-path and data-path
  signal binary_1102_inst_ack_1 : boolean;
  signal simple_obj_ref_1087_inst_ack_0 : boolean;
  signal binary_1115_inst_req_1 : boolean;
  signal binary_1115_inst_req_0 : boolean;
  signal if_stmt_1104_branch_ack_1 : boolean;
  signal simple_obj_ref_1096_inst_req_0 : boolean;
  signal binary_1102_inst_ack_0 : boolean;
  signal simple_obj_ref_1096_inst_ack_0 : boolean;
  signal if_stmt_1104_branch_ack_0 : boolean;
  signal binary_1115_inst_ack_1 : boolean;
  signal binary_1115_inst_ack_0 : boolean;
  signal if_stmt_1104_branch_req_0 : boolean;
  signal binary_1102_inst_req_1 : boolean;
  signal binary_1102_inst_req_0 : boolean;
  signal simple_obj_ref_1087_inst_req_0 : boolean;
  signal type_cast_1119_inst_req_0 : boolean;
  signal type_cast_1119_inst_ack_0 : boolean;
  signal binary_1125_inst_req_0 : boolean;
  signal binary_1125_inst_ack_0 : boolean;
  signal binary_1125_inst_req_1 : boolean;
  signal binary_1125_inst_ack_1 : boolean;
  signal binary_1131_inst_req_0 : boolean;
  signal binary_1131_inst_ack_0 : boolean;
  signal binary_1131_inst_req_1 : boolean;
  signal binary_1131_inst_ack_1 : boolean;
  signal binary_1137_inst_req_0 : boolean;
  signal binary_1137_inst_ack_0 : boolean;
  signal binary_1137_inst_req_1 : boolean;
  signal binary_1137_inst_ack_1 : boolean;
  signal type_cast_1142_inst_req_0 : boolean;
  signal type_cast_1142_inst_ack_0 : boolean;
  signal binary_1146_inst_req_0 : boolean;
  signal binary_1146_inst_ack_0 : boolean;
  signal binary_1146_inst_req_1 : boolean;
  signal binary_1146_inst_ack_1 : boolean;
  signal binary_1152_inst_req_0 : boolean;
  signal binary_1152_inst_ack_0 : boolean;
  signal binary_1152_inst_req_1 : boolean;
  signal binary_1152_inst_ack_1 : boolean;
  signal binary_1158_inst_req_0 : boolean;
  signal binary_1158_inst_ack_0 : boolean;
  signal binary_1158_inst_req_1 : boolean;
  signal binary_1158_inst_ack_1 : boolean;
  signal binary_1164_inst_req_0 : boolean;
  signal binary_1164_inst_ack_0 : boolean;
  signal binary_1164_inst_req_1 : boolean;
  signal binary_1164_inst_ack_1 : boolean;
  signal ternary_1170_inst_req_0 : boolean;
  signal ternary_1170_inst_ack_0 : boolean;
  signal type_cast_1174_inst_req_0 : boolean;
  signal type_cast_1174_inst_ack_0 : boolean;
  signal binary_1180_inst_req_0 : boolean;
  signal binary_1180_inst_ack_0 : boolean;
  signal binary_1180_inst_req_1 : boolean;
  signal binary_1180_inst_ack_1 : boolean;
  signal binary_1186_inst_req_0 : boolean;
  signal binary_1186_inst_ack_0 : boolean;
  signal binary_1186_inst_req_1 : boolean;
  signal binary_1186_inst_ack_1 : boolean;
  signal binary_1191_inst_req_0 : boolean;
  signal binary_1191_inst_ack_0 : boolean;
  signal binary_1191_inst_req_1 : boolean;
  signal binary_1191_inst_ack_1 : boolean;
  signal simple_obj_ref_1208_inst_req_0 : boolean;
  signal simple_obj_ref_1208_inst_ack_0 : boolean;
  signal simple_obj_ref_1217_inst_req_0 : boolean;
  signal simple_obj_ref_1217_inst_ack_0 : boolean;
  signal type_cast_1200_inst_req_0 : boolean;
  signal type_cast_1200_inst_ack_0 : boolean;
  signal phi_stmt_1195_req_1 : boolean;
  signal type_cast_1198_inst_req_0 : boolean;
  signal type_cast_1198_inst_ack_0 : boolean;
  signal phi_stmt_1195_req_0 : boolean;
  signal phi_stmt_1195_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  output_port_lookup_CP_5084: Block -- control-path 
    signal cp_elements: BooleanArray(99 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= OrReduce(cp_elements(17) & cp_elements(88));
    cp_elements(3) <= simple_obj_ref_1087_inst_ack_0;
    simple_obj_ref_1096_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= simple_obj_ref_1096_inst_ack_0;
    cp_elements(5) <= cp_elements(4);
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(7) & cp_elements(8));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1102_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= cp_elements(5);
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= binary_1102_inst_ack_0;
    binary_1102_inst_req_1 <= cp_elements(9);
    cp_elements(10) <= binary_1102_inst_ack_1;
    cp_elements(11) <= cp_elements(10);
    cp_elements(12) <= false;
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= cp_elements(10);
    if_stmt_1104_branch_req_0 <= cp_elements(14);
    cp_elements(15) <= cp_elements(14);
    cp_elements(16) <= cp_elements(15);
    cp_elements(17) <= if_stmt_1104_branch_ack_1;
    cp_elements(18) <= cp_elements(15);
    cp_elements(19) <= if_stmt_1104_branch_ack_0;
    cp_elements(20) <= cp_elements(2);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(23));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1115_inst_req_0 <= cp_elements(21);
    cp_elements(22) <= cp_elements(20);
    cp_elements(23) <= cp_elements(20);
    cp_elements(24) <= binary_1115_inst_ack_0;
    binary_1115_inst_req_1 <= cp_elements(24);
    cp_elements(25) <= binary_1115_inst_ack_1;
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(28));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1119_inst_req_0 <= cp_elements(26);
    cp_elements(27) <= cp_elements(20);
    cp_elements(28) <= cp_elements(25);
    cp_elements(29) <= type_cast_1119_inst_ack_0;
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(29) & cp_elements(31));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1125_inst_req_0 <= cp_elements(30);
    cp_elements(31) <= cp_elements(20);
    cp_elements(32) <= binary_1125_inst_ack_0;
    binary_1125_inst_req_1 <= cp_elements(32);
    cp_elements(33) <= binary_1125_inst_ack_1;
    cpelement_group_34 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(33) & cp_elements(35));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(34),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1131_inst_req_0 <= cp_elements(34);
    cp_elements(35) <= cp_elements(20);
    cp_elements(36) <= binary_1131_inst_ack_0;
    binary_1131_inst_req_1 <= cp_elements(36);
    cp_elements(37) <= binary_1131_inst_ack_1;
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(39) & cp_elements(40));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1137_inst_req_0 <= cp_elements(38);
    cp_elements(39) <= cp_elements(20);
    cp_elements(40) <= cp_elements(25);
    cp_elements(41) <= binary_1137_inst_ack_0;
    binary_1137_inst_req_1 <= cp_elements(41);
    cp_elements(42) <= binary_1137_inst_ack_1;
    cpelement_group_43 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(44) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(43),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1146_inst_req_0 <= cp_elements(43);
    cp_elements(44) <= cp_elements(20);
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(46));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1142_inst_req_0 <= cp_elements(45);
    cp_elements(46) <= cp_elements(20);
    cp_elements(47) <= type_cast_1142_inst_ack_0;
    cp_elements(48) <= binary_1146_inst_ack_0;
    binary_1146_inst_req_1 <= cp_elements(48);
    cp_elements(49) <= binary_1146_inst_ack_1;
    cpelement_group_50 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(52));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(50),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1152_inst_req_0 <= cp_elements(50);
    cp_elements(51) <= cp_elements(20);
    cp_elements(52) <= cp_elements(37);
    cp_elements(53) <= binary_1152_inst_ack_0;
    binary_1152_inst_req_1 <= cp_elements(53);
    cp_elements(54) <= binary_1152_inst_ack_1;
    cpelement_group_55 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(54) & cp_elements(56));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(55),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1158_inst_req_0 <= cp_elements(55);
    cp_elements(56) <= cp_elements(20);
    cp_elements(57) <= binary_1158_inst_ack_0;
    binary_1158_inst_req_1 <= cp_elements(57);
    cp_elements(58) <= binary_1158_inst_ack_1;
    cpelement_group_59 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(61));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(59),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1164_inst_req_0 <= cp_elements(59);
    cp_elements(60) <= cp_elements(20);
    cp_elements(61) <= cp_elements(37);
    cp_elements(62) <= binary_1164_inst_ack_0;
    binary_1164_inst_req_1 <= cp_elements(62);
    cp_elements(63) <= binary_1164_inst_ack_1;
    cp_elements(64) <= cp_elements(20);
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(49) & cp_elements(58) & cp_elements(63) & cp_elements(64));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ternary_1170_inst_req_0 <= cp_elements(65);
    cp_elements(66) <= ternary_1170_inst_ack_0;
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1174_inst_req_0 <= cp_elements(67);
    cp_elements(68) <= cp_elements(20);
    cp_elements(69) <= type_cast_1174_inst_ack_0;
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(72));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1180_inst_req_0 <= cp_elements(70);
    cp_elements(71) <= cp_elements(20);
    cp_elements(72) <= cp_elements(20);
    cp_elements(73) <= binary_1180_inst_ack_0;
    binary_1180_inst_req_1 <= cp_elements(73);
    cp_elements(74) <= binary_1180_inst_ack_1;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(69) & cp_elements(76));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1186_inst_req_0 <= cp_elements(75);
    cp_elements(76) <= cp_elements(20);
    cp_elements(77) <= binary_1186_inst_ack_0;
    binary_1186_inst_req_1 <= cp_elements(77);
    cp_elements(78) <= binary_1186_inst_ack_1;
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(78) & cp_elements(80));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1191_inst_req_0 <= cp_elements(79);
    cp_elements(80) <= cp_elements(20);
    cp_elements(81) <= binary_1191_inst_ack_0;
    binary_1191_inst_req_1 <= cp_elements(81);
    cp_elements(82) <= binary_1191_inst_ack_1;
    cp_elements(83) <= simple_obj_ref_1208_inst_ack_0;
    simple_obj_ref_1217_inst_req_0 <= cp_elements(83);
    cp_elements(84) <= simple_obj_ref_1217_inst_ack_0;
    cp_elements(85) <= OrReduce(cp_elements(0) & cp_elements(84));
    cp_elements(86) <= cp_elements(85);
    simple_obj_ref_1087_inst_req_0 <= cp_elements(86);
    cp_elements(87) <= false;
    cp_elements(88) <= cp_elements(87);
    cp_elements(89) <= cp_elements(19);
    cp_elements(90) <= cp_elements(19);
    type_cast_1200_inst_req_0 <= cp_elements(90);
    cp_elements(91) <= type_cast_1200_inst_ack_0;
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(91));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1195_req_1 <= cp_elements(92);
    cp_elements(93) <= cp_elements(82);
    type_cast_1198_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= type_cast_1198_inst_ack_0;
    cp_elements(95) <= cp_elements(82);
    cpelement_group_96 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(94) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(96),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1195_req_0 <= cp_elements(96);
    cp_elements(97) <= OrReduce(cp_elements(92) & cp_elements(96));
    cp_elements(98) <= cp_elements(97);
    cp_elements(99) <= phi_stmt_1195_ack_0;
    simple_obj_ref_1208_inst_req_0 <= cp_elements(99);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal datax_x0_1195 : std_logic_vector(63 downto 0);
    signal iNsTr_1_1085 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1094 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1207 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1216 : std_logic_vector(31 downto 0);
    signal tmp10_1147 : std_logic_vector(0 downto 0);
    signal tmp11_1153 : std_logic_vector(31 downto 0);
    signal tmp12_1159 : std_logic_vector(31 downto 0);
    signal tmp13_1165 : std_logic_vector(31 downto 0);
    signal tmp14_1171 : std_logic_vector(31 downto 0);
    signal tmp15_1175 : std_logic_vector(63 downto 0);
    signal tmp16_1181 : std_logic_vector(63 downto 0);
    signal tmp17_1187 : std_logic_vector(63 downto 0);
    signal tmp18_1192 : std_logic_vector(63 downto 0);
    signal tmp2_1088 : std_logic_vector(7 downto 0);
    signal tmp3_1097 : std_logic_vector(63 downto 0);
    signal tmp4_1103 : std_logic_vector(0 downto 0);
    signal tmp6_1116 : std_logic_vector(63 downto 0);
    signal tmp7_1126 : std_logic_vector(31 downto 0);
    signal tmp8_1132 : std_logic_vector(31 downto 0);
    signal tmp9_1138 : std_logic_vector(63 downto 0);
    signal tmp_1120 : std_logic_vector(31 downto 0);
    signal type_cast_1101_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1114_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1129_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1136_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1142_wire : std_logic_vector(63 downto 0);
    signal type_cast_1145_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1151_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1157_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1179_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1185_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1198_wire : std_logic_vector(63 downto 0);
    signal type_cast_1200_wire : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    iNsTr_1_1085 <= "00000000000000000000000000000000";
    iNsTr_2_1094 <= "00000000000000000000000000000000";
    iNsTr_5_1207 <= "00000000000000000000000000000000";
    iNsTr_7_1216 <= "00000000000000000000000000000000";
    type_cast_1101_wire_constant <= "11111111";
    type_cast_1114_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1124_wire_constant <= "00000000000000001111111111111111";
    type_cast_1129_wire_constant <= "00000000000000000000000000000001";
    type_cast_1136_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000001";
    type_cast_1145_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1151_wire_constant <= "00000000000000000000000000000001";
    type_cast_1157_wire_constant <= "00000000000000000111111111111111";
    type_cast_1163_wire_constant <= "00000000000000000000000000000001";
    type_cast_1179_wire_constant <= "0000000000000000111111111111111111111111111111111111111111111111";
    type_cast_1185_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    phi_stmt_1195: Block -- phi operator 
      signal idata: std_logic_vector(127 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1198_wire & type_cast_1200_wire;
      req <= phi_stmt_1195_req_0 & phi_stmt_1195_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 64) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1195_ack_0,
          idata => idata,
          odata => datax_x0_1195,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1195
    ternary_1170_inst: SelectBase generic map(data_width => 32) -- 
      port map( x => tmp12_1159, y => tmp13_1165, sel => tmp10_1147, z => tmp14_1171, req => ternary_1170_inst_req_0, ack => ternary_1170_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1119_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 32, flow_through => false ) 
      port map( din => tmp6_1116, dout => tmp_1120, req => type_cast_1119_inst_req_0, ack => type_cast_1119_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1142_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp9_1138, dout => type_cast_1142_wire, req => type_cast_1142_inst_req_0, ack => type_cast_1142_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1174_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 64, flow_through => false ) 
      port map( din => tmp14_1171, dout => tmp15_1175, req => type_cast_1174_inst_req_0, ack => type_cast_1174_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1198_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp18_1192, dout => type_cast_1198_wire, req => type_cast_1198_inst_req_0, ack => type_cast_1198_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1200_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 64, flow_through => true ) 
      port map( din => tmp3_1097, dout => type_cast_1200_wire, req => type_cast_1200_inst_req_0, ack => type_cast_1200_inst_ack_0, clk => clk, reset => reset); -- 
    if_stmt_1104_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp4_1103;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1104_branch_req_0,
          ack0 => if_stmt_1104_branch_ack_0,
          ack1 => if_stmt_1104_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : binary_1102_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_1088;
      tmp4_1103 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1102_inst_req_0,
          ackL => binary_1102_inst_ack_0,
          reqR => binary_1102_inst_req_1,
          ackR => binary_1102_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_1115_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp3_1097;
      tmp6_1116 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1115_inst_req_0,
          ackL => binary_1115_inst_ack_0,
          reqR => binary_1115_inst_req_1,
          ackR => binary_1115_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_1125_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1120;
      tmp7_1126 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1125_inst_req_0,
          ackL => binary_1125_inst_ack_0,
          reqR => binary_1125_inst_req_1,
          ackR => binary_1125_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_1131_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1129_wire_constant & tmp7_1126;
      tmp8_1132 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1131_inst_req_0,
          ackL => binary_1131_inst_ack_0,
          reqR => binary_1131_inst_req_1,
          ackR => binary_1131_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_1137_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_1116;
      tmp9_1138 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000001",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1137_inst_req_0,
          ackL => binary_1137_inst_ack_0,
          reqR => binary_1137_inst_req_1,
          ackR => binary_1137_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_1146_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1142_wire;
      tmp10_1147 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000000000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1146_inst_req_0,
          ackL => binary_1146_inst_ack_0,
          reqR => binary_1146_inst_req_1,
          ackR => binary_1146_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_1152_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp8_1132;
      tmp11_1153 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1152_inst_req_0,
          ackL => binary_1152_inst_ack_0,
          reqR => binary_1152_inst_req_1,
          ackR => binary_1152_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_1158_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_1153;
      tmp12_1159 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1158_inst_req_0,
          ackL => binary_1158_inst_ack_0,
          reqR => binary_1158_inst_req_1,
          ackR => binary_1158_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_1164_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp8_1132;
      tmp13_1165 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1164_inst_req_0,
          ackL => binary_1164_inst_ack_0,
          reqR => binary_1164_inst_req_1,
          ackR => binary_1164_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_1180_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp3_1097;
      tmp16_1181 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000111111111111111111111111111111111111111111111111",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1180_inst_req_0,
          ackL => binary_1180_inst_ack_0,
          reqR => binary_1180_inst_req_1,
          ackR => binary_1180_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_1186_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_1175;
      tmp17_1187 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1186_inst_req_0,
          ackL => binary_1186_inst_ack_0,
          reqR => binary_1186_inst_req_1,
          ackR => binary_1186_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_1191_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp17_1187 & tmp16_1181;
      tmp18_1192 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1191_inst_req_0,
          ackL => binary_1191_inst_ack_0,
          reqR => binary_1191_inst_req_1,
          ackR => binary_1191_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared inport operator group (0) : simple_obj_ref_1087_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1087_inst_req_0;
      simple_obj_ref_1087_inst_ack_0 <= ack(0);
      tmp2_1088 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => op_lut_ctrl_pipe_read_req(0),
          oack => op_lut_ctrl_pipe_read_ack(0),
          odata => op_lut_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1096_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1096_inst_req_0;
      simple_obj_ref_1096_inst_ack_0 <= ack(0);
      tmp3_1097 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => op_lut_data_pipe_read_req(0),
          oack => op_lut_data_pipe_read_ack(0),
          odata => op_lut_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared outport operator group (0) : simple_obj_ref_1208_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1208_inst_req_0;
      simple_obj_ref_1208_inst_ack_0 <= ack(0);
      data_in <= tmp2_1088;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_ctrl_pipe_write_req(0),
          oack => out_ctrl_pipe_write_ack(0),
          odata => out_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_1217_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1217_inst_req_0;
      simple_obj_ref_1217_inst_ack_0 <= ack(0);
      data_in <= datax_x0_1195;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_3_sr_req : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(87 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(7 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(15 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
    free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
    in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    last_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    last_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    last_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    pkt_length_pipe_write_req : out  std_logic_vector(0 downto 0);
    pkt_length_pipe_write_ack : in   std_logic_vector(0 downto 0);
    pkt_length_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_input;
architecture Default of wrapper_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_input_CP_5456_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_1472_addr_0_req_0 : boolean;
  signal array_obj_ref_1307_root_address_inst_req_0 : boolean;
  signal binary_1489_inst_ack_1 : boolean;
  signal array_obj_ref_1807_root_address_inst_ack_0 : boolean;
  signal binary_1525_inst_ack_0 : boolean;
  signal array_obj_ref_1302_root_address_inst_ack_1 : boolean;
  signal type_cast_1469_inst_ack_0 : boolean;
  signal binary_1519_inst_ack_1 : boolean;
  signal ptr_deref_1232_gather_scatter_req_0 : boolean;
  signal ptr_deref_1852_store_0_req_1 : boolean;
  signal array_obj_ref_1307_base_resize_ack_0 : boolean;
  signal ptr_deref_1458_store_0_ack_0 : boolean;
  signal ptr_deref_1458_store_0_req_1 : boolean;
  signal ptr_deref_1444_gather_scatter_ack_0 : boolean;
  signal binary_1525_inst_req_1 : boolean;
  signal array_obj_ref_1533_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1292_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1292_final_reg_req_0 : boolean;
  signal binary_1525_inst_ack_1 : boolean;
  signal array_obj_ref_1297_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1302_final_reg_ack_0 : boolean;
  signal ptr_deref_1480_store_0_req_1 : boolean;
  signal ptr_deref_1458_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1232_store_0_req_0 : boolean;
  signal ptr_deref_1232_store_0_req_1 : boolean;
  signal array_obj_ref_1292_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1316_root_address_inst_req_0 : boolean;
  signal binary_1519_inst_req_0 : boolean;
  signal array_obj_ref_1292_root_address_inst_ack_1 : boolean;
  signal binary_1489_inst_ack_0 : boolean;
  signal binary_1489_inst_req_0 : boolean;
  signal simple_obj_ref_1255_inst_ack_0 : boolean;
  signal binary_1501_inst_ack_0 : boolean;
  signal array_obj_ref_1807_root_address_inst_req_0 : boolean;
  signal ptr_deref_1458_addr_0_ack_0 : boolean;
  signal binary_1519_inst_ack_0 : boolean;
  signal array_obj_ref_1292_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1537_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1307_base_resize_req_0 : boolean;
  signal binary_1451_inst_req_0 : boolean;
  signal array_obj_ref_1307_root_address_inst_req_1 : boolean;
  signal binary_1501_inst_req_0 : boolean;
  signal array_obj_ref_1297_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1302_root_address_inst_req_1 : boolean;
  signal ptr_deref_1444_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1297_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_store_0_ack_0 : boolean;
  signal binary_1519_inst_req_1 : boolean;
  signal ptr_deref_1472_base_resize_ack_0 : boolean;
  signal ptr_deref_1458_store_0_ack_1 : boolean;
  signal ptr_deref_1232_store_0_ack_1 : boolean;
  signal binary_1501_inst_ack_1 : boolean;
  signal ptr_deref_1232_store_0_ack_0 : boolean;
  signal array_obj_ref_1529_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1537_offset_inst_req_0 : boolean;
  signal array_obj_ref_1292_base_resize_ack_0 : boolean;
  signal if_stmt_1263_branch_req_0 : boolean;
  signal array_obj_ref_1302_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1292_base_resize_req_0 : boolean;
  signal ptr_deref_1444_addr_0_ack_0 : boolean;
  signal array_obj_ref_1529_final_reg_ack_0 : boolean;
  signal binary_1501_inst_req_1 : boolean;
  signal binary_1489_inst_req_1 : boolean;
  signal array_obj_ref_1292_final_reg_ack_0 : boolean;
  signal ptr_deref_1458_gather_scatter_req_0 : boolean;
  signal binary_1525_inst_req_0 : boolean;
  signal simple_obj_ref_1255_inst_req_0 : boolean;
  signal simple_obj_ref_1277_inst_ack_0 : boolean;
  signal array_obj_ref_1307_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1537_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1316_base_resize_req_0 : boolean;
  signal array_obj_ref_1529_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1232_gather_scatter_ack_0 : boolean;
  signal type_cast_1469_inst_req_0 : boolean;
  signal binary_1793_inst_ack_1 : boolean;
  signal binary_1817_inst_ack_1 : boolean;
  signal array_obj_ref_1316_base_resize_ack_0 : boolean;
  signal array_obj_ref_1326_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1472_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1297_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1533_final_reg_ack_0 : boolean;
  signal ptr_deref_1458_base_resize_req_0 : boolean;
  signal array_obj_ref_1529_base_resize_req_0 : boolean;
  signal array_obj_ref_1316_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1541_base_resize_ack_0 : boolean;
  signal ptr_deref_1444_addr_0_req_0 : boolean;
  signal array_obj_ref_1316_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1297_base_resize_req_0 : boolean;
  signal array_obj_ref_1302_final_reg_req_0 : boolean;
  signal array_obj_ref_1529_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1541_offset_inst_req_0 : boolean;
  signal binary_1817_inst_req_0 : boolean;
  signal type_cast_1311_inst_req_0 : boolean;
  signal ptr_deref_1834_store_0_ack_1 : boolean;
  signal array_obj_ref_1316_root_address_inst_ack_1 : boolean;
  signal binary_1495_inst_ack_1 : boolean;
  signal array_obj_ref_1307_final_reg_ack_0 : boolean;
  signal array_obj_ref_1297_base_resize_ack_0 : boolean;
  signal ptr_deref_1458_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_store_0_req_0 : boolean;
  signal array_obj_ref_1316_final_reg_ack_0 : boolean;
  signal array_obj_ref_1307_final_reg_req_0 : boolean;
  signal binary_1451_inst_req_1 : boolean;
  signal binary_1495_inst_req_1 : boolean;
  signal type_cast_1311_inst_ack_0 : boolean;
  signal simple_obj_ref_1244_inst_req_0 : boolean;
  signal ptr_deref_1458_root_address_inst_req_0 : boolean;
  signal if_stmt_1263_branch_ack_1 : boolean;
  signal simple_obj_ref_1244_inst_ack_0 : boolean;
  signal binary_1495_inst_ack_0 : boolean;
  signal binary_1495_inst_req_0 : boolean;
  signal array_obj_ref_1533_root_address_inst_req_1 : boolean;
  signal ptr_deref_1480_store_0_ack_1 : boolean;
  signal ptr_deref_1472_root_address_inst_req_0 : boolean;
  signal type_cast_1797_inst_req_0 : boolean;
  signal binary_1451_inst_ack_0 : boolean;
  signal array_obj_ref_1533_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1302_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1297_final_reg_req_0 : boolean;
  signal if_stmt_1263_branch_ack_0 : boolean;
  signal array_obj_ref_1541_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1537_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1326_root_address_inst_req_1 : boolean;
  signal ptr_deref_1444_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1277_inst_req_0 : boolean;
  signal array_obj_ref_1326_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1529_offset_inst_ack_0 : boolean;
  signal binary_1261_inst_ack_1 : boolean;
  signal array_obj_ref_1529_final_reg_req_0 : boolean;
  signal ptr_deref_1480_addr_0_ack_0 : boolean;
  signal array_obj_ref_1533_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1537_base_resize_ack_0 : boolean;
  signal binary_1261_inst_req_1 : boolean;
  signal ptr_deref_1480_root_address_inst_req_0 : boolean;
  signal binary_1261_inst_ack_0 : boolean;
  signal type_cast_1287_inst_ack_0 : boolean;
  signal binary_1859_inst_ack_0 : boolean;
  signal array_obj_ref_1533_offset_inst_req_0 : boolean;
  signal binary_1507_inst_req_0 : boolean;
  signal type_cast_1287_inst_req_0 : boolean;
  signal array_obj_ref_1326_final_reg_ack_0 : boolean;
  signal ptr_deref_1852_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_base_resize_ack_0 : boolean;
  signal binary_1261_inst_req_0 : boolean;
  signal array_obj_ref_1321_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1321_base_resize_req_0 : boolean;
  signal array_obj_ref_1533_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1326_final_reg_req_0 : boolean;
  signal array_obj_ref_1529_offset_inst_req_0 : boolean;
  signal binary_1507_inst_ack_0 : boolean;
  signal binary_1507_inst_req_1 : boolean;
  signal array_obj_ref_1533_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1321_root_address_inst_req_1 : boolean;
  signal ptr_deref_1444_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1326_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_base_resize_req_0 : boolean;
  signal binary_1817_inst_req_1 : boolean;
  signal array_obj_ref_1831_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1834_store_0_req_1 : boolean;
  signal binary_1507_inst_ack_1 : boolean;
  signal binary_1465_inst_req_0 : boolean;
  signal array_obj_ref_1321_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1480_addr_0_req_0 : boolean;
  signal ptr_deref_1472_addr_0_ack_0 : boolean;
  signal ptr_deref_1458_store_0_req_0 : boolean;
  signal ptr_deref_1458_base_resize_ack_0 : boolean;
  signal array_obj_ref_1529_base_resize_ack_0 : boolean;
  signal array_obj_ref_1321_root_address_inst_req_0 : boolean;
  signal binary_1465_inst_ack_0 : boolean;
  signal array_obj_ref_1326_base_resize_ack_0 : boolean;
  signal array_obj_ref_1831_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1297_final_reg_ack_0 : boolean;
  signal array_obj_ref_1302_base_resize_ack_0 : boolean;
  signal array_obj_ref_1537_index_0_resize_ack_0 : boolean;
  signal binary_1465_inst_req_1 : boolean;
  signal ptr_deref_1444_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1321_final_reg_ack_0 : boolean;
  signal array_obj_ref_1321_final_reg_req_0 : boolean;
  signal ptr_deref_1458_addr_0_req_0 : boolean;
  signal array_obj_ref_1326_base_resize_req_0 : boolean;
  signal array_obj_ref_1302_base_resize_req_0 : boolean;
  signal binary_1465_inst_ack_1 : boolean;
  signal array_obj_ref_1533_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1852_base_resize_req_0 : boolean;
  signal type_cast_1282_inst_ack_0 : boolean;
  signal type_cast_1282_inst_req_0 : boolean;
  signal ptr_deref_1444_store_0_req_0 : boolean;
  signal binary_1451_inst_ack_1 : boolean;
  signal array_obj_ref_1529_root_address_inst_req_1 : boolean;
  signal ptr_deref_1852_base_resize_ack_0 : boolean;
  signal array_obj_ref_1316_final_reg_req_0 : boolean;
  signal ptr_deref_1444_store_0_ack_0 : boolean;
  signal array_obj_ref_1533_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1472_base_resize_req_0 : boolean;
  signal array_obj_ref_1537_root_address_inst_req_0 : boolean;
  signal ptr_deref_1472_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1321_base_resize_ack_0 : boolean;
  signal array_obj_ref_1831_root_address_inst_req_1 : boolean;
  signal ptr_deref_1480_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1307_root_address_inst_ack_0 : boolean;
  signal binary_1513_inst_req_0 : boolean;
  signal binary_1513_inst_ack_0 : boolean;
  signal ptr_deref_1444_store_0_req_1 : boolean;
  signal binary_1513_inst_req_1 : boolean;
  signal array_obj_ref_1541_root_address_inst_ack_0 : boolean;
  signal type_cast_1797_inst_ack_0 : boolean;
  signal ptr_deref_1472_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1537_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1537_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1537_final_reg_req_0 : boolean;
  signal binary_1513_inst_ack_1 : boolean;
  signal ptr_deref_1444_store_0_ack_1 : boolean;
  signal binary_1859_inst_req_0 : boolean;
  signal array_obj_ref_1541_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1537_final_reg_ack_0 : boolean;
  signal array_obj_ref_1533_base_resize_req_0 : boolean;
  signal ptr_deref_1834_store_0_ack_0 : boolean;
  signal array_obj_ref_1533_base_resize_ack_0 : boolean;
  signal array_obj_ref_1537_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1831_offset_inst_req_0 : boolean;
  signal array_obj_ref_1533_index_0_resize_req_0 : boolean;
  signal ptr_deref_1852_addr_0_ack_0 : boolean;
  signal binary_1342_inst_req_0 : boolean;
  signal array_obj_ref_1529_index_0_rename_ack_0 : boolean;
  signal binary_1342_inst_ack_0 : boolean;
  signal binary_1342_inst_req_1 : boolean;
  signal ptr_deref_1444_base_resize_req_0 : boolean;
  signal binary_1342_inst_ack_1 : boolean;
  signal array_obj_ref_1541_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1529_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1541_index_0_rename_ack_0 : boolean;
  signal simple_obj_ref_1351_inst_req_0 : boolean;
  signal simple_obj_ref_1351_inst_ack_0 : boolean;
  signal array_obj_ref_1533_final_reg_req_0 : boolean;
  signal array_obj_ref_1541_final_reg_ack_0 : boolean;
  signal ptr_deref_1834_store_0_req_0 : boolean;
  signal array_obj_ref_1541_final_reg_req_0 : boolean;
  signal array_obj_ref_1541_index_0_rename_req_0 : boolean;
  signal simple_obj_ref_1885_inst_req_0 : boolean;
  signal simple_obj_ref_1360_inst_req_0 : boolean;
  signal simple_obj_ref_1360_inst_ack_0 : boolean;
  signal array_obj_ref_1537_base_resize_req_0 : boolean;
  signal array_obj_ref_1529_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1537_index_0_resize_req_0 : boolean;
  signal type_cast_1364_inst_req_0 : boolean;
  signal array_obj_ref_1529_index_0_resize_req_0 : boolean;
  signal type_cast_1364_inst_ack_0 : boolean;
  signal type_cast_1336_inst_req_0 : boolean;
  signal switch_stmt_1366_branch_default_req_0 : boolean;
  signal binary_1793_inst_req_1 : boolean;
  signal switch_stmt_1366_select_expr_0_req_0 : boolean;
  signal switch_stmt_1366_select_expr_0_ack_0 : boolean;
  signal switch_stmt_1366_select_expr_0_req_1 : boolean;
  signal switch_stmt_1366_select_expr_0_ack_1 : boolean;
  signal type_cast_1477_inst_ack_0 : boolean;
  signal switch_stmt_1366_branch_0_req_0 : boolean;
  signal binary_1817_inst_ack_0 : boolean;
  signal switch_stmt_1366_select_expr_1_req_0 : boolean;
  signal switch_stmt_1366_select_expr_1_ack_0 : boolean;
  signal type_cast_1477_inst_req_0 : boolean;
  signal switch_stmt_1366_select_expr_1_req_1 : boolean;
  signal switch_stmt_1366_select_expr_1_ack_1 : boolean;
  signal switch_stmt_1366_branch_1_req_0 : boolean;
  signal switch_stmt_1366_branch_0_ack_1 : boolean;
  signal binary_1859_inst_req_1 : boolean;
  signal switch_stmt_1366_branch_1_ack_1 : boolean;
  signal ptr_deref_1852_addr_0_req_0 : boolean;
  signal array_obj_ref_1541_index_0_resize_ack_0 : boolean;
  signal switch_stmt_1366_branch_default_ack_0 : boolean;
  signal array_obj_ref_1541_index_0_resize_req_0 : boolean;
  signal binary_1793_inst_ack_0 : boolean;
  signal type_cast_1455_inst_ack_0 : boolean;
  signal binary_1381_inst_req_0 : boolean;
  signal binary_1381_inst_ack_0 : boolean;
  signal binary_1793_inst_req_0 : boolean;
  signal binary_1381_inst_req_1 : boolean;
  signal binary_1381_inst_ack_1 : boolean;
  signal type_cast_1455_inst_req_0 : boolean;
  signal type_cast_1385_inst_req_0 : boolean;
  signal type_cast_1385_inst_ack_0 : boolean;
  signal ptr_deref_1472_store_0_ack_1 : boolean;
  signal ptr_deref_1472_store_0_req_1 : boolean;
  signal array_obj_ref_1831_base_resize_req_0 : boolean;
  signal ptr_deref_1388_base_resize_req_0 : boolean;
  signal ptr_deref_1388_base_resize_ack_0 : boolean;
  signal array_obj_ref_1541_base_resize_req_0 : boolean;
  signal ptr_deref_1388_root_address_inst_req_0 : boolean;
  signal ptr_deref_1388_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1388_addr_0_req_0 : boolean;
  signal ptr_deref_1388_addr_0_ack_0 : boolean;
  signal ptr_deref_1388_gather_scatter_req_0 : boolean;
  signal ptr_deref_1388_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1472_store_0_ack_0 : boolean;
  signal array_obj_ref_1541_offset_inst_ack_0 : boolean;
  signal ptr_deref_1388_store_0_req_0 : boolean;
  signal ptr_deref_1472_store_0_req_0 : boolean;
  signal ptr_deref_1388_store_0_ack_0 : boolean;
  signal ptr_deref_1388_store_0_req_1 : boolean;
  signal ptr_deref_1388_store_0_ack_1 : boolean;
  signal array_obj_ref_1831_base_resize_ack_0 : boolean;
  signal binary_1395_inst_req_0 : boolean;
  signal binary_1395_inst_ack_0 : boolean;
  signal binary_1395_inst_req_1 : boolean;
  signal array_obj_ref_1711_offset_inst_req_0 : boolean;
  signal binary_1395_inst_ack_1 : boolean;
  signal binary_1731_inst_req_0 : boolean;
  signal ptr_deref_1714_store_0_ack_1 : boolean;
  signal array_obj_ref_1711_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1711_root_address_inst_ack_1 : boolean;
  signal type_cast_1399_inst_req_0 : boolean;
  signal type_cast_1399_inst_ack_0 : boolean;
  signal array_obj_ref_1711_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1711_final_reg_req_0 : boolean;
  signal array_obj_ref_1711_final_reg_ack_0 : boolean;
  signal binary_1721_inst_ack_0 : boolean;
  signal ptr_deref_1714_addr_0_ack_0 : boolean;
  signal ptr_deref_1402_base_resize_req_0 : boolean;
  signal ptr_deref_1402_base_resize_ack_0 : boolean;
  signal ptr_deref_1714_store_0_req_1 : boolean;
  signal ptr_deref_1402_root_address_inst_req_0 : boolean;
  signal ptr_deref_1402_root_address_inst_ack_0 : boolean;
  signal binary_1731_inst_ack_1 : boolean;
  signal ptr_deref_1402_addr_0_req_0 : boolean;
  signal array_obj_ref_1711_base_resize_req_0 : boolean;
  signal ptr_deref_1402_addr_0_ack_0 : boolean;
  signal ptr_deref_1402_gather_scatter_req_0 : boolean;
  signal ptr_deref_1714_gather_scatter_req_0 : boolean;
  signal ptr_deref_1402_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1714_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1402_store_0_req_0 : boolean;
  signal ptr_deref_1402_store_0_ack_0 : boolean;
  signal array_obj_ref_1711_base_resize_ack_0 : boolean;
  signal binary_1721_inst_req_1 : boolean;
  signal ptr_deref_1402_store_0_req_1 : boolean;
  signal ptr_deref_1402_store_0_ack_1 : boolean;
  signal binary_1731_inst_ack_0 : boolean;
  signal array_obj_ref_1735_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1852_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1711_root_address_inst_req_0 : boolean;
  signal binary_1731_inst_req_1 : boolean;
  signal binary_1409_inst_req_0 : boolean;
  signal binary_1409_inst_ack_0 : boolean;
  signal binary_1409_inst_req_1 : boolean;
  signal binary_1409_inst_ack_1 : boolean;
  signal array_obj_ref_1735_index_0_resize_req_0 : boolean;
  signal binary_1721_inst_ack_1 : boolean;
  signal array_obj_ref_1711_index_0_resize_req_0 : boolean;
  signal ptr_deref_1714_store_0_req_0 : boolean;
  signal array_obj_ref_1711_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1714_store_0_ack_0 : boolean;
  signal ptr_deref_1714_addr_0_req_0 : boolean;
  signal type_cast_1413_inst_req_0 : boolean;
  signal type_cast_1413_inst_ack_0 : boolean;
  signal binary_1721_inst_req_0 : boolean;
  signal ptr_deref_1714_base_resize_req_0 : boolean;
  signal ptr_deref_1714_base_resize_ack_0 : boolean;
  signal ptr_deref_1416_base_resize_req_0 : boolean;
  signal ptr_deref_1714_root_address_inst_req_0 : boolean;
  signal ptr_deref_1416_base_resize_ack_0 : boolean;
  signal type_cast_1725_inst_req_0 : boolean;
  signal ptr_deref_1416_root_address_inst_req_0 : boolean;
  signal ptr_deref_1416_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1714_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1416_addr_0_req_0 : boolean;
  signal ptr_deref_1416_addr_0_ack_0 : boolean;
  signal type_cast_1725_inst_ack_0 : boolean;
  signal array_obj_ref_1711_index_0_rename_req_0 : boolean;
  signal ptr_deref_1416_gather_scatter_req_0 : boolean;
  signal ptr_deref_1416_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1416_store_0_req_0 : boolean;
  signal ptr_deref_1416_store_0_ack_0 : boolean;
  signal ptr_deref_1416_store_0_req_1 : boolean;
  signal ptr_deref_1416_store_0_ack_1 : boolean;
  signal array_obj_ref_1807_root_address_inst_ack_1 : boolean;
  signal binary_1423_inst_req_0 : boolean;
  signal binary_1423_inst_ack_0 : boolean;
  signal binary_1423_inst_req_1 : boolean;
  signal binary_1423_inst_ack_1 : boolean;
  signal type_cast_1427_inst_req_0 : boolean;
  signal type_cast_1427_inst_ack_0 : boolean;
  signal ptr_deref_1430_base_resize_req_0 : boolean;
  signal ptr_deref_1430_base_resize_ack_0 : boolean;
  signal ptr_deref_1430_root_address_inst_req_0 : boolean;
  signal ptr_deref_1430_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1430_addr_0_req_0 : boolean;
  signal ptr_deref_1430_addr_0_ack_0 : boolean;
  signal ptr_deref_1430_gather_scatter_req_0 : boolean;
  signal ptr_deref_1430_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1430_store_0_req_0 : boolean;
  signal ptr_deref_1430_store_0_ack_0 : boolean;
  signal ptr_deref_1430_store_0_req_1 : boolean;
  signal ptr_deref_1430_store_0_ack_1 : boolean;
  signal binary_1437_inst_req_0 : boolean;
  signal binary_1437_inst_ack_0 : boolean;
  signal binary_1437_inst_req_1 : boolean;
  signal binary_1437_inst_ack_1 : boolean;
  signal type_cast_1441_inst_req_0 : boolean;
  signal type_cast_1441_inst_ack_0 : boolean;
  signal array_obj_ref_1545_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1545_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1545_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1545_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1545_offset_inst_req_0 : boolean;
  signal array_obj_ref_1545_offset_inst_ack_0 : boolean;
  signal binary_1859_inst_ack_1 : boolean;
  signal array_obj_ref_1545_base_resize_req_0 : boolean;
  signal array_obj_ref_1545_base_resize_ack_0 : boolean;
  signal binary_1803_inst_req_0 : boolean;
  signal array_obj_ref_1545_root_address_inst_req_0 : boolean;
  signal binary_1803_inst_ack_0 : boolean;
  signal array_obj_ref_1545_root_address_inst_ack_0 : boolean;
  signal type_cast_1839_inst_req_0 : boolean;
  signal array_obj_ref_1545_root_address_inst_req_1 : boolean;
  signal binary_1803_inst_req_1 : boolean;
  signal array_obj_ref_1545_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1545_final_reg_req_0 : boolean;
  signal simple_obj_ref_1876_inst_req_0 : boolean;
  signal array_obj_ref_1545_final_reg_ack_0 : boolean;
  signal binary_1803_inst_ack_1 : boolean;
  signal type_cast_1839_inst_ack_0 : boolean;
  signal simple_obj_ref_1876_inst_ack_0 : boolean;
  signal array_obj_ref_1831_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1549_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1549_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1549_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1549_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1549_offset_inst_req_0 : boolean;
  signal array_obj_ref_1549_offset_inst_ack_0 : boolean;
  signal type_cast_1821_inst_req_0 : boolean;
  signal type_cast_1821_inst_ack_0 : boolean;
  signal array_obj_ref_1549_base_resize_req_0 : boolean;
  signal array_obj_ref_1549_base_resize_ack_0 : boolean;
  signal array_obj_ref_1807_final_reg_req_0 : boolean;
  signal array_obj_ref_1549_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1549_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1549_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1549_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1549_final_reg_req_0 : boolean;
  signal array_obj_ref_1549_final_reg_ack_0 : boolean;
  signal binary_1845_inst_req_0 : boolean;
  signal binary_1845_inst_ack_0 : boolean;
  signal binary_1845_inst_req_1 : boolean;
  signal binary_1845_inst_ack_1 : boolean;
  signal array_obj_ref_1553_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1553_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1807_final_reg_ack_0 : boolean;
  signal array_obj_ref_1553_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1553_index_0_rename_ack_0 : boolean;
  signal simple_obj_ref_1885_inst_ack_0 : boolean;
  signal array_obj_ref_1553_offset_inst_req_0 : boolean;
  signal array_obj_ref_1553_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1553_base_resize_req_0 : boolean;
  signal array_obj_ref_1553_base_resize_ack_0 : boolean;
  signal array_obj_ref_1553_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1553_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1553_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1553_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1553_final_reg_req_0 : boolean;
  signal array_obj_ref_1553_final_reg_ack_0 : boolean;
  signal binary_1827_inst_req_0 : boolean;
  signal binary_1827_inst_ack_0 : boolean;
  signal array_obj_ref_1557_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1557_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1852_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1557_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1557_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1849_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1557_offset_inst_req_0 : boolean;
  signal array_obj_ref_1557_offset_inst_ack_0 : boolean;
  signal binary_1827_inst_req_1 : boolean;
  signal array_obj_ref_1557_base_resize_req_0 : boolean;
  signal array_obj_ref_1557_base_resize_ack_0 : boolean;
  signal array_obj_ref_1849_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1557_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1557_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1557_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1557_root_address_inst_ack_1 : boolean;
  signal phi_stmt_1330_ack_0 : boolean;
  signal array_obj_ref_1849_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1557_final_reg_req_0 : boolean;
  signal array_obj_ref_1557_final_reg_ack_0 : boolean;
  signal binary_1827_inst_ack_1 : boolean;
  signal array_obj_ref_1849_index_0_rename_ack_0 : boolean;
  signal binary_1563_inst_req_0 : boolean;
  signal binary_1563_inst_ack_0 : boolean;
  signal binary_1563_inst_req_1 : boolean;
  signal array_obj_ref_1849_offset_inst_req_0 : boolean;
  signal binary_1563_inst_ack_1 : boolean;
  signal ptr_deref_1852_store_0_ack_1 : boolean;
  signal array_obj_ref_1849_offset_inst_ack_0 : boolean;
  signal type_cast_1567_inst_req_0 : boolean;
  signal ptr_deref_1852_store_0_req_0 : boolean;
  signal type_cast_1567_inst_ack_0 : boolean;
  signal array_obj_ref_1807_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1807_index_0_resize_req_0 : boolean;
  signal ptr_deref_1852_store_0_ack_0 : boolean;
  signal array_obj_ref_1849_base_resize_req_0 : boolean;
  signal array_obj_ref_1849_base_resize_ack_0 : boolean;
  signal ptr_deref_1570_base_resize_req_0 : boolean;
  signal ptr_deref_1570_base_resize_ack_0 : boolean;
  signal array_obj_ref_1807_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1570_root_address_inst_req_0 : boolean;
  signal ptr_deref_1570_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1570_addr_0_req_0 : boolean;
  signal ptr_deref_1570_addr_0_ack_0 : boolean;
  signal ptr_deref_1570_gather_scatter_req_0 : boolean;
  signal ptr_deref_1570_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1807_index_0_rename_req_0 : boolean;
  signal ptr_deref_1570_store_0_req_0 : boolean;
  signal ptr_deref_1570_store_0_ack_0 : boolean;
  signal array_obj_ref_1807_index_0_rename_ack_0 : boolean;
  signal ptr_deref_1570_store_0_req_1 : boolean;
  signal ptr_deref_1570_store_0_ack_1 : boolean;
  signal array_obj_ref_1849_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1849_root_address_inst_ack_0 : boolean;
  signal binary_1577_inst_req_0 : boolean;
  signal binary_1577_inst_ack_0 : boolean;
  signal binary_1577_inst_req_1 : boolean;
  signal array_obj_ref_1807_offset_inst_req_0 : boolean;
  signal binary_1577_inst_ack_1 : boolean;
  signal array_obj_ref_1849_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1849_root_address_inst_ack_1 : boolean;
  signal type_cast_1581_inst_req_0 : boolean;
  signal type_cast_1581_inst_ack_0 : boolean;
  signal array_obj_ref_1807_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1849_final_reg_req_0 : boolean;
  signal ptr_deref_1584_base_resize_req_0 : boolean;
  signal array_obj_ref_1849_final_reg_ack_0 : boolean;
  signal ptr_deref_1584_base_resize_ack_0 : boolean;
  signal ptr_deref_1584_root_address_inst_req_0 : boolean;
  signal ptr_deref_1584_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1852_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1584_addr_0_req_0 : boolean;
  signal ptr_deref_1584_addr_0_ack_0 : boolean;
  signal array_obj_ref_1831_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1831_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1584_gather_scatter_req_0 : boolean;
  signal ptr_deref_1584_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1584_store_0_req_0 : boolean;
  signal ptr_deref_1584_store_0_ack_0 : boolean;
  signal ptr_deref_1584_store_0_req_1 : boolean;
  signal ptr_deref_1584_store_0_ack_1 : boolean;
  signal array_obj_ref_1831_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1807_base_resize_req_0 : boolean;
  signal array_obj_ref_1831_index_0_rename_ack_0 : boolean;
  signal binary_1591_inst_req_0 : boolean;
  signal binary_1591_inst_ack_0 : boolean;
  signal array_obj_ref_1807_base_resize_ack_0 : boolean;
  signal binary_1591_inst_req_1 : boolean;
  signal binary_1591_inst_ack_1 : boolean;
  signal type_cast_1595_inst_req_0 : boolean;
  signal type_cast_1595_inst_ack_0 : boolean;
  signal ptr_deref_1598_base_resize_req_0 : boolean;
  signal ptr_deref_1598_base_resize_ack_0 : boolean;
  signal ptr_deref_1598_root_address_inst_req_0 : boolean;
  signal ptr_deref_1598_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1598_addr_0_req_0 : boolean;
  signal ptr_deref_1598_addr_0_ack_0 : boolean;
  signal ptr_deref_1598_gather_scatter_req_0 : boolean;
  signal ptr_deref_1598_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1598_store_0_req_0 : boolean;
  signal ptr_deref_1598_store_0_ack_0 : boolean;
  signal ptr_deref_1598_store_0_req_1 : boolean;
  signal ptr_deref_1598_store_0_ack_1 : boolean;
  signal binary_1605_inst_req_0 : boolean;
  signal binary_1605_inst_ack_0 : boolean;
  signal binary_1605_inst_req_1 : boolean;
  signal binary_1605_inst_ack_1 : boolean;
  signal type_cast_1609_inst_req_0 : boolean;
  signal type_cast_1609_inst_ack_0 : boolean;
  signal ptr_deref_1612_base_resize_req_0 : boolean;
  signal ptr_deref_1612_base_resize_ack_0 : boolean;
  signal ptr_deref_1612_root_address_inst_req_0 : boolean;
  signal ptr_deref_1612_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1612_addr_0_req_0 : boolean;
  signal ptr_deref_1612_addr_0_ack_0 : boolean;
  signal ptr_deref_1612_gather_scatter_req_0 : boolean;
  signal ptr_deref_1612_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1612_store_0_req_0 : boolean;
  signal ptr_deref_1612_store_0_ack_0 : boolean;
  signal ptr_deref_1612_store_0_req_1 : boolean;
  signal ptr_deref_1612_store_0_ack_1 : boolean;
  signal binary_1619_inst_req_0 : boolean;
  signal binary_1619_inst_ack_0 : boolean;
  signal binary_1619_inst_req_1 : boolean;
  signal binary_1619_inst_ack_1 : boolean;
  signal type_cast_1623_inst_req_0 : boolean;
  signal type_cast_1623_inst_ack_0 : boolean;
  signal ptr_deref_1626_base_resize_req_0 : boolean;
  signal ptr_deref_1626_base_resize_ack_0 : boolean;
  signal ptr_deref_1626_root_address_inst_req_0 : boolean;
  signal ptr_deref_1626_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1626_addr_0_req_0 : boolean;
  signal ptr_deref_1626_addr_0_ack_0 : boolean;
  signal ptr_deref_1626_gather_scatter_req_0 : boolean;
  signal ptr_deref_1626_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1626_store_0_req_0 : boolean;
  signal ptr_deref_1626_store_0_ack_0 : boolean;
  signal ptr_deref_1626_store_0_req_1 : boolean;
  signal ptr_deref_1626_store_0_ack_1 : boolean;
  signal binary_1633_inst_req_0 : boolean;
  signal binary_1633_inst_ack_0 : boolean;
  signal binary_1633_inst_req_1 : boolean;
  signal binary_1633_inst_ack_1 : boolean;
  signal type_cast_1637_inst_req_0 : boolean;
  signal type_cast_1637_inst_ack_0 : boolean;
  signal ptr_deref_1640_base_resize_req_0 : boolean;
  signal ptr_deref_1640_base_resize_ack_0 : boolean;
  signal ptr_deref_1640_root_address_inst_req_0 : boolean;
  signal ptr_deref_1640_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1640_addr_0_req_0 : boolean;
  signal ptr_deref_1640_addr_0_ack_0 : boolean;
  signal ptr_deref_1640_gather_scatter_req_0 : boolean;
  signal ptr_deref_1640_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1640_store_0_req_0 : boolean;
  signal ptr_deref_1640_store_0_ack_0 : boolean;
  signal ptr_deref_1640_store_0_req_1 : boolean;
  signal ptr_deref_1640_store_0_ack_1 : boolean;
  signal binary_1647_inst_req_0 : boolean;
  signal binary_1647_inst_ack_0 : boolean;
  signal binary_1647_inst_req_1 : boolean;
  signal binary_1647_inst_ack_1 : boolean;
  signal type_cast_1651_inst_req_0 : boolean;
  signal type_cast_1651_inst_ack_0 : boolean;
  signal ptr_deref_1654_base_resize_req_0 : boolean;
  signal ptr_deref_1654_base_resize_ack_0 : boolean;
  signal ptr_deref_1654_root_address_inst_req_0 : boolean;
  signal ptr_deref_1654_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1654_addr_0_req_0 : boolean;
  signal ptr_deref_1654_addr_0_ack_0 : boolean;
  signal ptr_deref_1654_gather_scatter_req_0 : boolean;
  signal ptr_deref_1654_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1654_store_0_req_0 : boolean;
  signal ptr_deref_1654_store_0_ack_0 : boolean;
  signal ptr_deref_1654_store_0_req_1 : boolean;
  signal ptr_deref_1654_store_0_ack_1 : boolean;
  signal type_cast_1659_inst_req_0 : boolean;
  signal type_cast_1659_inst_ack_0 : boolean;
  signal ptr_deref_1662_base_resize_req_0 : boolean;
  signal ptr_deref_1662_base_resize_ack_0 : boolean;
  signal ptr_deref_1662_root_address_inst_req_0 : boolean;
  signal ptr_deref_1662_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1662_addr_0_req_0 : boolean;
  signal ptr_deref_1662_addr_0_ack_0 : boolean;
  signal ptr_deref_1662_gather_scatter_req_0 : boolean;
  signal ptr_deref_1662_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1662_store_0_req_0 : boolean;
  signal ptr_deref_1662_store_0_ack_0 : boolean;
  signal ptr_deref_1662_store_0_req_1 : boolean;
  signal ptr_deref_1662_store_0_ack_1 : boolean;
  signal binary_1671_inst_req_0 : boolean;
  signal binary_1671_inst_ack_0 : boolean;
  signal binary_1671_inst_req_1 : boolean;
  signal binary_1671_inst_ack_1 : boolean;
  signal binary_1679_inst_req_0 : boolean;
  signal binary_1679_inst_ack_0 : boolean;
  signal binary_1679_inst_req_1 : boolean;
  signal binary_1679_inst_ack_1 : boolean;
  signal type_cast_1683_inst_req_0 : boolean;
  signal type_cast_1683_inst_ack_0 : boolean;
  signal array_obj_ref_1687_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1687_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1687_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1687_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1687_offset_inst_req_0 : boolean;
  signal array_obj_ref_1687_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1687_base_resize_req_0 : boolean;
  signal array_obj_ref_1687_base_resize_ack_0 : boolean;
  signal array_obj_ref_1687_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1687_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1687_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1687_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1687_final_reg_req_0 : boolean;
  signal array_obj_ref_1687_final_reg_ack_0 : boolean;
  signal ptr_deref_1690_base_resize_req_0 : boolean;
  signal ptr_deref_1690_base_resize_ack_0 : boolean;
  signal ptr_deref_1690_root_address_inst_req_0 : boolean;
  signal ptr_deref_1690_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1690_addr_0_req_0 : boolean;
  signal ptr_deref_1690_addr_0_ack_0 : boolean;
  signal ptr_deref_1690_gather_scatter_req_0 : boolean;
  signal ptr_deref_1690_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1690_store_0_req_0 : boolean;
  signal ptr_deref_1690_store_0_ack_0 : boolean;
  signal ptr_deref_1690_store_0_req_1 : boolean;
  signal ptr_deref_1690_store_0_ack_1 : boolean;
  signal binary_1697_inst_req_0 : boolean;
  signal binary_1697_inst_ack_0 : boolean;
  signal binary_1697_inst_req_1 : boolean;
  signal binary_1697_inst_ack_1 : boolean;
  signal type_cast_1701_inst_req_0 : boolean;
  signal type_cast_1701_inst_ack_0 : boolean;
  signal binary_1707_inst_req_0 : boolean;
  signal binary_1707_inst_ack_0 : boolean;
  signal binary_1707_inst_req_1 : boolean;
  signal binary_1707_inst_ack_1 : boolean;
  signal array_obj_ref_1735_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1735_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1735_offset_inst_req_0 : boolean;
  signal array_obj_ref_1735_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1735_base_resize_req_0 : boolean;
  signal array_obj_ref_1735_base_resize_ack_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1735_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1735_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1810_store_0_ack_1 : boolean;
  signal array_obj_ref_1735_final_reg_req_0 : boolean;
  signal ptr_deref_1810_store_0_req_1 : boolean;
  signal array_obj_ref_1735_final_reg_ack_0 : boolean;
  signal ptr_deref_1810_store_0_ack_0 : boolean;
  signal ptr_deref_1738_base_resize_req_0 : boolean;
  signal ptr_deref_1810_store_0_req_0 : boolean;
  signal ptr_deref_1738_base_resize_ack_0 : boolean;
  signal ptr_deref_1834_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1738_root_address_inst_req_0 : boolean;
  signal ptr_deref_1738_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1834_gather_scatter_req_0 : boolean;
  signal ptr_deref_1738_addr_0_req_0 : boolean;
  signal ptr_deref_1738_addr_0_ack_0 : boolean;
  signal ptr_deref_1834_addr_0_ack_0 : boolean;
  signal ptr_deref_1810_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1738_gather_scatter_req_0 : boolean;
  signal ptr_deref_1810_gather_scatter_req_0 : boolean;
  signal ptr_deref_1738_gather_scatter_ack_0 : boolean;
  signal phi_stmt_1330_req_1 : boolean;
  signal ptr_deref_1738_store_0_req_0 : boolean;
  signal ptr_deref_1738_store_0_ack_0 : boolean;
  signal type_cast_1336_inst_ack_0 : boolean;
  signal ptr_deref_1810_addr_0_ack_0 : boolean;
  signal ptr_deref_1738_store_0_req_1 : boolean;
  signal ptr_deref_1810_addr_0_req_0 : boolean;
  signal ptr_deref_1738_store_0_ack_1 : boolean;
  signal ptr_deref_1834_addr_0_req_0 : boolean;
  signal ptr_deref_1810_root_address_inst_ack_0 : boolean;
  signal binary_1745_inst_req_0 : boolean;
  signal binary_1745_inst_ack_0 : boolean;
  signal ptr_deref_1834_root_address_inst_ack_0 : boolean;
  signal binary_1745_inst_req_1 : boolean;
  signal binary_1745_inst_ack_1 : boolean;
  signal ptr_deref_1810_root_address_inst_req_0 : boolean;
  signal ptr_deref_1834_root_address_inst_req_0 : boolean;
  signal ptr_deref_1834_base_resize_ack_0 : boolean;
  signal type_cast_1749_inst_req_0 : boolean;
  signal type_cast_1749_inst_ack_0 : boolean;
  signal ptr_deref_1810_base_resize_ack_0 : boolean;
  signal ptr_deref_1834_base_resize_req_0 : boolean;
  signal ptr_deref_1810_base_resize_req_0 : boolean;
  signal binary_1755_inst_req_0 : boolean;
  signal binary_1755_inst_ack_0 : boolean;
  signal binary_1755_inst_req_1 : boolean;
  signal binary_1755_inst_ack_1 : boolean;
  signal array_obj_ref_1831_final_reg_ack_0 : boolean;
  signal array_obj_ref_1831_final_reg_req_0 : boolean;
  signal array_obj_ref_1759_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1759_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1759_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1759_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1759_offset_inst_req_0 : boolean;
  signal array_obj_ref_1759_offset_inst_ack_0 : boolean;
  signal simple_obj_ref_1867_inst_ack_0 : boolean;
  signal array_obj_ref_1759_base_resize_req_0 : boolean;
  signal simple_obj_ref_1867_inst_req_0 : boolean;
  signal array_obj_ref_1759_base_resize_ack_0 : boolean;
  signal array_obj_ref_1759_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1759_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1831_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1759_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1759_root_address_inst_ack_1 : boolean;
  signal phi_stmt_1330_req_0 : boolean;
  signal array_obj_ref_1759_final_reg_req_0 : boolean;
  signal array_obj_ref_1759_final_reg_ack_0 : boolean;
  signal ptr_deref_1762_base_resize_req_0 : boolean;
  signal ptr_deref_1762_base_resize_ack_0 : boolean;
  signal ptr_deref_1762_root_address_inst_req_0 : boolean;
  signal ptr_deref_1762_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1762_addr_0_req_0 : boolean;
  signal ptr_deref_1762_addr_0_ack_0 : boolean;
  signal ptr_deref_1762_gather_scatter_req_0 : boolean;
  signal ptr_deref_1762_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1762_store_0_req_0 : boolean;
  signal ptr_deref_1762_store_0_ack_0 : boolean;
  signal ptr_deref_1762_store_0_req_1 : boolean;
  signal ptr_deref_1762_store_0_ack_1 : boolean;
  signal binary_1769_inst_req_0 : boolean;
  signal binary_1769_inst_ack_0 : boolean;
  signal binary_1769_inst_req_1 : boolean;
  signal binary_1769_inst_ack_1 : boolean;
  signal type_cast_1773_inst_req_0 : boolean;
  signal type_cast_1773_inst_ack_0 : boolean;
  signal binary_1779_inst_req_0 : boolean;
  signal binary_1779_inst_ack_0 : boolean;
  signal binary_1779_inst_req_1 : boolean;
  signal binary_1779_inst_ack_1 : boolean;
  signal array_obj_ref_1783_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1783_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1783_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1783_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1783_offset_inst_req_0 : boolean;
  signal array_obj_ref_1783_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1783_base_resize_req_0 : boolean;
  signal array_obj_ref_1783_base_resize_ack_0 : boolean;
  signal array_obj_ref_1783_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1783_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1783_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1783_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1783_final_reg_req_0 : boolean;
  signal array_obj_ref_1783_final_reg_ack_0 : boolean;
  signal ptr_deref_1786_base_resize_req_0 : boolean;
  signal ptr_deref_1786_base_resize_ack_0 : boolean;
  signal ptr_deref_1786_root_address_inst_req_0 : boolean;
  signal ptr_deref_1786_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1786_addr_0_req_0 : boolean;
  signal ptr_deref_1786_addr_0_ack_0 : boolean;
  signal ptr_deref_1786_gather_scatter_req_0 : boolean;
  signal ptr_deref_1786_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1786_store_0_req_0 : boolean;
  signal ptr_deref_1786_store_0_ack_0 : boolean;
  signal ptr_deref_1786_store_0_req_1 : boolean;
  signal ptr_deref_1786_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_input_CP_5456: Block -- control-path 
    signal cp_elements: BooleanArray(809 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(17);
    cp_elements(3) <= OrReduce(cp_elements(32) & cp_elements(801));
    simple_obj_ref_1277_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= cp_elements(96);
    phi_stmt_1330_req_0 <= cp_elements(4);
    cp_elements(5) <= OrReduce(cp_elements(124) & cp_elements(807));
    cp_elements(6) <= cp_elements(269);
    cp_elements(7) <= cp_elements(526);
    cp_elements(8) <= cp_elements(794);
    simple_obj_ref_1867_inst_req_0 <= cp_elements(8);
    cp_elements(9) <= cp_elements(0);
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(10) & cp_elements(13));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1232_gather_scatter_req_0 <= cp_elements(11);
    cp_elements(12) <= cp_elements(9);
    cp_elements(13) <= cp_elements(9);
    cp_elements(14) <= ptr_deref_1232_gather_scatter_ack_0;
    ptr_deref_1232_store_0_req_0 <= cp_elements(14);
    cp_elements(15) <= ptr_deref_1232_store_0_ack_0;
    ptr_deref_1232_store_0_req_1 <= cp_elements(15);
    cp_elements(16) <= ptr_deref_1232_store_0_ack_1;
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(16));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(18) <= simple_obj_ref_1244_inst_ack_0;
    simple_obj_ref_1255_inst_req_0 <= cp_elements(18);
    cp_elements(19) <= simple_obj_ref_1255_inst_ack_0;
    cp_elements(20) <= cp_elements(19);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(23));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1261_inst_req_0 <= cp_elements(21);
    cp_elements(22) <= cp_elements(20);
    cp_elements(23) <= cp_elements(20);
    cp_elements(24) <= binary_1261_inst_ack_0;
    binary_1261_inst_req_1 <= cp_elements(24);
    cp_elements(25) <= binary_1261_inst_ack_1;
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= false;
    cp_elements(28) <= cp_elements(27);
    cp_elements(29) <= cp_elements(25);
    if_stmt_1263_branch_req_0 <= cp_elements(29);
    cp_elements(30) <= cp_elements(29);
    cp_elements(31) <= cp_elements(30);
    cp_elements(32) <= if_stmt_1263_branch_ack_1;
    cp_elements(33) <= cp_elements(30);
    cp_elements(34) <= if_stmt_1263_branch_ack_0;
    cp_elements(35) <= simple_obj_ref_1277_inst_ack_0;
    cp_elements(36) <= cp_elements(35);
    cpelement_group_37 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(38) & cp_elements(39));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(37),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1282_inst_req_0 <= cp_elements(37);
    cp_elements(38) <= cp_elements(36);
    cp_elements(39) <= cp_elements(36);
    cp_elements(40) <= type_cast_1282_inst_ack_0;
    array_obj_ref_1307_base_resize_req_0 <= cp_elements(40);
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(43));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1287_inst_req_0 <= cp_elements(41);
    cp_elements(42) <= cp_elements(36);
    cp_elements(43) <= cp_elements(36);
    cp_elements(44) <= type_cast_1287_inst_ack_0;
    cp_elements(45) <= cp_elements(36);
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(50));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1292_final_reg_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(44);
    array_obj_ref_1292_base_resize_req_0 <= cp_elements(47);
    cp_elements(48) <= array_obj_ref_1292_base_resize_ack_0;
    array_obj_ref_1292_root_address_inst_req_0 <= cp_elements(48);
    cp_elements(49) <= array_obj_ref_1292_root_address_inst_ack_0;
    array_obj_ref_1292_root_address_inst_req_1 <= cp_elements(49);
    cp_elements(50) <= array_obj_ref_1292_root_address_inst_ack_1;
    cp_elements(51) <= array_obj_ref_1292_final_reg_ack_0;
    cp_elements(52) <= cp_elements(36);
    cpelement_group_53 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(52) & cp_elements(57));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(53),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1297_final_reg_req_0 <= cp_elements(53);
    cp_elements(54) <= cp_elements(44);
    array_obj_ref_1297_base_resize_req_0 <= cp_elements(54);
    cp_elements(55) <= array_obj_ref_1297_base_resize_ack_0;
    array_obj_ref_1297_root_address_inst_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_1297_root_address_inst_ack_0;
    array_obj_ref_1297_root_address_inst_req_1 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_1297_root_address_inst_ack_1;
    cp_elements(58) <= array_obj_ref_1297_final_reg_ack_0;
    cp_elements(59) <= cp_elements(36);
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(59) & cp_elements(64));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1302_final_reg_req_0 <= cp_elements(60);
    cp_elements(61) <= cp_elements(44);
    array_obj_ref_1302_base_resize_req_0 <= cp_elements(61);
    cp_elements(62) <= array_obj_ref_1302_base_resize_ack_0;
    array_obj_ref_1302_root_address_inst_req_0 <= cp_elements(62);
    cp_elements(63) <= array_obj_ref_1302_root_address_inst_ack_0;
    array_obj_ref_1302_root_address_inst_req_1 <= cp_elements(63);
    cp_elements(64) <= array_obj_ref_1302_root_address_inst_ack_1;
    cp_elements(65) <= array_obj_ref_1302_final_reg_ack_0;
    cp_elements(66) <= cp_elements(36);
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(70));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1307_final_reg_req_0 <= cp_elements(67);
    cp_elements(68) <= array_obj_ref_1307_base_resize_ack_0;
    array_obj_ref_1307_root_address_inst_req_0 <= cp_elements(68);
    cp_elements(69) <= array_obj_ref_1307_root_address_inst_ack_0;
    array_obj_ref_1307_root_address_inst_req_1 <= cp_elements(69);
    cp_elements(70) <= array_obj_ref_1307_root_address_inst_ack_1;
    cp_elements(71) <= array_obj_ref_1307_final_reg_ack_0;
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(73));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1311_inst_req_0 <= cp_elements(72);
    cp_elements(73) <= cp_elements(36);
    cp_elements(74) <= type_cast_1311_inst_ack_0;
    cp_elements(75) <= cp_elements(36);
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(80));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1316_final_reg_req_0 <= cp_elements(76);
    cp_elements(77) <= cp_elements(44);
    array_obj_ref_1316_base_resize_req_0 <= cp_elements(77);
    cp_elements(78) <= array_obj_ref_1316_base_resize_ack_0;
    array_obj_ref_1316_root_address_inst_req_0 <= cp_elements(78);
    cp_elements(79) <= array_obj_ref_1316_root_address_inst_ack_0;
    array_obj_ref_1316_root_address_inst_req_1 <= cp_elements(79);
    cp_elements(80) <= array_obj_ref_1316_root_address_inst_ack_1;
    cp_elements(81) <= array_obj_ref_1316_final_reg_ack_0;
    cp_elements(82) <= cp_elements(36);
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(87));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1321_final_reg_req_0 <= cp_elements(83);
    cp_elements(84) <= cp_elements(44);
    array_obj_ref_1321_base_resize_req_0 <= cp_elements(84);
    cp_elements(85) <= array_obj_ref_1321_base_resize_ack_0;
    array_obj_ref_1321_root_address_inst_req_0 <= cp_elements(85);
    cp_elements(86) <= array_obj_ref_1321_root_address_inst_ack_0;
    array_obj_ref_1321_root_address_inst_req_1 <= cp_elements(86);
    cp_elements(87) <= array_obj_ref_1321_root_address_inst_ack_1;
    cp_elements(88) <= array_obj_ref_1321_final_reg_ack_0;
    cp_elements(89) <= cp_elements(36);
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(94));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1326_final_reg_req_0 <= cp_elements(90);
    cp_elements(91) <= cp_elements(44);
    array_obj_ref_1326_base_resize_req_0 <= cp_elements(91);
    cp_elements(92) <= array_obj_ref_1326_base_resize_ack_0;
    array_obj_ref_1326_root_address_inst_req_0 <= cp_elements(92);
    cp_elements(93) <= array_obj_ref_1326_root_address_inst_ack_0;
    array_obj_ref_1326_root_address_inst_req_1 <= cp_elements(93);
    cp_elements(94) <= array_obj_ref_1326_root_address_inst_ack_1;
    cp_elements(95) <= array_obj_ref_1326_final_reg_ack_0;
    cpelement_group_96 : Block -- 
      signal predecessors: BooleanArray(6 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(58) & cp_elements(65) & cp_elements(74) & cp_elements(81) & cp_elements(88) & cp_elements(95));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(96),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(97) <= cp_elements(805);
    cpelement_group_98 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(99) & cp_elements(100));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(98),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1342_inst_req_0 <= cp_elements(98);
    cp_elements(99) <= cp_elements(97);
    cp_elements(100) <= cp_elements(97);
    cp_elements(101) <= binary_1342_inst_ack_0;
    binary_1342_inst_req_1 <= cp_elements(101);
    cp_elements(102) <= binary_1342_inst_ack_1;
    simple_obj_ref_1351_inst_req_0 <= cp_elements(102);
    cp_elements(103) <= simple_obj_ref_1351_inst_ack_0;
    simple_obj_ref_1360_inst_req_0 <= cp_elements(103);
    cp_elements(104) <= simple_obj_ref_1360_inst_ack_0;
    cp_elements(105) <= cp_elements(104);
    cpelement_group_106 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(107) & cp_elements(108));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(106),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1364_inst_req_0 <= cp_elements(106);
    cp_elements(107) <= cp_elements(105);
    cp_elements(108) <= cp_elements(105);
    cp_elements(109) <= type_cast_1364_inst_ack_0;
    cp_elements(110) <= cp_elements(109);
    cp_elements(111) <= false;
    cp_elements(112) <= cp_elements(111);
    cp_elements(113) <= cp_elements(109);
    cp_elements(114) <= cp_elements(113);
    cp_elements(115) <= cp_elements(114);
    switch_stmt_1366_select_expr_0_req_0 <= cp_elements(115);
    cp_elements(116) <= switch_stmt_1366_select_expr_0_ack_0;
    switch_stmt_1366_select_expr_0_req_1 <= cp_elements(116);
    cp_elements(117) <= switch_stmt_1366_select_expr_0_ack_1;
    switch_stmt_1366_branch_0_req_0 <= cp_elements(117);
    cp_elements(118) <= cp_elements(114);
    switch_stmt_1366_select_expr_1_req_0 <= cp_elements(118);
    cp_elements(119) <= switch_stmt_1366_select_expr_1_ack_0;
    switch_stmt_1366_select_expr_1_req_1 <= cp_elements(119);
    cp_elements(120) <= switch_stmt_1366_select_expr_1_ack_1;
    switch_stmt_1366_branch_1_req_0 <= cp_elements(120);
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(117) & cp_elements(120));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    switch_stmt_1366_branch_default_req_0 <= cp_elements(121);
    cp_elements(122) <= cp_elements(121);
    cp_elements(123) <= cp_elements(122);
    cp_elements(124) <= switch_stmt_1366_branch_0_ack_1;
    cp_elements(125) <= cp_elements(122);
    cp_elements(126) <= switch_stmt_1366_branch_1_ack_1;
    cp_elements(127) <= cp_elements(122);
    cp_elements(128) <= switch_stmt_1366_branch_default_ack_0;
    cp_elements(129) <= cp_elements(5);
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(131) & cp_elements(132));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1381_inst_req_0 <= cp_elements(130);
    cp_elements(131) <= cp_elements(129);
    cp_elements(132) <= cp_elements(129);
    cp_elements(133) <= binary_1381_inst_ack_0;
    binary_1381_inst_req_1 <= cp_elements(133);
    cp_elements(134) <= binary_1381_inst_ack_1;
    cpelement_group_135 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(136));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(135),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1385_inst_req_0 <= cp_elements(135);
    cp_elements(136) <= cp_elements(129);
    cp_elements(137) <= type_cast_1385_inst_ack_0;
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(139) & cp_elements(143));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1388_gather_scatter_req_0 <= cp_elements(138);
    cp_elements(139) <= cp_elements(129);
    cp_elements(140) <= cp_elements(139);
    ptr_deref_1388_base_resize_req_0 <= cp_elements(140);
    cp_elements(141) <= ptr_deref_1388_base_resize_ack_0;
    ptr_deref_1388_root_address_inst_req_0 <= cp_elements(141);
    cp_elements(142) <= ptr_deref_1388_root_address_inst_ack_0;
    ptr_deref_1388_addr_0_req_0 <= cp_elements(142);
    cp_elements(143) <= ptr_deref_1388_addr_0_ack_0;
    cp_elements(144) <= ptr_deref_1388_gather_scatter_ack_0;
    ptr_deref_1388_store_0_req_0 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_1388_store_0_ack_0;
    cp_elements(146) <= cp_elements(145);
    ptr_deref_1388_store_0_req_1 <= cp_elements(146);
    cp_elements(147) <= ptr_deref_1388_store_0_ack_1;
    cpelement_group_148 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(150));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(148),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1395_inst_req_0 <= cp_elements(148);
    cp_elements(149) <= cp_elements(129);
    cp_elements(150) <= cp_elements(129);
    cp_elements(151) <= binary_1395_inst_ack_0;
    binary_1395_inst_req_1 <= cp_elements(151);
    cp_elements(152) <= binary_1395_inst_ack_1;
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1399_inst_req_0 <= cp_elements(153);
    cp_elements(154) <= cp_elements(129);
    cp_elements(155) <= type_cast_1399_inst_ack_0;
    cpelement_group_156 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(145) & cp_elements(155) & cp_elements(157) & cp_elements(161));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(156),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1402_gather_scatter_req_0 <= cp_elements(156);
    cp_elements(157) <= cp_elements(129);
    cp_elements(158) <= cp_elements(157);
    ptr_deref_1402_base_resize_req_0 <= cp_elements(158);
    cp_elements(159) <= ptr_deref_1402_base_resize_ack_0;
    ptr_deref_1402_root_address_inst_req_0 <= cp_elements(159);
    cp_elements(160) <= ptr_deref_1402_root_address_inst_ack_0;
    ptr_deref_1402_addr_0_req_0 <= cp_elements(160);
    cp_elements(161) <= ptr_deref_1402_addr_0_ack_0;
    cp_elements(162) <= ptr_deref_1402_gather_scatter_ack_0;
    ptr_deref_1402_store_0_req_0 <= cp_elements(162);
    cp_elements(163) <= ptr_deref_1402_store_0_ack_0;
    cp_elements(164) <= cp_elements(163);
    ptr_deref_1402_store_0_req_1 <= cp_elements(164);
    cp_elements(165) <= ptr_deref_1402_store_0_ack_1;
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(167) & cp_elements(168));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1409_inst_req_0 <= cp_elements(166);
    cp_elements(167) <= cp_elements(129);
    cp_elements(168) <= cp_elements(129);
    cp_elements(169) <= binary_1409_inst_ack_0;
    binary_1409_inst_req_1 <= cp_elements(169);
    cp_elements(170) <= binary_1409_inst_ack_1;
    cpelement_group_171 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(170) & cp_elements(172));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(171),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1413_inst_req_0 <= cp_elements(171);
    cp_elements(172) <= cp_elements(129);
    cp_elements(173) <= type_cast_1413_inst_ack_0;
    cpelement_group_174 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(163) & cp_elements(173) & cp_elements(175) & cp_elements(179));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(174),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1416_gather_scatter_req_0 <= cp_elements(174);
    cp_elements(175) <= cp_elements(129);
    cp_elements(176) <= cp_elements(175);
    ptr_deref_1416_base_resize_req_0 <= cp_elements(176);
    cp_elements(177) <= ptr_deref_1416_base_resize_ack_0;
    ptr_deref_1416_root_address_inst_req_0 <= cp_elements(177);
    cp_elements(178) <= ptr_deref_1416_root_address_inst_ack_0;
    ptr_deref_1416_addr_0_req_0 <= cp_elements(178);
    cp_elements(179) <= ptr_deref_1416_addr_0_ack_0;
    cp_elements(180) <= ptr_deref_1416_gather_scatter_ack_0;
    ptr_deref_1416_store_0_req_0 <= cp_elements(180);
    cp_elements(181) <= ptr_deref_1416_store_0_ack_0;
    cp_elements(182) <= cp_elements(181);
    ptr_deref_1416_store_0_req_1 <= cp_elements(182);
    cp_elements(183) <= ptr_deref_1416_store_0_ack_1;
    cpelement_group_184 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(185) & cp_elements(186));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(184),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1423_inst_req_0 <= cp_elements(184);
    cp_elements(185) <= cp_elements(129);
    cp_elements(186) <= cp_elements(129);
    cp_elements(187) <= binary_1423_inst_ack_0;
    binary_1423_inst_req_1 <= cp_elements(187);
    cp_elements(188) <= binary_1423_inst_ack_1;
    cpelement_group_189 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(188) & cp_elements(190));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(189),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1427_inst_req_0 <= cp_elements(189);
    cp_elements(190) <= cp_elements(129);
    cp_elements(191) <= type_cast_1427_inst_ack_0;
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(191) & cp_elements(193) & cp_elements(197));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1430_gather_scatter_req_0 <= cp_elements(192);
    cp_elements(193) <= cp_elements(129);
    cp_elements(194) <= cp_elements(193);
    ptr_deref_1430_base_resize_req_0 <= cp_elements(194);
    cp_elements(195) <= ptr_deref_1430_base_resize_ack_0;
    ptr_deref_1430_root_address_inst_req_0 <= cp_elements(195);
    cp_elements(196) <= ptr_deref_1430_root_address_inst_ack_0;
    ptr_deref_1430_addr_0_req_0 <= cp_elements(196);
    cp_elements(197) <= ptr_deref_1430_addr_0_ack_0;
    cp_elements(198) <= ptr_deref_1430_gather_scatter_ack_0;
    ptr_deref_1430_store_0_req_0 <= cp_elements(198);
    cp_elements(199) <= ptr_deref_1430_store_0_ack_0;
    cp_elements(200) <= cp_elements(199);
    ptr_deref_1430_store_0_req_1 <= cp_elements(200);
    cp_elements(201) <= ptr_deref_1430_store_0_ack_1;
    cpelement_group_202 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(204));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(202),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1437_inst_req_0 <= cp_elements(202);
    cp_elements(203) <= cp_elements(129);
    cp_elements(204) <= cp_elements(129);
    cp_elements(205) <= binary_1437_inst_ack_0;
    binary_1437_inst_req_1 <= cp_elements(205);
    cp_elements(206) <= binary_1437_inst_ack_1;
    cpelement_group_207 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(206) & cp_elements(208));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(207),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1441_inst_req_0 <= cp_elements(207);
    cp_elements(208) <= cp_elements(129);
    cp_elements(209) <= type_cast_1441_inst_ack_0;
    cpelement_group_210 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(209) & cp_elements(211) & cp_elements(215));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(210),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1444_gather_scatter_req_0 <= cp_elements(210);
    cp_elements(211) <= cp_elements(129);
    cp_elements(212) <= cp_elements(211);
    ptr_deref_1444_base_resize_req_0 <= cp_elements(212);
    cp_elements(213) <= ptr_deref_1444_base_resize_ack_0;
    ptr_deref_1444_root_address_inst_req_0 <= cp_elements(213);
    cp_elements(214) <= ptr_deref_1444_root_address_inst_ack_0;
    ptr_deref_1444_addr_0_req_0 <= cp_elements(214);
    cp_elements(215) <= ptr_deref_1444_addr_0_ack_0;
    cp_elements(216) <= ptr_deref_1444_gather_scatter_ack_0;
    ptr_deref_1444_store_0_req_0 <= cp_elements(216);
    cp_elements(217) <= ptr_deref_1444_store_0_ack_0;
    cp_elements(218) <= cp_elements(217);
    ptr_deref_1444_store_0_req_1 <= cp_elements(218);
    cp_elements(219) <= ptr_deref_1444_store_0_ack_1;
    cpelement_group_220 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(221) & cp_elements(222));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(220),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1451_inst_req_0 <= cp_elements(220);
    cp_elements(221) <= cp_elements(129);
    cp_elements(222) <= cp_elements(129);
    cp_elements(223) <= binary_1451_inst_ack_0;
    binary_1451_inst_req_1 <= cp_elements(223);
    cp_elements(224) <= binary_1451_inst_ack_1;
    cpelement_group_225 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(224) & cp_elements(226));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(225),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1455_inst_req_0 <= cp_elements(225);
    cp_elements(226) <= cp_elements(129);
    cp_elements(227) <= type_cast_1455_inst_ack_0;
    cpelement_group_228 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(217) & cp_elements(227) & cp_elements(229) & cp_elements(233));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1458_gather_scatter_req_0 <= cp_elements(228);
    cp_elements(229) <= cp_elements(129);
    cp_elements(230) <= cp_elements(229);
    ptr_deref_1458_base_resize_req_0 <= cp_elements(230);
    cp_elements(231) <= ptr_deref_1458_base_resize_ack_0;
    ptr_deref_1458_root_address_inst_req_0 <= cp_elements(231);
    cp_elements(232) <= ptr_deref_1458_root_address_inst_ack_0;
    ptr_deref_1458_addr_0_req_0 <= cp_elements(232);
    cp_elements(233) <= ptr_deref_1458_addr_0_ack_0;
    cp_elements(234) <= ptr_deref_1458_gather_scatter_ack_0;
    ptr_deref_1458_store_0_req_0 <= cp_elements(234);
    cp_elements(235) <= ptr_deref_1458_store_0_ack_0;
    cp_elements(236) <= cp_elements(235);
    ptr_deref_1458_store_0_req_1 <= cp_elements(236);
    cp_elements(237) <= ptr_deref_1458_store_0_ack_1;
    cpelement_group_238 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(239) & cp_elements(240));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(238),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1465_inst_req_0 <= cp_elements(238);
    cp_elements(239) <= cp_elements(129);
    cp_elements(240) <= cp_elements(129);
    cp_elements(241) <= binary_1465_inst_ack_0;
    binary_1465_inst_req_1 <= cp_elements(241);
    cp_elements(242) <= binary_1465_inst_ack_1;
    cpelement_group_243 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(242) & cp_elements(244));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(243),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1469_inst_req_0 <= cp_elements(243);
    cp_elements(244) <= cp_elements(129);
    cp_elements(245) <= type_cast_1469_inst_ack_0;
    cpelement_group_246 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(235) & cp_elements(245) & cp_elements(247) & cp_elements(251));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(246),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1472_gather_scatter_req_0 <= cp_elements(246);
    cp_elements(247) <= cp_elements(129);
    cp_elements(248) <= cp_elements(247);
    ptr_deref_1472_base_resize_req_0 <= cp_elements(248);
    cp_elements(249) <= ptr_deref_1472_base_resize_ack_0;
    ptr_deref_1472_root_address_inst_req_0 <= cp_elements(249);
    cp_elements(250) <= ptr_deref_1472_root_address_inst_ack_0;
    ptr_deref_1472_addr_0_req_0 <= cp_elements(250);
    cp_elements(251) <= ptr_deref_1472_addr_0_ack_0;
    cp_elements(252) <= ptr_deref_1472_gather_scatter_ack_0;
    ptr_deref_1472_store_0_req_0 <= cp_elements(252);
    cp_elements(253) <= ptr_deref_1472_store_0_ack_0;
    cp_elements(254) <= cp_elements(253);
    ptr_deref_1472_store_0_req_1 <= cp_elements(254);
    cp_elements(255) <= ptr_deref_1472_store_0_ack_1;
    cpelement_group_256 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(257) & cp_elements(258));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(256),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1477_inst_req_0 <= cp_elements(256);
    cp_elements(257) <= cp_elements(129);
    cp_elements(258) <= cp_elements(129);
    cp_elements(259) <= type_cast_1477_inst_ack_0;
    cpelement_group_260 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(253) & cp_elements(259) & cp_elements(261) & cp_elements(265));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(260),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1480_gather_scatter_req_0 <= cp_elements(260);
    cp_elements(261) <= cp_elements(129);
    cp_elements(262) <= cp_elements(261);
    ptr_deref_1480_base_resize_req_0 <= cp_elements(262);
    cp_elements(263) <= ptr_deref_1480_base_resize_ack_0;
    ptr_deref_1480_root_address_inst_req_0 <= cp_elements(263);
    cp_elements(264) <= ptr_deref_1480_root_address_inst_ack_0;
    ptr_deref_1480_addr_0_req_0 <= cp_elements(264);
    cp_elements(265) <= ptr_deref_1480_addr_0_ack_0;
    cp_elements(266) <= ptr_deref_1480_gather_scatter_ack_0;
    ptr_deref_1480_store_0_req_0 <= cp_elements(266);
    cp_elements(267) <= ptr_deref_1480_store_0_ack_0;
    ptr_deref_1480_store_0_req_1 <= cp_elements(267);
    cp_elements(268) <= ptr_deref_1480_store_0_ack_1;
    cpelement_group_269 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(147) & cp_elements(165) & cp_elements(183) & cp_elements(201) & cp_elements(219) & cp_elements(237) & cp_elements(255) & cp_elements(268));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(269),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(270) <= cp_elements(126);
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(272) & cp_elements(273));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1489_inst_req_0 <= cp_elements(271);
    cp_elements(272) <= cp_elements(270);
    cp_elements(273) <= cp_elements(270);
    cp_elements(274) <= binary_1489_inst_ack_0;
    binary_1489_inst_req_1 <= cp_elements(274);
    cp_elements(275) <= binary_1489_inst_ack_1;
    array_obj_ref_1533_index_0_resize_req_0 <= cp_elements(275);
    cpelement_group_276 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(277) & cp_elements(278));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1495_inst_req_0 <= cp_elements(276);
    cp_elements(277) <= cp_elements(270);
    cp_elements(278) <= cp_elements(270);
    cp_elements(279) <= binary_1495_inst_ack_0;
    binary_1495_inst_req_1 <= cp_elements(279);
    cp_elements(280) <= binary_1495_inst_ack_1;
    array_obj_ref_1537_index_0_resize_req_0 <= cp_elements(280);
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(282) & cp_elements(283));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1501_inst_req_0 <= cp_elements(281);
    cp_elements(282) <= cp_elements(270);
    cp_elements(283) <= cp_elements(270);
    cp_elements(284) <= binary_1501_inst_ack_0;
    binary_1501_inst_req_1 <= cp_elements(284);
    cp_elements(285) <= binary_1501_inst_ack_1;
    array_obj_ref_1541_index_0_resize_req_0 <= cp_elements(285);
    cpelement_group_286 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(287) & cp_elements(288));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(286),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1507_inst_req_0 <= cp_elements(286);
    cp_elements(287) <= cp_elements(270);
    cp_elements(288) <= cp_elements(270);
    cp_elements(289) <= binary_1507_inst_ack_0;
    binary_1507_inst_req_1 <= cp_elements(289);
    cp_elements(290) <= binary_1507_inst_ack_1;
    array_obj_ref_1545_index_0_resize_req_0 <= cp_elements(290);
    cpelement_group_291 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(292) & cp_elements(293));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(291),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1513_inst_req_0 <= cp_elements(291);
    cp_elements(292) <= cp_elements(270);
    cp_elements(293) <= cp_elements(270);
    cp_elements(294) <= binary_1513_inst_ack_0;
    binary_1513_inst_req_1 <= cp_elements(294);
    cp_elements(295) <= binary_1513_inst_ack_1;
    array_obj_ref_1549_index_0_resize_req_0 <= cp_elements(295);
    cpelement_group_296 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(297) & cp_elements(298));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(296),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1519_inst_req_0 <= cp_elements(296);
    cp_elements(297) <= cp_elements(270);
    cp_elements(298) <= cp_elements(270);
    cp_elements(299) <= binary_1519_inst_ack_0;
    binary_1519_inst_req_1 <= cp_elements(299);
    cp_elements(300) <= binary_1519_inst_ack_1;
    array_obj_ref_1553_index_0_resize_req_0 <= cp_elements(300);
    cpelement_group_301 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(302) & cp_elements(303));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(301),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1525_inst_req_0 <= cp_elements(301);
    cp_elements(302) <= cp_elements(270);
    cp_elements(303) <= cp_elements(270);
    cp_elements(304) <= binary_1525_inst_ack_0;
    binary_1525_inst_req_1 <= cp_elements(304);
    cp_elements(305) <= binary_1525_inst_ack_1;
    array_obj_ref_1557_index_0_resize_req_0 <= cp_elements(305);
    cp_elements(306) <= cp_elements(270);
    cpelement_group_307 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(306) & cp_elements(316));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(307),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1529_final_reg_req_0 <= cp_elements(307);
    cp_elements(308) <= cp_elements(270);
    array_obj_ref_1529_base_resize_req_0 <= cp_elements(308);
    cp_elements(309) <= cp_elements(270);
    array_obj_ref_1529_index_0_resize_req_0 <= cp_elements(309);
    cp_elements(310) <= array_obj_ref_1529_index_0_resize_ack_0;
    array_obj_ref_1529_index_0_rename_req_0 <= cp_elements(310);
    cp_elements(311) <= array_obj_ref_1529_index_0_rename_ack_0;
    array_obj_ref_1529_offset_inst_req_0 <= cp_elements(311);
    cp_elements(312) <= array_obj_ref_1529_offset_inst_ack_0;
    cp_elements(313) <= array_obj_ref_1529_base_resize_ack_0;
    cpelement_group_314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(312) & cp_elements(313));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1529_root_address_inst_req_0 <= cp_elements(314);
    cp_elements(315) <= array_obj_ref_1529_root_address_inst_ack_0;
    array_obj_ref_1529_root_address_inst_req_1 <= cp_elements(315);
    cp_elements(316) <= array_obj_ref_1529_root_address_inst_ack_1;
    cp_elements(317) <= array_obj_ref_1529_final_reg_ack_0;
    cp_elements(318) <= cp_elements(270);
    cpelement_group_319 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(318) & cp_elements(327));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(319),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1533_final_reg_req_0 <= cp_elements(319);
    cp_elements(320) <= cp_elements(270);
    array_obj_ref_1533_base_resize_req_0 <= cp_elements(320);
    cp_elements(321) <= array_obj_ref_1533_index_0_resize_ack_0;
    array_obj_ref_1533_index_0_rename_req_0 <= cp_elements(321);
    cp_elements(322) <= array_obj_ref_1533_index_0_rename_ack_0;
    array_obj_ref_1533_offset_inst_req_0 <= cp_elements(322);
    cp_elements(323) <= array_obj_ref_1533_offset_inst_ack_0;
    cp_elements(324) <= array_obj_ref_1533_base_resize_ack_0;
    cpelement_group_325 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(323) & cp_elements(324));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(325),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1533_root_address_inst_req_0 <= cp_elements(325);
    cp_elements(326) <= array_obj_ref_1533_root_address_inst_ack_0;
    array_obj_ref_1533_root_address_inst_req_1 <= cp_elements(326);
    cp_elements(327) <= array_obj_ref_1533_root_address_inst_ack_1;
    cp_elements(328) <= array_obj_ref_1533_final_reg_ack_0;
    cp_elements(329) <= cp_elements(270);
    cpelement_group_330 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(338));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(330),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1537_final_reg_req_0 <= cp_elements(330);
    cp_elements(331) <= cp_elements(270);
    array_obj_ref_1537_base_resize_req_0 <= cp_elements(331);
    cp_elements(332) <= array_obj_ref_1537_index_0_resize_ack_0;
    array_obj_ref_1537_index_0_rename_req_0 <= cp_elements(332);
    cp_elements(333) <= array_obj_ref_1537_index_0_rename_ack_0;
    array_obj_ref_1537_offset_inst_req_0 <= cp_elements(333);
    cp_elements(334) <= array_obj_ref_1537_offset_inst_ack_0;
    cp_elements(335) <= array_obj_ref_1537_base_resize_ack_0;
    cpelement_group_336 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(334) & cp_elements(335));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(336),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1537_root_address_inst_req_0 <= cp_elements(336);
    cp_elements(337) <= array_obj_ref_1537_root_address_inst_ack_0;
    array_obj_ref_1537_root_address_inst_req_1 <= cp_elements(337);
    cp_elements(338) <= array_obj_ref_1537_root_address_inst_ack_1;
    cp_elements(339) <= array_obj_ref_1537_final_reg_ack_0;
    cp_elements(340) <= cp_elements(270);
    cpelement_group_341 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(340) & cp_elements(349));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1541_final_reg_req_0 <= cp_elements(341);
    cp_elements(342) <= cp_elements(270);
    array_obj_ref_1541_base_resize_req_0 <= cp_elements(342);
    cp_elements(343) <= array_obj_ref_1541_index_0_resize_ack_0;
    array_obj_ref_1541_index_0_rename_req_0 <= cp_elements(343);
    cp_elements(344) <= array_obj_ref_1541_index_0_rename_ack_0;
    array_obj_ref_1541_offset_inst_req_0 <= cp_elements(344);
    cp_elements(345) <= array_obj_ref_1541_offset_inst_ack_0;
    cp_elements(346) <= array_obj_ref_1541_base_resize_ack_0;
    cpelement_group_347 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(345) & cp_elements(346));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(347),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1541_root_address_inst_req_0 <= cp_elements(347);
    cp_elements(348) <= array_obj_ref_1541_root_address_inst_ack_0;
    array_obj_ref_1541_root_address_inst_req_1 <= cp_elements(348);
    cp_elements(349) <= array_obj_ref_1541_root_address_inst_ack_1;
    cp_elements(350) <= array_obj_ref_1541_final_reg_ack_0;
    cp_elements(351) <= cp_elements(270);
    cpelement_group_352 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(351) & cp_elements(360));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(352),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1545_final_reg_req_0 <= cp_elements(352);
    cp_elements(353) <= cp_elements(270);
    array_obj_ref_1545_base_resize_req_0 <= cp_elements(353);
    cp_elements(354) <= array_obj_ref_1545_index_0_resize_ack_0;
    array_obj_ref_1545_index_0_rename_req_0 <= cp_elements(354);
    cp_elements(355) <= array_obj_ref_1545_index_0_rename_ack_0;
    array_obj_ref_1545_offset_inst_req_0 <= cp_elements(355);
    cp_elements(356) <= array_obj_ref_1545_offset_inst_ack_0;
    cp_elements(357) <= array_obj_ref_1545_base_resize_ack_0;
    cpelement_group_358 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(356) & cp_elements(357));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(358),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1545_root_address_inst_req_0 <= cp_elements(358);
    cp_elements(359) <= array_obj_ref_1545_root_address_inst_ack_0;
    array_obj_ref_1545_root_address_inst_req_1 <= cp_elements(359);
    cp_elements(360) <= array_obj_ref_1545_root_address_inst_ack_1;
    cp_elements(361) <= array_obj_ref_1545_final_reg_ack_0;
    cp_elements(362) <= cp_elements(270);
    cpelement_group_363 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(362) & cp_elements(371));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1549_final_reg_req_0 <= cp_elements(363);
    cp_elements(364) <= cp_elements(270);
    array_obj_ref_1549_base_resize_req_0 <= cp_elements(364);
    cp_elements(365) <= array_obj_ref_1549_index_0_resize_ack_0;
    array_obj_ref_1549_index_0_rename_req_0 <= cp_elements(365);
    cp_elements(366) <= array_obj_ref_1549_index_0_rename_ack_0;
    array_obj_ref_1549_offset_inst_req_0 <= cp_elements(366);
    cp_elements(367) <= array_obj_ref_1549_offset_inst_ack_0;
    cp_elements(368) <= array_obj_ref_1549_base_resize_ack_0;
    cpelement_group_369 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(367) & cp_elements(368));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(369),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1549_root_address_inst_req_0 <= cp_elements(369);
    cp_elements(370) <= array_obj_ref_1549_root_address_inst_ack_0;
    array_obj_ref_1549_root_address_inst_req_1 <= cp_elements(370);
    cp_elements(371) <= array_obj_ref_1549_root_address_inst_ack_1;
    cp_elements(372) <= array_obj_ref_1549_final_reg_ack_0;
    cp_elements(373) <= cp_elements(270);
    cpelement_group_374 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(373) & cp_elements(382));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1553_final_reg_req_0 <= cp_elements(374);
    cp_elements(375) <= cp_elements(270);
    array_obj_ref_1553_base_resize_req_0 <= cp_elements(375);
    cp_elements(376) <= array_obj_ref_1553_index_0_resize_ack_0;
    array_obj_ref_1553_index_0_rename_req_0 <= cp_elements(376);
    cp_elements(377) <= array_obj_ref_1553_index_0_rename_ack_0;
    array_obj_ref_1553_offset_inst_req_0 <= cp_elements(377);
    cp_elements(378) <= array_obj_ref_1553_offset_inst_ack_0;
    cp_elements(379) <= array_obj_ref_1553_base_resize_ack_0;
    cpelement_group_380 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(378) & cp_elements(379));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(380),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1553_root_address_inst_req_0 <= cp_elements(380);
    cp_elements(381) <= array_obj_ref_1553_root_address_inst_ack_0;
    array_obj_ref_1553_root_address_inst_req_1 <= cp_elements(381);
    cp_elements(382) <= array_obj_ref_1553_root_address_inst_ack_1;
    cp_elements(383) <= array_obj_ref_1553_final_reg_ack_0;
    cp_elements(384) <= cp_elements(270);
    cpelement_group_385 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(384) & cp_elements(393));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(385),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1557_final_reg_req_0 <= cp_elements(385);
    cp_elements(386) <= cp_elements(270);
    array_obj_ref_1557_base_resize_req_0 <= cp_elements(386);
    cp_elements(387) <= array_obj_ref_1557_index_0_resize_ack_0;
    array_obj_ref_1557_index_0_rename_req_0 <= cp_elements(387);
    cp_elements(388) <= array_obj_ref_1557_index_0_rename_ack_0;
    array_obj_ref_1557_offset_inst_req_0 <= cp_elements(388);
    cp_elements(389) <= array_obj_ref_1557_offset_inst_ack_0;
    cp_elements(390) <= array_obj_ref_1557_base_resize_ack_0;
    cpelement_group_391 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(389) & cp_elements(390));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(391),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1557_root_address_inst_req_0 <= cp_elements(391);
    cp_elements(392) <= array_obj_ref_1557_root_address_inst_ack_0;
    array_obj_ref_1557_root_address_inst_req_1 <= cp_elements(392);
    cp_elements(393) <= array_obj_ref_1557_root_address_inst_ack_1;
    cp_elements(394) <= array_obj_ref_1557_final_reg_ack_0;
    cpelement_group_395 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(396) & cp_elements(397));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(395),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1563_inst_req_0 <= cp_elements(395);
    cp_elements(396) <= cp_elements(270);
    cp_elements(397) <= cp_elements(270);
    cp_elements(398) <= binary_1563_inst_ack_0;
    binary_1563_inst_req_1 <= cp_elements(398);
    cp_elements(399) <= binary_1563_inst_ack_1;
    cpelement_group_400 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(399) & cp_elements(401));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(400),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1567_inst_req_0 <= cp_elements(400);
    cp_elements(401) <= cp_elements(270);
    cp_elements(402) <= type_cast_1567_inst_ack_0;
    cpelement_group_403 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(317) & cp_elements(402) & cp_elements(407));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(403),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1570_gather_scatter_req_0 <= cp_elements(403);
    cp_elements(404) <= cp_elements(317);
    ptr_deref_1570_base_resize_req_0 <= cp_elements(404);
    cp_elements(405) <= ptr_deref_1570_base_resize_ack_0;
    ptr_deref_1570_root_address_inst_req_0 <= cp_elements(405);
    cp_elements(406) <= ptr_deref_1570_root_address_inst_ack_0;
    ptr_deref_1570_addr_0_req_0 <= cp_elements(406);
    cp_elements(407) <= ptr_deref_1570_addr_0_ack_0;
    cp_elements(408) <= ptr_deref_1570_gather_scatter_ack_0;
    ptr_deref_1570_store_0_req_0 <= cp_elements(408);
    cp_elements(409) <= ptr_deref_1570_store_0_ack_0;
    cp_elements(410) <= cp_elements(409);
    ptr_deref_1570_store_0_req_1 <= cp_elements(410);
    cp_elements(411) <= ptr_deref_1570_store_0_ack_1;
    cpelement_group_412 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(413) & cp_elements(414));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(412),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1577_inst_req_0 <= cp_elements(412);
    cp_elements(413) <= cp_elements(270);
    cp_elements(414) <= cp_elements(270);
    cp_elements(415) <= binary_1577_inst_ack_0;
    binary_1577_inst_req_1 <= cp_elements(415);
    cp_elements(416) <= binary_1577_inst_ack_1;
    cpelement_group_417 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(416) & cp_elements(418));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(417),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1581_inst_req_0 <= cp_elements(417);
    cp_elements(418) <= cp_elements(270);
    cp_elements(419) <= type_cast_1581_inst_ack_0;
    cpelement_group_420 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(328) & cp_elements(409) & cp_elements(419) & cp_elements(424));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(420),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1584_gather_scatter_req_0 <= cp_elements(420);
    cp_elements(421) <= cp_elements(328);
    ptr_deref_1584_base_resize_req_0 <= cp_elements(421);
    cp_elements(422) <= ptr_deref_1584_base_resize_ack_0;
    ptr_deref_1584_root_address_inst_req_0 <= cp_elements(422);
    cp_elements(423) <= ptr_deref_1584_root_address_inst_ack_0;
    ptr_deref_1584_addr_0_req_0 <= cp_elements(423);
    cp_elements(424) <= ptr_deref_1584_addr_0_ack_0;
    cp_elements(425) <= ptr_deref_1584_gather_scatter_ack_0;
    ptr_deref_1584_store_0_req_0 <= cp_elements(425);
    cp_elements(426) <= ptr_deref_1584_store_0_ack_0;
    cp_elements(427) <= cp_elements(426);
    ptr_deref_1584_store_0_req_1 <= cp_elements(427);
    cp_elements(428) <= ptr_deref_1584_store_0_ack_1;
    cpelement_group_429 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(430) & cp_elements(431));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(429),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1591_inst_req_0 <= cp_elements(429);
    cp_elements(430) <= cp_elements(270);
    cp_elements(431) <= cp_elements(270);
    cp_elements(432) <= binary_1591_inst_ack_0;
    binary_1591_inst_req_1 <= cp_elements(432);
    cp_elements(433) <= binary_1591_inst_ack_1;
    cpelement_group_434 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(433) & cp_elements(435));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(434),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1595_inst_req_0 <= cp_elements(434);
    cp_elements(435) <= cp_elements(270);
    cp_elements(436) <= type_cast_1595_inst_ack_0;
    cpelement_group_437 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(339) & cp_elements(426) & cp_elements(436) & cp_elements(441));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(437),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1598_gather_scatter_req_0 <= cp_elements(437);
    cp_elements(438) <= cp_elements(339);
    ptr_deref_1598_base_resize_req_0 <= cp_elements(438);
    cp_elements(439) <= ptr_deref_1598_base_resize_ack_0;
    ptr_deref_1598_root_address_inst_req_0 <= cp_elements(439);
    cp_elements(440) <= ptr_deref_1598_root_address_inst_ack_0;
    ptr_deref_1598_addr_0_req_0 <= cp_elements(440);
    cp_elements(441) <= ptr_deref_1598_addr_0_ack_0;
    cp_elements(442) <= ptr_deref_1598_gather_scatter_ack_0;
    ptr_deref_1598_store_0_req_0 <= cp_elements(442);
    cp_elements(443) <= ptr_deref_1598_store_0_ack_0;
    cp_elements(444) <= cp_elements(443);
    ptr_deref_1598_store_0_req_1 <= cp_elements(444);
    cp_elements(445) <= ptr_deref_1598_store_0_ack_1;
    cpelement_group_446 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(447) & cp_elements(448));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(446),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1605_inst_req_0 <= cp_elements(446);
    cp_elements(447) <= cp_elements(270);
    cp_elements(448) <= cp_elements(270);
    cp_elements(449) <= binary_1605_inst_ack_0;
    binary_1605_inst_req_1 <= cp_elements(449);
    cp_elements(450) <= binary_1605_inst_ack_1;
    cpelement_group_451 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(450) & cp_elements(452));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(451),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1609_inst_req_0 <= cp_elements(451);
    cp_elements(452) <= cp_elements(270);
    cp_elements(453) <= type_cast_1609_inst_ack_0;
    cpelement_group_454 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(350) & cp_elements(443) & cp_elements(453) & cp_elements(458));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(454),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1612_gather_scatter_req_0 <= cp_elements(454);
    cp_elements(455) <= cp_elements(350);
    ptr_deref_1612_base_resize_req_0 <= cp_elements(455);
    cp_elements(456) <= ptr_deref_1612_base_resize_ack_0;
    ptr_deref_1612_root_address_inst_req_0 <= cp_elements(456);
    cp_elements(457) <= ptr_deref_1612_root_address_inst_ack_0;
    ptr_deref_1612_addr_0_req_0 <= cp_elements(457);
    cp_elements(458) <= ptr_deref_1612_addr_0_ack_0;
    cp_elements(459) <= ptr_deref_1612_gather_scatter_ack_0;
    ptr_deref_1612_store_0_req_0 <= cp_elements(459);
    cp_elements(460) <= ptr_deref_1612_store_0_ack_0;
    cp_elements(461) <= cp_elements(460);
    ptr_deref_1612_store_0_req_1 <= cp_elements(461);
    cp_elements(462) <= ptr_deref_1612_store_0_ack_1;
    cpelement_group_463 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(464) & cp_elements(465));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(463),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1619_inst_req_0 <= cp_elements(463);
    cp_elements(464) <= cp_elements(270);
    cp_elements(465) <= cp_elements(270);
    cp_elements(466) <= binary_1619_inst_ack_0;
    binary_1619_inst_req_1 <= cp_elements(466);
    cp_elements(467) <= binary_1619_inst_ack_1;
    cpelement_group_468 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(467) & cp_elements(469));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(468),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1623_inst_req_0 <= cp_elements(468);
    cp_elements(469) <= cp_elements(270);
    cp_elements(470) <= type_cast_1623_inst_ack_0;
    cpelement_group_471 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(460) & cp_elements(470) & cp_elements(475));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(471),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1626_gather_scatter_req_0 <= cp_elements(471);
    cp_elements(472) <= cp_elements(361);
    ptr_deref_1626_base_resize_req_0 <= cp_elements(472);
    cp_elements(473) <= ptr_deref_1626_base_resize_ack_0;
    ptr_deref_1626_root_address_inst_req_0 <= cp_elements(473);
    cp_elements(474) <= ptr_deref_1626_root_address_inst_ack_0;
    ptr_deref_1626_addr_0_req_0 <= cp_elements(474);
    cp_elements(475) <= ptr_deref_1626_addr_0_ack_0;
    cp_elements(476) <= ptr_deref_1626_gather_scatter_ack_0;
    ptr_deref_1626_store_0_req_0 <= cp_elements(476);
    cp_elements(477) <= ptr_deref_1626_store_0_ack_0;
    cp_elements(478) <= cp_elements(477);
    ptr_deref_1626_store_0_req_1 <= cp_elements(478);
    cp_elements(479) <= ptr_deref_1626_store_0_ack_1;
    cpelement_group_480 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(481) & cp_elements(482));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(480),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1633_inst_req_0 <= cp_elements(480);
    cp_elements(481) <= cp_elements(270);
    cp_elements(482) <= cp_elements(270);
    cp_elements(483) <= binary_1633_inst_ack_0;
    binary_1633_inst_req_1 <= cp_elements(483);
    cp_elements(484) <= binary_1633_inst_ack_1;
    cpelement_group_485 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(484) & cp_elements(486));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(485),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1637_inst_req_0 <= cp_elements(485);
    cp_elements(486) <= cp_elements(270);
    cp_elements(487) <= type_cast_1637_inst_ack_0;
    cpelement_group_488 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(372) & cp_elements(477) & cp_elements(487) & cp_elements(492));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(488),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1640_gather_scatter_req_0 <= cp_elements(488);
    cp_elements(489) <= cp_elements(372);
    ptr_deref_1640_base_resize_req_0 <= cp_elements(489);
    cp_elements(490) <= ptr_deref_1640_base_resize_ack_0;
    ptr_deref_1640_root_address_inst_req_0 <= cp_elements(490);
    cp_elements(491) <= ptr_deref_1640_root_address_inst_ack_0;
    ptr_deref_1640_addr_0_req_0 <= cp_elements(491);
    cp_elements(492) <= ptr_deref_1640_addr_0_ack_0;
    cp_elements(493) <= ptr_deref_1640_gather_scatter_ack_0;
    ptr_deref_1640_store_0_req_0 <= cp_elements(493);
    cp_elements(494) <= ptr_deref_1640_store_0_ack_0;
    cp_elements(495) <= cp_elements(494);
    ptr_deref_1640_store_0_req_1 <= cp_elements(495);
    cp_elements(496) <= ptr_deref_1640_store_0_ack_1;
    cpelement_group_497 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(498) & cp_elements(499));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(497),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1647_inst_req_0 <= cp_elements(497);
    cp_elements(498) <= cp_elements(270);
    cp_elements(499) <= cp_elements(270);
    cp_elements(500) <= binary_1647_inst_ack_0;
    binary_1647_inst_req_1 <= cp_elements(500);
    cp_elements(501) <= binary_1647_inst_ack_1;
    cpelement_group_502 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(501) & cp_elements(503));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(502),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1651_inst_req_0 <= cp_elements(502);
    cp_elements(503) <= cp_elements(270);
    cp_elements(504) <= type_cast_1651_inst_ack_0;
    cpelement_group_505 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(383) & cp_elements(494) & cp_elements(504) & cp_elements(509));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(505),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1654_gather_scatter_req_0 <= cp_elements(505);
    cp_elements(506) <= cp_elements(383);
    ptr_deref_1654_base_resize_req_0 <= cp_elements(506);
    cp_elements(507) <= ptr_deref_1654_base_resize_ack_0;
    ptr_deref_1654_root_address_inst_req_0 <= cp_elements(507);
    cp_elements(508) <= ptr_deref_1654_root_address_inst_ack_0;
    ptr_deref_1654_addr_0_req_0 <= cp_elements(508);
    cp_elements(509) <= ptr_deref_1654_addr_0_ack_0;
    cp_elements(510) <= ptr_deref_1654_gather_scatter_ack_0;
    ptr_deref_1654_store_0_req_0 <= cp_elements(510);
    cp_elements(511) <= ptr_deref_1654_store_0_ack_0;
    cp_elements(512) <= cp_elements(511);
    ptr_deref_1654_store_0_req_1 <= cp_elements(512);
    cp_elements(513) <= ptr_deref_1654_store_0_ack_1;
    cpelement_group_514 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(515) & cp_elements(516));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(514),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1659_inst_req_0 <= cp_elements(514);
    cp_elements(515) <= cp_elements(270);
    cp_elements(516) <= cp_elements(270);
    cp_elements(517) <= type_cast_1659_inst_ack_0;
    cpelement_group_518 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(394) & cp_elements(511) & cp_elements(517) & cp_elements(522));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1662_gather_scatter_req_0 <= cp_elements(518);
    cp_elements(519) <= cp_elements(394);
    ptr_deref_1662_base_resize_req_0 <= cp_elements(519);
    cp_elements(520) <= ptr_deref_1662_base_resize_ack_0;
    ptr_deref_1662_root_address_inst_req_0 <= cp_elements(520);
    cp_elements(521) <= ptr_deref_1662_root_address_inst_ack_0;
    ptr_deref_1662_addr_0_req_0 <= cp_elements(521);
    cp_elements(522) <= ptr_deref_1662_addr_0_ack_0;
    cp_elements(523) <= ptr_deref_1662_gather_scatter_ack_0;
    ptr_deref_1662_store_0_req_0 <= cp_elements(523);
    cp_elements(524) <= ptr_deref_1662_store_0_ack_0;
    ptr_deref_1662_store_0_req_1 <= cp_elements(524);
    cp_elements(525) <= ptr_deref_1662_store_0_ack_1;
    cpelement_group_526 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(411) & cp_elements(428) & cp_elements(445) & cp_elements(462) & cp_elements(479) & cp_elements(496) & cp_elements(513) & cp_elements(525));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(526),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(527) <= cp_elements(809);
    cpelement_group_528 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(529) & cp_elements(530));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(528),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1671_inst_req_0 <= cp_elements(528);
    cp_elements(529) <= cp_elements(527);
    cp_elements(530) <= cp_elements(527);
    cp_elements(531) <= binary_1671_inst_ack_0;
    binary_1671_inst_req_1 <= cp_elements(531);
    cp_elements(532) <= binary_1671_inst_ack_1;
    type_cast_1336_inst_req_0 <= cp_elements(532);
    cp_elements(533) <= cp_elements(128);
    cpelement_group_534 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(535) & cp_elements(536));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(534),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1679_inst_req_0 <= cp_elements(534);
    cp_elements(535) <= cp_elements(533);
    cp_elements(536) <= cp_elements(533);
    cp_elements(537) <= binary_1679_inst_ack_0;
    binary_1679_inst_req_1 <= cp_elements(537);
    cp_elements(538) <= binary_1679_inst_ack_1;
    cpelement_group_539 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(538) & cp_elements(540));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(539),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1683_inst_req_0 <= cp_elements(539);
    cp_elements(540) <= cp_elements(533);
    cp_elements(541) <= type_cast_1683_inst_ack_0;
    cp_elements(542) <= cp_elements(533);
    cpelement_group_543 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(542) & cp_elements(552));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(543),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1687_final_reg_req_0 <= cp_elements(543);
    cp_elements(544) <= cp_elements(533);
    array_obj_ref_1687_base_resize_req_0 <= cp_elements(544);
    cp_elements(545) <= cp_elements(533);
    array_obj_ref_1687_index_0_resize_req_0 <= cp_elements(545);
    cp_elements(546) <= array_obj_ref_1687_index_0_resize_ack_0;
    array_obj_ref_1687_index_0_rename_req_0 <= cp_elements(546);
    cp_elements(547) <= array_obj_ref_1687_index_0_rename_ack_0;
    array_obj_ref_1687_offset_inst_req_0 <= cp_elements(547);
    cp_elements(548) <= array_obj_ref_1687_offset_inst_ack_0;
    cp_elements(549) <= array_obj_ref_1687_base_resize_ack_0;
    cpelement_group_550 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(548) & cp_elements(549));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(550),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1687_root_address_inst_req_0 <= cp_elements(550);
    cp_elements(551) <= array_obj_ref_1687_root_address_inst_ack_0;
    array_obj_ref_1687_root_address_inst_req_1 <= cp_elements(551);
    cp_elements(552) <= array_obj_ref_1687_root_address_inst_ack_1;
    cp_elements(553) <= array_obj_ref_1687_final_reg_ack_0;
    cpelement_group_554 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(541) & cp_elements(553) & cp_elements(558));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(554),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1690_gather_scatter_req_0 <= cp_elements(554);
    cp_elements(555) <= cp_elements(553);
    ptr_deref_1690_base_resize_req_0 <= cp_elements(555);
    cp_elements(556) <= ptr_deref_1690_base_resize_ack_0;
    ptr_deref_1690_root_address_inst_req_0 <= cp_elements(556);
    cp_elements(557) <= ptr_deref_1690_root_address_inst_ack_0;
    ptr_deref_1690_addr_0_req_0 <= cp_elements(557);
    cp_elements(558) <= ptr_deref_1690_addr_0_ack_0;
    cp_elements(559) <= ptr_deref_1690_gather_scatter_ack_0;
    ptr_deref_1690_store_0_req_0 <= cp_elements(559);
    cp_elements(560) <= ptr_deref_1690_store_0_ack_0;
    cp_elements(561) <= cp_elements(560);
    ptr_deref_1690_store_0_req_1 <= cp_elements(561);
    cp_elements(562) <= ptr_deref_1690_store_0_ack_1;
    cpelement_group_563 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(564) & cp_elements(565));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(563),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1697_inst_req_0 <= cp_elements(563);
    cp_elements(564) <= cp_elements(533);
    cp_elements(565) <= cp_elements(533);
    cp_elements(566) <= binary_1697_inst_ack_0;
    binary_1697_inst_req_1 <= cp_elements(566);
    cp_elements(567) <= binary_1697_inst_ack_1;
    cpelement_group_568 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(567) & cp_elements(569));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(568),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1701_inst_req_0 <= cp_elements(568);
    cp_elements(569) <= cp_elements(533);
    cp_elements(570) <= type_cast_1701_inst_ack_0;
    cpelement_group_571 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(572) & cp_elements(573));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(571),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1707_inst_req_0 <= cp_elements(571);
    cp_elements(572) <= cp_elements(533);
    cp_elements(573) <= cp_elements(533);
    cp_elements(574) <= binary_1707_inst_ack_0;
    binary_1707_inst_req_1 <= cp_elements(574);
    cp_elements(575) <= binary_1707_inst_ack_1;
    array_obj_ref_1711_index_0_resize_req_0 <= cp_elements(575);
    cp_elements(576) <= cp_elements(533);
    cpelement_group_577 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(576) & cp_elements(585));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(577),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1711_final_reg_req_0 <= cp_elements(577);
    cp_elements(578) <= cp_elements(533);
    array_obj_ref_1711_base_resize_req_0 <= cp_elements(578);
    cp_elements(579) <= array_obj_ref_1711_index_0_resize_ack_0;
    array_obj_ref_1711_index_0_rename_req_0 <= cp_elements(579);
    cp_elements(580) <= array_obj_ref_1711_index_0_rename_ack_0;
    array_obj_ref_1711_offset_inst_req_0 <= cp_elements(580);
    cp_elements(581) <= array_obj_ref_1711_offset_inst_ack_0;
    cp_elements(582) <= array_obj_ref_1711_base_resize_ack_0;
    cpelement_group_583 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(581) & cp_elements(582));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(583),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1711_root_address_inst_req_0 <= cp_elements(583);
    cp_elements(584) <= array_obj_ref_1711_root_address_inst_ack_0;
    array_obj_ref_1711_root_address_inst_req_1 <= cp_elements(584);
    cp_elements(585) <= array_obj_ref_1711_root_address_inst_ack_1;
    cp_elements(586) <= array_obj_ref_1711_final_reg_ack_0;
    cpelement_group_587 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(560) & cp_elements(570) & cp_elements(586) & cp_elements(591));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(587),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1714_gather_scatter_req_0 <= cp_elements(587);
    cp_elements(588) <= cp_elements(586);
    ptr_deref_1714_base_resize_req_0 <= cp_elements(588);
    cp_elements(589) <= ptr_deref_1714_base_resize_ack_0;
    ptr_deref_1714_root_address_inst_req_0 <= cp_elements(589);
    cp_elements(590) <= ptr_deref_1714_root_address_inst_ack_0;
    ptr_deref_1714_addr_0_req_0 <= cp_elements(590);
    cp_elements(591) <= ptr_deref_1714_addr_0_ack_0;
    cp_elements(592) <= ptr_deref_1714_gather_scatter_ack_0;
    ptr_deref_1714_store_0_req_0 <= cp_elements(592);
    cp_elements(593) <= ptr_deref_1714_store_0_ack_0;
    cp_elements(594) <= cp_elements(593);
    ptr_deref_1714_store_0_req_1 <= cp_elements(594);
    cp_elements(595) <= ptr_deref_1714_store_0_ack_1;
    cpelement_group_596 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(597) & cp_elements(598));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(596),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1721_inst_req_0 <= cp_elements(596);
    cp_elements(597) <= cp_elements(533);
    cp_elements(598) <= cp_elements(533);
    cp_elements(599) <= binary_1721_inst_ack_0;
    binary_1721_inst_req_1 <= cp_elements(599);
    cp_elements(600) <= binary_1721_inst_ack_1;
    cpelement_group_601 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(600) & cp_elements(602));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(601),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1725_inst_req_0 <= cp_elements(601);
    cp_elements(602) <= cp_elements(533);
    cp_elements(603) <= type_cast_1725_inst_ack_0;
    cpelement_group_604 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(605) & cp_elements(606));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(604),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1731_inst_req_0 <= cp_elements(604);
    cp_elements(605) <= cp_elements(533);
    cp_elements(606) <= cp_elements(533);
    cp_elements(607) <= binary_1731_inst_ack_0;
    binary_1731_inst_req_1 <= cp_elements(607);
    cp_elements(608) <= binary_1731_inst_ack_1;
    array_obj_ref_1735_index_0_resize_req_0 <= cp_elements(608);
    cp_elements(609) <= cp_elements(533);
    cpelement_group_610 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(609) & cp_elements(618));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(610),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1735_final_reg_req_0 <= cp_elements(610);
    cp_elements(611) <= cp_elements(533);
    array_obj_ref_1735_base_resize_req_0 <= cp_elements(611);
    cp_elements(612) <= array_obj_ref_1735_index_0_resize_ack_0;
    array_obj_ref_1735_index_0_rename_req_0 <= cp_elements(612);
    cp_elements(613) <= array_obj_ref_1735_index_0_rename_ack_0;
    array_obj_ref_1735_offset_inst_req_0 <= cp_elements(613);
    cp_elements(614) <= array_obj_ref_1735_offset_inst_ack_0;
    cp_elements(615) <= array_obj_ref_1735_base_resize_ack_0;
    cpelement_group_616 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(614) & cp_elements(615));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(616),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1735_root_address_inst_req_0 <= cp_elements(616);
    cp_elements(617) <= array_obj_ref_1735_root_address_inst_ack_0;
    array_obj_ref_1735_root_address_inst_req_1 <= cp_elements(617);
    cp_elements(618) <= array_obj_ref_1735_root_address_inst_ack_1;
    cp_elements(619) <= array_obj_ref_1735_final_reg_ack_0;
    cpelement_group_620 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(593) & cp_elements(603) & cp_elements(619) & cp_elements(624));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(620),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1738_gather_scatter_req_0 <= cp_elements(620);
    cp_elements(621) <= cp_elements(619);
    ptr_deref_1738_base_resize_req_0 <= cp_elements(621);
    cp_elements(622) <= ptr_deref_1738_base_resize_ack_0;
    ptr_deref_1738_root_address_inst_req_0 <= cp_elements(622);
    cp_elements(623) <= ptr_deref_1738_root_address_inst_ack_0;
    ptr_deref_1738_addr_0_req_0 <= cp_elements(623);
    cp_elements(624) <= ptr_deref_1738_addr_0_ack_0;
    cp_elements(625) <= ptr_deref_1738_gather_scatter_ack_0;
    ptr_deref_1738_store_0_req_0 <= cp_elements(625);
    cp_elements(626) <= ptr_deref_1738_store_0_ack_0;
    cp_elements(627) <= cp_elements(626);
    ptr_deref_1738_store_0_req_1 <= cp_elements(627);
    cp_elements(628) <= ptr_deref_1738_store_0_ack_1;
    cpelement_group_629 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(630) & cp_elements(631));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(629),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1745_inst_req_0 <= cp_elements(629);
    cp_elements(630) <= cp_elements(533);
    cp_elements(631) <= cp_elements(533);
    cp_elements(632) <= binary_1745_inst_ack_0;
    binary_1745_inst_req_1 <= cp_elements(632);
    cp_elements(633) <= binary_1745_inst_ack_1;
    cpelement_group_634 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(633) & cp_elements(635));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(634),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1749_inst_req_0 <= cp_elements(634);
    cp_elements(635) <= cp_elements(533);
    cp_elements(636) <= type_cast_1749_inst_ack_0;
    cpelement_group_637 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(638) & cp_elements(639));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(637),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1755_inst_req_0 <= cp_elements(637);
    cp_elements(638) <= cp_elements(533);
    cp_elements(639) <= cp_elements(533);
    cp_elements(640) <= binary_1755_inst_ack_0;
    binary_1755_inst_req_1 <= cp_elements(640);
    cp_elements(641) <= binary_1755_inst_ack_1;
    array_obj_ref_1759_index_0_resize_req_0 <= cp_elements(641);
    cp_elements(642) <= cp_elements(533);
    cpelement_group_643 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(642) & cp_elements(651));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(643),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1759_final_reg_req_0 <= cp_elements(643);
    cp_elements(644) <= cp_elements(533);
    array_obj_ref_1759_base_resize_req_0 <= cp_elements(644);
    cp_elements(645) <= array_obj_ref_1759_index_0_resize_ack_0;
    array_obj_ref_1759_index_0_rename_req_0 <= cp_elements(645);
    cp_elements(646) <= array_obj_ref_1759_index_0_rename_ack_0;
    array_obj_ref_1759_offset_inst_req_0 <= cp_elements(646);
    cp_elements(647) <= array_obj_ref_1759_offset_inst_ack_0;
    cp_elements(648) <= array_obj_ref_1759_base_resize_ack_0;
    cpelement_group_649 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(647) & cp_elements(648));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(649),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1759_root_address_inst_req_0 <= cp_elements(649);
    cp_elements(650) <= array_obj_ref_1759_root_address_inst_ack_0;
    array_obj_ref_1759_root_address_inst_req_1 <= cp_elements(650);
    cp_elements(651) <= array_obj_ref_1759_root_address_inst_ack_1;
    cp_elements(652) <= array_obj_ref_1759_final_reg_ack_0;
    cpelement_group_653 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(626) & cp_elements(636) & cp_elements(652) & cp_elements(657));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(653),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1762_gather_scatter_req_0 <= cp_elements(653);
    cp_elements(654) <= cp_elements(652);
    ptr_deref_1762_base_resize_req_0 <= cp_elements(654);
    cp_elements(655) <= ptr_deref_1762_base_resize_ack_0;
    ptr_deref_1762_root_address_inst_req_0 <= cp_elements(655);
    cp_elements(656) <= ptr_deref_1762_root_address_inst_ack_0;
    ptr_deref_1762_addr_0_req_0 <= cp_elements(656);
    cp_elements(657) <= ptr_deref_1762_addr_0_ack_0;
    cp_elements(658) <= ptr_deref_1762_gather_scatter_ack_0;
    ptr_deref_1762_store_0_req_0 <= cp_elements(658);
    cp_elements(659) <= ptr_deref_1762_store_0_ack_0;
    cp_elements(660) <= cp_elements(659);
    ptr_deref_1762_store_0_req_1 <= cp_elements(660);
    cp_elements(661) <= ptr_deref_1762_store_0_ack_1;
    cpelement_group_662 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(663) & cp_elements(664));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(662),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1769_inst_req_0 <= cp_elements(662);
    cp_elements(663) <= cp_elements(533);
    cp_elements(664) <= cp_elements(533);
    cp_elements(665) <= binary_1769_inst_ack_0;
    binary_1769_inst_req_1 <= cp_elements(665);
    cp_elements(666) <= binary_1769_inst_ack_1;
    cpelement_group_667 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(666) & cp_elements(668));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(667),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1773_inst_req_0 <= cp_elements(667);
    cp_elements(668) <= cp_elements(533);
    cp_elements(669) <= type_cast_1773_inst_ack_0;
    cpelement_group_670 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(671) & cp_elements(672));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(670),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1779_inst_req_0 <= cp_elements(670);
    cp_elements(671) <= cp_elements(533);
    cp_elements(672) <= cp_elements(533);
    cp_elements(673) <= binary_1779_inst_ack_0;
    binary_1779_inst_req_1 <= cp_elements(673);
    cp_elements(674) <= binary_1779_inst_ack_1;
    array_obj_ref_1783_index_0_resize_req_0 <= cp_elements(674);
    cp_elements(675) <= cp_elements(533);
    cpelement_group_676 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(675) & cp_elements(684));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(676),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1783_final_reg_req_0 <= cp_elements(676);
    cp_elements(677) <= cp_elements(533);
    array_obj_ref_1783_base_resize_req_0 <= cp_elements(677);
    cp_elements(678) <= array_obj_ref_1783_index_0_resize_ack_0;
    array_obj_ref_1783_index_0_rename_req_0 <= cp_elements(678);
    cp_elements(679) <= array_obj_ref_1783_index_0_rename_ack_0;
    array_obj_ref_1783_offset_inst_req_0 <= cp_elements(679);
    cp_elements(680) <= array_obj_ref_1783_offset_inst_ack_0;
    cp_elements(681) <= array_obj_ref_1783_base_resize_ack_0;
    cpelement_group_682 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(680) & cp_elements(681));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(682),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1783_root_address_inst_req_0 <= cp_elements(682);
    cp_elements(683) <= array_obj_ref_1783_root_address_inst_ack_0;
    array_obj_ref_1783_root_address_inst_req_1 <= cp_elements(683);
    cp_elements(684) <= array_obj_ref_1783_root_address_inst_ack_1;
    cp_elements(685) <= array_obj_ref_1783_final_reg_ack_0;
    cpelement_group_686 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(659) & cp_elements(669) & cp_elements(685) & cp_elements(690));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(686),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1786_gather_scatter_req_0 <= cp_elements(686);
    cp_elements(687) <= cp_elements(685);
    ptr_deref_1786_base_resize_req_0 <= cp_elements(687);
    cp_elements(688) <= ptr_deref_1786_base_resize_ack_0;
    ptr_deref_1786_root_address_inst_req_0 <= cp_elements(688);
    cp_elements(689) <= ptr_deref_1786_root_address_inst_ack_0;
    ptr_deref_1786_addr_0_req_0 <= cp_elements(689);
    cp_elements(690) <= ptr_deref_1786_addr_0_ack_0;
    cp_elements(691) <= ptr_deref_1786_gather_scatter_ack_0;
    ptr_deref_1786_store_0_req_0 <= cp_elements(691);
    cp_elements(692) <= ptr_deref_1786_store_0_ack_0;
    cp_elements(693) <= cp_elements(692);
    ptr_deref_1786_store_0_req_1 <= cp_elements(693);
    cp_elements(694) <= ptr_deref_1786_store_0_ack_1;
    cpelement_group_695 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(696) & cp_elements(697));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(695),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1793_inst_req_0 <= cp_elements(695);
    cp_elements(696) <= cp_elements(533);
    cp_elements(697) <= cp_elements(533);
    cp_elements(698) <= binary_1793_inst_ack_0;
    binary_1793_inst_req_1 <= cp_elements(698);
    cp_elements(699) <= binary_1793_inst_ack_1;
    cpelement_group_700 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(699) & cp_elements(701));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(700),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1797_inst_req_0 <= cp_elements(700);
    cp_elements(701) <= cp_elements(533);
    cp_elements(702) <= type_cast_1797_inst_ack_0;
    cpelement_group_703 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(704) & cp_elements(705));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(703),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1803_inst_req_0 <= cp_elements(703);
    cp_elements(704) <= cp_elements(533);
    cp_elements(705) <= cp_elements(533);
    cp_elements(706) <= binary_1803_inst_ack_0;
    binary_1803_inst_req_1 <= cp_elements(706);
    cp_elements(707) <= binary_1803_inst_ack_1;
    array_obj_ref_1807_index_0_resize_req_0 <= cp_elements(707);
    cp_elements(708) <= cp_elements(533);
    cpelement_group_709 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(708) & cp_elements(717));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(709),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1807_final_reg_req_0 <= cp_elements(709);
    cp_elements(710) <= cp_elements(533);
    array_obj_ref_1807_base_resize_req_0 <= cp_elements(710);
    cp_elements(711) <= array_obj_ref_1807_index_0_resize_ack_0;
    array_obj_ref_1807_index_0_rename_req_0 <= cp_elements(711);
    cp_elements(712) <= array_obj_ref_1807_index_0_rename_ack_0;
    array_obj_ref_1807_offset_inst_req_0 <= cp_elements(712);
    cp_elements(713) <= array_obj_ref_1807_offset_inst_ack_0;
    cp_elements(714) <= array_obj_ref_1807_base_resize_ack_0;
    cpelement_group_715 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(713) & cp_elements(714));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(715),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1807_root_address_inst_req_0 <= cp_elements(715);
    cp_elements(716) <= array_obj_ref_1807_root_address_inst_ack_0;
    array_obj_ref_1807_root_address_inst_req_1 <= cp_elements(716);
    cp_elements(717) <= array_obj_ref_1807_root_address_inst_ack_1;
    cp_elements(718) <= array_obj_ref_1807_final_reg_ack_0;
    cpelement_group_719 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(692) & cp_elements(702) & cp_elements(718) & cp_elements(723));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(719),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1810_gather_scatter_req_0 <= cp_elements(719);
    cp_elements(720) <= cp_elements(718);
    ptr_deref_1810_base_resize_req_0 <= cp_elements(720);
    cp_elements(721) <= ptr_deref_1810_base_resize_ack_0;
    ptr_deref_1810_root_address_inst_req_0 <= cp_elements(721);
    cp_elements(722) <= ptr_deref_1810_root_address_inst_ack_0;
    ptr_deref_1810_addr_0_req_0 <= cp_elements(722);
    cp_elements(723) <= ptr_deref_1810_addr_0_ack_0;
    cp_elements(724) <= ptr_deref_1810_gather_scatter_ack_0;
    ptr_deref_1810_store_0_req_0 <= cp_elements(724);
    cp_elements(725) <= ptr_deref_1810_store_0_ack_0;
    cp_elements(726) <= cp_elements(725);
    ptr_deref_1810_store_0_req_1 <= cp_elements(726);
    cp_elements(727) <= ptr_deref_1810_store_0_ack_1;
    cpelement_group_728 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(729) & cp_elements(730));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(728),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1817_inst_req_0 <= cp_elements(728);
    cp_elements(729) <= cp_elements(533);
    cp_elements(730) <= cp_elements(533);
    cp_elements(731) <= binary_1817_inst_ack_0;
    binary_1817_inst_req_1 <= cp_elements(731);
    cp_elements(732) <= binary_1817_inst_ack_1;
    cpelement_group_733 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(732) & cp_elements(734));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(733),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1821_inst_req_0 <= cp_elements(733);
    cp_elements(734) <= cp_elements(533);
    cp_elements(735) <= type_cast_1821_inst_ack_0;
    cpelement_group_736 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(737) & cp_elements(738));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(736),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1827_inst_req_0 <= cp_elements(736);
    cp_elements(737) <= cp_elements(533);
    cp_elements(738) <= cp_elements(533);
    cp_elements(739) <= binary_1827_inst_ack_0;
    binary_1827_inst_req_1 <= cp_elements(739);
    cp_elements(740) <= binary_1827_inst_ack_1;
    array_obj_ref_1831_index_0_resize_req_0 <= cp_elements(740);
    cp_elements(741) <= cp_elements(533);
    cpelement_group_742 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(741) & cp_elements(750));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(742),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1831_final_reg_req_0 <= cp_elements(742);
    cp_elements(743) <= cp_elements(533);
    array_obj_ref_1831_base_resize_req_0 <= cp_elements(743);
    cp_elements(744) <= array_obj_ref_1831_index_0_resize_ack_0;
    array_obj_ref_1831_index_0_rename_req_0 <= cp_elements(744);
    cp_elements(745) <= array_obj_ref_1831_index_0_rename_ack_0;
    array_obj_ref_1831_offset_inst_req_0 <= cp_elements(745);
    cp_elements(746) <= array_obj_ref_1831_offset_inst_ack_0;
    cp_elements(747) <= array_obj_ref_1831_base_resize_ack_0;
    cpelement_group_748 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(746) & cp_elements(747));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(748),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1831_root_address_inst_req_0 <= cp_elements(748);
    cp_elements(749) <= array_obj_ref_1831_root_address_inst_ack_0;
    array_obj_ref_1831_root_address_inst_req_1 <= cp_elements(749);
    cp_elements(750) <= array_obj_ref_1831_root_address_inst_ack_1;
    cp_elements(751) <= array_obj_ref_1831_final_reg_ack_0;
    cpelement_group_752 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(725) & cp_elements(735) & cp_elements(751) & cp_elements(756));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(752),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1834_gather_scatter_req_0 <= cp_elements(752);
    cp_elements(753) <= cp_elements(751);
    ptr_deref_1834_base_resize_req_0 <= cp_elements(753);
    cp_elements(754) <= ptr_deref_1834_base_resize_ack_0;
    ptr_deref_1834_root_address_inst_req_0 <= cp_elements(754);
    cp_elements(755) <= ptr_deref_1834_root_address_inst_ack_0;
    ptr_deref_1834_addr_0_req_0 <= cp_elements(755);
    cp_elements(756) <= ptr_deref_1834_addr_0_ack_0;
    cp_elements(757) <= ptr_deref_1834_gather_scatter_ack_0;
    ptr_deref_1834_store_0_req_0 <= cp_elements(757);
    cp_elements(758) <= ptr_deref_1834_store_0_ack_0;
    cp_elements(759) <= cp_elements(758);
    ptr_deref_1834_store_0_req_1 <= cp_elements(759);
    cp_elements(760) <= ptr_deref_1834_store_0_ack_1;
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(762) & cp_elements(763));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1839_inst_req_0 <= cp_elements(761);
    cp_elements(762) <= cp_elements(533);
    cp_elements(763) <= cp_elements(533);
    cp_elements(764) <= type_cast_1839_inst_ack_0;
    cpelement_group_765 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(766) & cp_elements(767));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(765),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1845_inst_req_0 <= cp_elements(765);
    cp_elements(766) <= cp_elements(533);
    cp_elements(767) <= cp_elements(533);
    cp_elements(768) <= binary_1845_inst_ack_0;
    binary_1845_inst_req_1 <= cp_elements(768);
    cp_elements(769) <= binary_1845_inst_ack_1;
    array_obj_ref_1849_index_0_resize_req_0 <= cp_elements(769);
    cp_elements(770) <= cp_elements(533);
    cpelement_group_771 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(770) & cp_elements(779));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(771),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1849_final_reg_req_0 <= cp_elements(771);
    cp_elements(772) <= cp_elements(533);
    array_obj_ref_1849_base_resize_req_0 <= cp_elements(772);
    cp_elements(773) <= array_obj_ref_1849_index_0_resize_ack_0;
    array_obj_ref_1849_index_0_rename_req_0 <= cp_elements(773);
    cp_elements(774) <= array_obj_ref_1849_index_0_rename_ack_0;
    array_obj_ref_1849_offset_inst_req_0 <= cp_elements(774);
    cp_elements(775) <= array_obj_ref_1849_offset_inst_ack_0;
    cp_elements(776) <= array_obj_ref_1849_base_resize_ack_0;
    cpelement_group_777 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(775) & cp_elements(776));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(777),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1849_root_address_inst_req_0 <= cp_elements(777);
    cp_elements(778) <= array_obj_ref_1849_root_address_inst_ack_0;
    array_obj_ref_1849_root_address_inst_req_1 <= cp_elements(778);
    cp_elements(779) <= array_obj_ref_1849_root_address_inst_ack_1;
    cp_elements(780) <= array_obj_ref_1849_final_reg_ack_0;
    cpelement_group_781 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(758) & cp_elements(764) & cp_elements(780) & cp_elements(785));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(781),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1852_gather_scatter_req_0 <= cp_elements(781);
    cp_elements(782) <= cp_elements(780);
    ptr_deref_1852_base_resize_req_0 <= cp_elements(782);
    cp_elements(783) <= ptr_deref_1852_base_resize_ack_0;
    ptr_deref_1852_root_address_inst_req_0 <= cp_elements(783);
    cp_elements(784) <= ptr_deref_1852_root_address_inst_ack_0;
    ptr_deref_1852_addr_0_req_0 <= cp_elements(784);
    cp_elements(785) <= ptr_deref_1852_addr_0_ack_0;
    cp_elements(786) <= ptr_deref_1852_gather_scatter_ack_0;
    ptr_deref_1852_store_0_req_0 <= cp_elements(786);
    cp_elements(787) <= ptr_deref_1852_store_0_ack_0;
    ptr_deref_1852_store_0_req_1 <= cp_elements(787);
    cp_elements(788) <= ptr_deref_1852_store_0_ack_1;
    cpelement_group_789 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(790) & cp_elements(791));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(789),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1859_inst_req_0 <= cp_elements(789);
    cp_elements(790) <= cp_elements(533);
    cp_elements(791) <= cp_elements(533);
    cp_elements(792) <= binary_1859_inst_ack_0;
    binary_1859_inst_req_1 <= cp_elements(792);
    cp_elements(793) <= binary_1859_inst_ack_1;
    cpelement_group_794 : Block -- 
      signal predecessors: BooleanArray(8 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(562) & cp_elements(595) & cp_elements(628) & cp_elements(661) & cp_elements(694) & cp_elements(727) & cp_elements(760) & cp_elements(788) & cp_elements(793));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(794),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(795) <= simple_obj_ref_1867_inst_ack_0;
    simple_obj_ref_1876_inst_req_0 <= cp_elements(795);
    cp_elements(796) <= simple_obj_ref_1876_inst_ack_0;
    simple_obj_ref_1885_inst_req_0 <= cp_elements(796);
    cp_elements(797) <= simple_obj_ref_1885_inst_ack_0;
    cp_elements(798) <= OrReduce(cp_elements(2) & cp_elements(34) & cp_elements(797));
    cp_elements(799) <= cp_elements(798);
    simple_obj_ref_1244_inst_req_0 <= cp_elements(799);
    cp_elements(800) <= false;
    cp_elements(801) <= cp_elements(800);
    cp_elements(802) <= type_cast_1336_inst_ack_0;
    phi_stmt_1330_req_1 <= cp_elements(802);
    cp_elements(803) <= OrReduce(cp_elements(4) & cp_elements(802));
    cp_elements(804) <= cp_elements(803);
    cp_elements(805) <= phi_stmt_1330_ack_0;
    cp_elements(806) <= false;
    cp_elements(807) <= cp_elements(806);
    cp_elements(808) <= OrReduce(cp_elements(6) & cp_elements(7));
    cp_elements(809) <= cp_elements(808);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1292_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1292_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1292_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1297_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1297_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1297_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1302_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1302_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1302_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1307_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1307_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1307_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1316_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1316_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1316_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1321_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1321_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1321_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1326_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1326_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1326_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1529_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1529_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1529_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1529_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1533_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1533_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1533_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1533_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1537_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1537_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1537_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1537_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1541_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1541_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1541_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1541_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1545_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1545_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1545_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1545_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1549_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1549_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1549_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1549_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1553_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1553_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1553_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1553_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1557_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1557_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1557_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1557_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1687_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1687_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1687_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1687_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1711_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1735_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1735_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1735_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1735_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1759_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1759_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1759_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1759_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1783_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1783_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1783_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1783_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1807_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1807_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1807_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1807_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1831_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1831_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1831_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1831_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1849_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1849_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_1849_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1849_root_address : std_logic_vector(10 downto 0);
    signal expr_1368_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1368_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_1371_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1371_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal iNsTr_0_1230 : std_logic_vector(31 downto 0);
    signal iNsTr_10_1349 : std_logic_vector(31 downto 0);
    signal iNsTr_11_1358 : std_logic_vector(31 downto 0);
    signal iNsTr_21_1866 : std_logic_vector(31 downto 0);
    signal iNsTr_23_1875 : std_logic_vector(31 downto 0);
    signal iNsTr_25_1884 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1243 : std_logic_vector(31 downto 0);
    signal iNsTr_5_1253 : std_logic_vector(31 downto 0);
    signal iNsTr_7_1275 : std_logic_vector(31 downto 0);
    signal iNsTr_9_1330 : std_logic_vector(31 downto 0);
    signal ptr_deref_1232_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1232_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1232_word_address_0 : std_logic_vector(3 downto 0);
    signal ptr_deref_1388_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1388_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1388_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1388_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1388_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1388_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1402_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1402_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1402_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1402_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1402_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1402_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1416_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1416_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1416_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1416_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1416_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1430_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1430_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1430_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1430_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1430_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1430_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1444_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1444_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1444_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1444_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1444_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1444_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1458_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1458_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1458_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1458_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1458_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1472_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1472_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1472_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1472_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1472_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1472_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1480_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1480_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1480_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1480_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1480_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1480_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1570_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1570_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1570_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1570_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1570_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1570_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1584_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1584_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1584_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1584_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1584_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1584_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1598_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1598_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1598_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1598_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1598_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1598_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1612_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1612_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1612_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1612_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1612_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1612_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1626_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1626_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1626_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1640_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1640_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1640_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1640_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1640_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1640_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1654_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1654_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1654_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1654_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1654_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1654_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1662_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1662_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1662_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1662_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1662_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1662_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1690_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1690_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1690_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1690_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1690_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1690_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1714_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1714_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1714_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1714_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1714_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1714_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1738_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1738_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1738_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1738_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1738_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1762_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1762_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1762_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1762_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1762_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1762_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1786_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1786_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1786_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1786_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1786_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1786_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1810_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1810_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1810_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1810_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1810_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1810_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1834_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1834_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1834_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1834_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1834_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1834_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1852_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1852_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1852_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1852_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1852_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1852_word_offset_0 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1528_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1528_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1532_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1532_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1536_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1536_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1540_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1540_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1544_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1544_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1548_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1548_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1552_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1552_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1556_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1556_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1686_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1686_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1710_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1710_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1734_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1734_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1758_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1758_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1782_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1782_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1806_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1806_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1830_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1830_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1848_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_1848_scaled : std_logic_vector(10 downto 0);
    signal tmp102_1550 : std_logic_vector(31 downto 0);
    signal tmp105_1554 : std_logic_vector(31 downto 0);
    signal tmp108_1558 : std_logic_vector(31 downto 0);
    signal tmp10_1424 : std_logic_vector(63 downto 0);
    signal tmp112_1688 : std_logic_vector(31 downto 0);
    signal tmp114_1708 : std_logic_vector(31 downto 0);
    signal tmp115_1712 : std_logic_vector(31 downto 0);
    signal tmp117_1732 : std_logic_vector(31 downto 0);
    signal tmp118_1736 : std_logic_vector(31 downto 0);
    signal tmp11_1428 : std_logic_vector(7 downto 0);
    signal tmp120_1756 : std_logic_vector(31 downto 0);
    signal tmp121_1760 : std_logic_vector(31 downto 0);
    signal tmp123_1780 : std_logic_vector(31 downto 0);
    signal tmp124_1784 : std_logic_vector(31 downto 0);
    signal tmp126_1804 : std_logic_vector(31 downto 0);
    signal tmp127_1808 : std_logic_vector(31 downto 0);
    signal tmp129_1828 : std_logic_vector(31 downto 0);
    signal tmp130_1832 : std_logic_vector(31 downto 0);
    signal tmp132_1846 : std_logic_vector(31 downto 0);
    signal tmp133_1850 : std_logic_vector(31 downto 0);
    signal tmp134_1860 : std_logic_vector(31 downto 0);
    signal tmp136143_1526 : std_logic_vector(31 downto 0);
    signal tmp137144_1520 : std_logic_vector(31 downto 0);
    signal tmp138145_1514 : std_logic_vector(31 downto 0);
    signal tmp139146_1508 : std_logic_vector(31 downto 0);
    signal tmp13_1438 : std_logic_vector(63 downto 0);
    signal tmp140147_1502 : std_logic_vector(31 downto 0);
    signal tmp141148_1496 : std_logic_vector(31 downto 0);
    signal tmp142149_1490 : std_logic_vector(31 downto 0);
    signal tmp14_1442 : std_logic_vector(7 downto 0);
    signal tmp16_1452 : std_logic_vector(63 downto 0);
    signal tmp17_1456 : std_logic_vector(7 downto 0);
    signal tmp19_1466 : std_logic_vector(63 downto 0);
    signal tmp1_1382 : std_logic_vector(63 downto 0);
    signal tmp20_1470 : std_logic_vector(7 downto 0);
    signal tmp22_1478 : std_logic_vector(7 downto 0);
    signal tmp24_1564 : std_logic_vector(63 downto 0);
    signal tmp25_1568 : std_logic_vector(7 downto 0);
    signal tmp27_1578 : std_logic_vector(63 downto 0);
    signal tmp28_1582 : std_logic_vector(7 downto 0);
    signal tmp2_1386 : std_logic_vector(7 downto 0);
    signal tmp2x_xi_1262 : std_logic_vector(0 downto 0);
    signal tmp30_1592 : std_logic_vector(63 downto 0);
    signal tmp31_1596 : std_logic_vector(7 downto 0);
    signal tmp33_1606 : std_logic_vector(63 downto 0);
    signal tmp34_1610 : std_logic_vector(7 downto 0);
    signal tmp36_1620 : std_logic_vector(63 downto 0);
    signal tmp37_1624 : std_logic_vector(7 downto 0);
    signal tmp39_1634 : std_logic_vector(63 downto 0);
    signal tmp40_1638 : std_logic_vector(7 downto 0);
    signal tmp42_1648 : std_logic_vector(63 downto 0);
    signal tmp43_1652 : std_logic_vector(7 downto 0);
    signal tmp45_1660 : std_logic_vector(7 downto 0);
    signal tmp47_1680 : std_logic_vector(63 downto 0);
    signal tmp48_1684 : std_logic_vector(7 downto 0);
    signal tmp4_1396 : std_logic_vector(63 downto 0);
    signal tmp4x_xi_1278 : std_logic_vector(31 downto 0);
    signal tmp50_1698 : std_logic_vector(63 downto 0);
    signal tmp51_1702 : std_logic_vector(7 downto 0);
    signal tmp53_1722 : std_logic_vector(63 downto 0);
    signal tmp54_1726 : std_logic_vector(7 downto 0);
    signal tmp56_1746 : std_logic_vector(63 downto 0);
    signal tmp57_1750 : std_logic_vector(7 downto 0);
    signal tmp59_1770 : std_logic_vector(63 downto 0);
    signal tmp5_1400 : std_logic_vector(7 downto 0);
    signal tmp5x_xi_1283 : std_logic_vector(31 downto 0);
    signal tmp60_1774 : std_logic_vector(7 downto 0);
    signal tmp62_1794 : std_logic_vector(63 downto 0);
    signal tmp63_1798 : std_logic_vector(7 downto 0);
    signal tmp65_1818 : std_logic_vector(63 downto 0);
    signal tmp66_1822 : std_logic_vector(7 downto 0);
    signal tmp68_1840 : std_logic_vector(7 downto 0);
    signal tmp70_1288 : std_logic_vector(31 downto 0);
    signal tmp72_1352 : std_logic_vector(63 downto 0);
    signal tmp73_1361 : std_logic_vector(7 downto 0);
    signal tmp74_1365 : std_logic_vector(31 downto 0);
    signal tmp76_1293 : std_logic_vector(31 downto 0);
    signal tmp77_1298 : std_logic_vector(31 downto 0);
    signal tmp78_1303 : std_logic_vector(31 downto 0);
    signal tmp79_1308 : std_logic_vector(31 downto 0);
    signal tmp7_1410 : std_logic_vector(63 downto 0);
    signal tmp80_1312 : std_logic_vector(31 downto 0);
    signal tmp81_1317 : std_logic_vector(31 downto 0);
    signal tmp82_1322 : std_logic_vector(31 downto 0);
    signal tmp83_1327 : std_logic_vector(31 downto 0);
    signal tmp87_1530 : std_logic_vector(31 downto 0);
    signal tmp8_1414 : std_logic_vector(7 downto 0);
    signal tmp90_1534 : std_logic_vector(31 downto 0);
    signal tmp93_1538 : std_logic_vector(31 downto 0);
    signal tmp96_1542 : std_logic_vector(31 downto 0);
    signal tmp99_1546 : std_logic_vector(31 downto 0);
    signal tmp_1343 : std_logic_vector(31 downto 0);
    signal tmpx_xi_1256 : std_logic_vector(7 downto 0);
    signal type_cast_1234_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1246_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1260_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1334_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1336_wire : std_logic_vector(31 downto 0);
    signal type_cast_1341_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1380_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1394_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1408_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1422_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1436_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1450_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1464_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1488_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1494_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1500_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1506_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1512_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1518_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1524_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1576_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1590_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1604_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1618_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1632_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1646_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1670_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1678_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1696_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1706_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1720_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1730_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1744_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1754_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1768_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1778_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1792_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1802_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1816_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1826_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1844_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1858_wire_constant : std_logic_vector(31 downto 0);
    signal wordx_x0x_xbe_1672 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1292_final_offset <= "00000000001";
    array_obj_ref_1297_final_offset <= "00000000010";
    array_obj_ref_1302_final_offset <= "00000000011";
    array_obj_ref_1307_final_offset <= "00000000100";
    array_obj_ref_1316_final_offset <= "00000000101";
    array_obj_ref_1321_final_offset <= "00000000110";
    array_obj_ref_1326_final_offset <= "00000000111";
    array_obj_ref_1529_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1533_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1537_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1541_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1545_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1549_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1553_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1557_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1687_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1711_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1735_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1759_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1783_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1807_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1831_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_1849_offset_scale_factor_0 <= "00000000001";
    expr_1368_wire_constant <= "00000000000000000000000011111111";
    expr_1371_wire_constant <= "00000000000000000000000000000000";
    iNsTr_0_1230 <= "00000000000000000000000000000000";
    iNsTr_10_1349 <= "00000000000000000000000000000000";
    iNsTr_11_1358 <= "00000000000000000000000000000000";
    iNsTr_21_1866 <= "00000000000000000000000000000000";
    iNsTr_23_1875 <= "00000000000000000000000000000000";
    iNsTr_25_1884 <= "00000000000000000000000000000000";
    iNsTr_3_1243 <= "00000000000000000000000000000000";
    iNsTr_5_1253 <= "00000000000000000000000000000000";
    iNsTr_7_1275 <= "00000000000000000000000000000000";
    ptr_deref_1232_word_address_0 <= "0000";
    ptr_deref_1388_word_offset_0 <= "00000000000";
    ptr_deref_1402_word_offset_0 <= "00000000000";
    ptr_deref_1416_word_offset_0 <= "00000000000";
    ptr_deref_1430_word_offset_0 <= "00000000000";
    ptr_deref_1444_word_offset_0 <= "00000000000";
    ptr_deref_1458_word_offset_0 <= "00000000000";
    ptr_deref_1472_word_offset_0 <= "00000000000";
    ptr_deref_1480_word_offset_0 <= "00000000000";
    ptr_deref_1570_word_offset_0 <= "00000000000";
    ptr_deref_1584_word_offset_0 <= "00000000000";
    ptr_deref_1598_word_offset_0 <= "00000000000";
    ptr_deref_1612_word_offset_0 <= "00000000000";
    ptr_deref_1626_word_offset_0 <= "00000000000";
    ptr_deref_1640_word_offset_0 <= "00000000000";
    ptr_deref_1654_word_offset_0 <= "00000000000";
    ptr_deref_1662_word_offset_0 <= "00000000000";
    ptr_deref_1690_word_offset_0 <= "00000000000";
    ptr_deref_1714_word_offset_0 <= "00000000000";
    ptr_deref_1738_word_offset_0 <= "00000000000";
    ptr_deref_1762_word_offset_0 <= "00000000000";
    ptr_deref_1786_word_offset_0 <= "00000000000";
    ptr_deref_1810_word_offset_0 <= "00000000000";
    ptr_deref_1834_word_offset_0 <= "00000000000";
    ptr_deref_1852_word_offset_0 <= "00000000000";
    type_cast_1234_wire_constant <= "00000001";
    type_cast_1246_wire_constant <= "00000010";
    type_cast_1260_wire_constant <= "00000011";
    type_cast_1334_wire_constant <= "00000000000000000000000000000000";
    type_cast_1341_wire_constant <= "00000000000000000000000000000011";
    type_cast_1380_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1394_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1408_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1422_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1436_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1450_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1464_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1488_wire_constant <= "00000000000000000000000000000001";
    type_cast_1494_wire_constant <= "00000000000000000000000000000010";
    type_cast_1500_wire_constant <= "00000000000000000000000000000011";
    type_cast_1506_wire_constant <= "00000000000000000000000000000100";
    type_cast_1512_wire_constant <= "00000000000000000000000000000101";
    type_cast_1518_wire_constant <= "00000000000000000000000000000110";
    type_cast_1524_wire_constant <= "00000000000000000000000000000111";
    type_cast_1562_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1576_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1590_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1604_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1618_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1632_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1646_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1670_wire_constant <= "00000000000000000000000000000001";
    type_cast_1678_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_1696_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_1706_wire_constant <= "00000000000000000000000000000001";
    type_cast_1720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_1730_wire_constant <= "00000000000000000000000000000010";
    type_cast_1744_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_1754_wire_constant <= "00000000000000000000000000000011";
    type_cast_1768_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_1778_wire_constant <= "00000000000000000000000000000100";
    type_cast_1792_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1802_wire_constant <= "00000000000000000000000000000101";
    type_cast_1816_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1826_wire_constant <= "00000000000000000000000000000110";
    type_cast_1844_wire_constant <= "00000000000000000000000000000111";
    type_cast_1858_wire_constant <= "00000000000000000000000000000001";
    phi_stmt_1330: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1334_wire_constant & type_cast_1336_wire;
      req <= phi_stmt_1330_req_0 & phi_stmt_1330_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1330_ack_0,
          idata => idata,
          odata => iNsTr_9_1330,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1330
    array_obj_ref_1292_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1292_resized_base_address, req => array_obj_ref_1292_base_resize_req_0, ack => array_obj_ref_1292_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1292_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1292_root_address, dout => tmp76_1293, req => array_obj_ref_1292_final_reg_req_0, ack => array_obj_ref_1292_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1297_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1297_resized_base_address, req => array_obj_ref_1297_base_resize_req_0, ack => array_obj_ref_1297_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1297_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1297_root_address, dout => tmp77_1298, req => array_obj_ref_1297_final_reg_req_0, ack => array_obj_ref_1297_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1302_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1302_resized_base_address, req => array_obj_ref_1302_base_resize_req_0, ack => array_obj_ref_1302_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1302_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1302_root_address, dout => tmp78_1303, req => array_obj_ref_1302_final_reg_req_0, ack => array_obj_ref_1302_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1307_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp5x_xi_1283, dout => array_obj_ref_1307_resized_base_address, req => array_obj_ref_1307_base_resize_req_0, ack => array_obj_ref_1307_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1307_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1307_root_address, dout => tmp79_1308, req => array_obj_ref_1307_final_reg_req_0, ack => array_obj_ref_1307_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1316_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1316_resized_base_address, req => array_obj_ref_1316_base_resize_req_0, ack => array_obj_ref_1316_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1316_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1316_root_address, dout => tmp81_1317, req => array_obj_ref_1316_final_reg_req_0, ack => array_obj_ref_1316_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1321_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1321_resized_base_address, req => array_obj_ref_1321_base_resize_req_0, ack => array_obj_ref_1321_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1321_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1321_root_address, dout => tmp82_1322, req => array_obj_ref_1321_final_reg_req_0, ack => array_obj_ref_1321_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1326_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1326_resized_base_address, req => array_obj_ref_1326_base_resize_req_0, ack => array_obj_ref_1326_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1326_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1326_root_address, dout => tmp83_1327, req => array_obj_ref_1326_final_reg_req_0, ack => array_obj_ref_1326_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1529_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1529_resized_base_address, req => array_obj_ref_1529_base_resize_req_0, ack => array_obj_ref_1529_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1529_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1529_root_address, dout => tmp87_1530, req => array_obj_ref_1529_final_reg_req_0, ack => array_obj_ref_1529_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1529_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp_1343, dout => simple_obj_ref_1528_resized, req => array_obj_ref_1529_index_0_resize_req_0, ack => array_obj_ref_1529_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1529_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1528_scaled, dout => array_obj_ref_1529_final_offset, req => array_obj_ref_1529_offset_inst_req_0, ack => array_obj_ref_1529_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1533_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1533_resized_base_address, req => array_obj_ref_1533_base_resize_req_0, ack => array_obj_ref_1533_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1533_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1533_root_address, dout => tmp90_1534, req => array_obj_ref_1533_final_reg_req_0, ack => array_obj_ref_1533_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1533_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp142149_1490, dout => simple_obj_ref_1532_resized, req => array_obj_ref_1533_index_0_resize_req_0, ack => array_obj_ref_1533_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1533_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1532_scaled, dout => array_obj_ref_1533_final_offset, req => array_obj_ref_1533_offset_inst_req_0, ack => array_obj_ref_1533_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1537_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1537_resized_base_address, req => array_obj_ref_1537_base_resize_req_0, ack => array_obj_ref_1537_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1537_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1537_root_address, dout => tmp93_1538, req => array_obj_ref_1537_final_reg_req_0, ack => array_obj_ref_1537_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1537_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp141148_1496, dout => simple_obj_ref_1536_resized, req => array_obj_ref_1537_index_0_resize_req_0, ack => array_obj_ref_1537_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1537_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1536_scaled, dout => array_obj_ref_1537_final_offset, req => array_obj_ref_1537_offset_inst_req_0, ack => array_obj_ref_1537_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1541_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1541_resized_base_address, req => array_obj_ref_1541_base_resize_req_0, ack => array_obj_ref_1541_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1541_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1541_root_address, dout => tmp96_1542, req => array_obj_ref_1541_final_reg_req_0, ack => array_obj_ref_1541_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1541_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp140147_1502, dout => simple_obj_ref_1540_resized, req => array_obj_ref_1541_index_0_resize_req_0, ack => array_obj_ref_1541_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1541_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1540_scaled, dout => array_obj_ref_1541_final_offset, req => array_obj_ref_1541_offset_inst_req_0, ack => array_obj_ref_1541_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1545_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1545_resized_base_address, req => array_obj_ref_1545_base_resize_req_0, ack => array_obj_ref_1545_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1545_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1545_root_address, dout => tmp99_1546, req => array_obj_ref_1545_final_reg_req_0, ack => array_obj_ref_1545_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1545_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp139146_1508, dout => simple_obj_ref_1544_resized, req => array_obj_ref_1545_index_0_resize_req_0, ack => array_obj_ref_1545_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1545_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1544_scaled, dout => array_obj_ref_1545_final_offset, req => array_obj_ref_1545_offset_inst_req_0, ack => array_obj_ref_1545_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1549_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1549_resized_base_address, req => array_obj_ref_1549_base_resize_req_0, ack => array_obj_ref_1549_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1549_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1549_root_address, dout => tmp102_1550, req => array_obj_ref_1549_final_reg_req_0, ack => array_obj_ref_1549_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1549_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp138145_1514, dout => simple_obj_ref_1548_resized, req => array_obj_ref_1549_index_0_resize_req_0, ack => array_obj_ref_1549_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1549_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1548_scaled, dout => array_obj_ref_1549_final_offset, req => array_obj_ref_1549_offset_inst_req_0, ack => array_obj_ref_1549_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1553_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1553_resized_base_address, req => array_obj_ref_1553_base_resize_req_0, ack => array_obj_ref_1553_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1553_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1553_root_address, dout => tmp105_1554, req => array_obj_ref_1553_final_reg_req_0, ack => array_obj_ref_1553_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1553_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp137144_1520, dout => simple_obj_ref_1552_resized, req => array_obj_ref_1553_index_0_resize_req_0, ack => array_obj_ref_1553_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1553_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1552_scaled, dout => array_obj_ref_1553_final_offset, req => array_obj_ref_1553_offset_inst_req_0, ack => array_obj_ref_1553_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1557_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1557_resized_base_address, req => array_obj_ref_1557_base_resize_req_0, ack => array_obj_ref_1557_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1557_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1557_root_address, dout => tmp108_1558, req => array_obj_ref_1557_final_reg_req_0, ack => array_obj_ref_1557_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1557_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp136143_1526, dout => simple_obj_ref_1556_resized, req => array_obj_ref_1557_index_0_resize_req_0, ack => array_obj_ref_1557_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1557_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1556_scaled, dout => array_obj_ref_1557_final_offset, req => array_obj_ref_1557_offset_inst_req_0, ack => array_obj_ref_1557_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1687_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1687_resized_base_address, req => array_obj_ref_1687_base_resize_req_0, ack => array_obj_ref_1687_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1687_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1687_root_address, dout => tmp112_1688, req => array_obj_ref_1687_final_reg_req_0, ack => array_obj_ref_1687_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1687_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp_1343, dout => simple_obj_ref_1686_resized, req => array_obj_ref_1687_index_0_resize_req_0, ack => array_obj_ref_1687_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1687_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1686_scaled, dout => array_obj_ref_1687_final_offset, req => array_obj_ref_1687_offset_inst_req_0, ack => array_obj_ref_1687_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1711_resized_base_address, req => array_obj_ref_1711_base_resize_req_0, ack => array_obj_ref_1711_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1711_root_address, dout => tmp115_1712, req => array_obj_ref_1711_final_reg_req_0, ack => array_obj_ref_1711_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp114_1708, dout => simple_obj_ref_1710_resized, req => array_obj_ref_1711_index_0_resize_req_0, ack => array_obj_ref_1711_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1711_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1710_scaled, dout => array_obj_ref_1711_final_offset, req => array_obj_ref_1711_offset_inst_req_0, ack => array_obj_ref_1711_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1735_resized_base_address, req => array_obj_ref_1735_base_resize_req_0, ack => array_obj_ref_1735_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1735_root_address, dout => tmp118_1736, req => array_obj_ref_1735_final_reg_req_0, ack => array_obj_ref_1735_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp117_1732, dout => simple_obj_ref_1734_resized, req => array_obj_ref_1735_index_0_resize_req_0, ack => array_obj_ref_1735_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1735_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1734_scaled, dout => array_obj_ref_1735_final_offset, req => array_obj_ref_1735_offset_inst_req_0, ack => array_obj_ref_1735_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1759_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1759_resized_base_address, req => array_obj_ref_1759_base_resize_req_0, ack => array_obj_ref_1759_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1759_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1759_root_address, dout => tmp121_1760, req => array_obj_ref_1759_final_reg_req_0, ack => array_obj_ref_1759_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1759_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp120_1756, dout => simple_obj_ref_1758_resized, req => array_obj_ref_1759_index_0_resize_req_0, ack => array_obj_ref_1759_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1759_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1758_scaled, dout => array_obj_ref_1759_final_offset, req => array_obj_ref_1759_offset_inst_req_0, ack => array_obj_ref_1759_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1783_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1783_resized_base_address, req => array_obj_ref_1783_base_resize_req_0, ack => array_obj_ref_1783_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1783_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1783_root_address, dout => tmp124_1784, req => array_obj_ref_1783_final_reg_req_0, ack => array_obj_ref_1783_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1783_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp123_1780, dout => simple_obj_ref_1782_resized, req => array_obj_ref_1783_index_0_resize_req_0, ack => array_obj_ref_1783_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1783_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1782_scaled, dout => array_obj_ref_1783_final_offset, req => array_obj_ref_1783_offset_inst_req_0, ack => array_obj_ref_1783_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1807_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1807_resized_base_address, req => array_obj_ref_1807_base_resize_req_0, ack => array_obj_ref_1807_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1807_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1807_root_address, dout => tmp127_1808, req => array_obj_ref_1807_final_reg_req_0, ack => array_obj_ref_1807_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1807_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp126_1804, dout => simple_obj_ref_1806_resized, req => array_obj_ref_1807_index_0_resize_req_0, ack => array_obj_ref_1807_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1807_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1806_scaled, dout => array_obj_ref_1807_final_offset, req => array_obj_ref_1807_offset_inst_req_0, ack => array_obj_ref_1807_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1831_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1831_resized_base_address, req => array_obj_ref_1831_base_resize_req_0, ack => array_obj_ref_1831_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1831_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1831_root_address, dout => tmp130_1832, req => array_obj_ref_1831_final_reg_req_0, ack => array_obj_ref_1831_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1831_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp129_1828, dout => simple_obj_ref_1830_resized, req => array_obj_ref_1831_index_0_resize_req_0, ack => array_obj_ref_1831_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1831_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1830_scaled, dout => array_obj_ref_1831_final_offset, req => array_obj_ref_1831_offset_inst_req_0, ack => array_obj_ref_1831_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1849_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => array_obj_ref_1849_resized_base_address, req => array_obj_ref_1849_base_resize_req_0, ack => array_obj_ref_1849_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1849_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1849_root_address, dout => tmp133_1850, req => array_obj_ref_1849_final_reg_req_0, ack => array_obj_ref_1849_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1849_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp132_1846, dout => simple_obj_ref_1848_resized, req => array_obj_ref_1849_index_0_resize_req_0, ack => array_obj_ref_1849_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1849_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_1848_scaled, dout => array_obj_ref_1849_final_offset, req => array_obj_ref_1849_offset_inst_req_0, ack => array_obj_ref_1849_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1388_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp70_1288, dout => ptr_deref_1388_resized_base_address, req => ptr_deref_1388_base_resize_req_0, ack => ptr_deref_1388_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1402_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp76_1293, dout => ptr_deref_1402_resized_base_address, req => ptr_deref_1402_base_resize_req_0, ack => ptr_deref_1402_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1416_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp77_1298, dout => ptr_deref_1416_resized_base_address, req => ptr_deref_1416_base_resize_req_0, ack => ptr_deref_1416_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1430_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp78_1303, dout => ptr_deref_1430_resized_base_address, req => ptr_deref_1430_base_resize_req_0, ack => ptr_deref_1430_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1444_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp80_1312, dout => ptr_deref_1444_resized_base_address, req => ptr_deref_1444_base_resize_req_0, ack => ptr_deref_1444_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1458_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp81_1317, dout => ptr_deref_1458_resized_base_address, req => ptr_deref_1458_base_resize_req_0, ack => ptr_deref_1458_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1472_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp82_1322, dout => ptr_deref_1472_resized_base_address, req => ptr_deref_1472_base_resize_req_0, ack => ptr_deref_1472_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1480_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp83_1327, dout => ptr_deref_1480_resized_base_address, req => ptr_deref_1480_base_resize_req_0, ack => ptr_deref_1480_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1570_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp87_1530, dout => ptr_deref_1570_resized_base_address, req => ptr_deref_1570_base_resize_req_0, ack => ptr_deref_1570_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1584_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp90_1534, dout => ptr_deref_1584_resized_base_address, req => ptr_deref_1584_base_resize_req_0, ack => ptr_deref_1584_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1598_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp93_1538, dout => ptr_deref_1598_resized_base_address, req => ptr_deref_1598_base_resize_req_0, ack => ptr_deref_1598_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1612_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp96_1542, dout => ptr_deref_1612_resized_base_address, req => ptr_deref_1612_base_resize_req_0, ack => ptr_deref_1612_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1626_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp99_1546, dout => ptr_deref_1626_resized_base_address, req => ptr_deref_1626_base_resize_req_0, ack => ptr_deref_1626_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1640_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp102_1550, dout => ptr_deref_1640_resized_base_address, req => ptr_deref_1640_base_resize_req_0, ack => ptr_deref_1640_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1654_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp105_1554, dout => ptr_deref_1654_resized_base_address, req => ptr_deref_1654_base_resize_req_0, ack => ptr_deref_1654_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1662_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp108_1558, dout => ptr_deref_1662_resized_base_address, req => ptr_deref_1662_base_resize_req_0, ack => ptr_deref_1662_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1690_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp112_1688, dout => ptr_deref_1690_resized_base_address, req => ptr_deref_1690_base_resize_req_0, ack => ptr_deref_1690_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1714_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp115_1712, dout => ptr_deref_1714_resized_base_address, req => ptr_deref_1714_base_resize_req_0, ack => ptr_deref_1714_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1738_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp118_1736, dout => ptr_deref_1738_resized_base_address, req => ptr_deref_1738_base_resize_req_0, ack => ptr_deref_1738_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1762_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp121_1760, dout => ptr_deref_1762_resized_base_address, req => ptr_deref_1762_base_resize_req_0, ack => ptr_deref_1762_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1786_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1784, dout => ptr_deref_1786_resized_base_address, req => ptr_deref_1786_base_resize_req_0, ack => ptr_deref_1786_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1810_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp127_1808, dout => ptr_deref_1810_resized_base_address, req => ptr_deref_1810_base_resize_req_0, ack => ptr_deref_1810_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1834_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp130_1832, dout => ptr_deref_1834_resized_base_address, req => ptr_deref_1834_base_resize_req_0, ack => ptr_deref_1834_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1852_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp133_1850, dout => ptr_deref_1852_resized_base_address, req => ptr_deref_1852_base_resize_req_0, ack => ptr_deref_1852_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1282_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1278, dout => tmp5x_xi_1283, req => type_cast_1282_inst_req_0, ack => type_cast_1282_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1287_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp4x_xi_1278, dout => tmp70_1288, req => type_cast_1287_inst_req_0, ack => type_cast_1287_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1311_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp79_1308, dout => tmp80_1312, req => type_cast_1311_inst_req_0, ack => type_cast_1311_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1336_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => wordx_x0x_xbe_1672, dout => type_cast_1336_wire, req => type_cast_1336_inst_req_0, ack => type_cast_1336_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1364_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp73_1361, dout => tmp74_1365, req => type_cast_1364_inst_req_0, ack => type_cast_1364_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1385_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp1_1382, dout => tmp2_1386, req => type_cast_1385_inst_req_0, ack => type_cast_1385_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1399_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp4_1396, dout => tmp5_1400, req => type_cast_1399_inst_req_0, ack => type_cast_1399_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1413_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp7_1410, dout => tmp8_1414, req => type_cast_1413_inst_req_0, ack => type_cast_1413_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1427_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp10_1424, dout => tmp11_1428, req => type_cast_1427_inst_req_0, ack => type_cast_1427_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1441_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp13_1438, dout => tmp14_1442, req => type_cast_1441_inst_req_0, ack => type_cast_1441_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1455_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp16_1452, dout => tmp17_1456, req => type_cast_1455_inst_req_0, ack => type_cast_1455_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1469_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp19_1466, dout => tmp20_1470, req => type_cast_1469_inst_req_0, ack => type_cast_1469_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1477_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp72_1352, dout => tmp22_1478, req => type_cast_1477_inst_req_0, ack => type_cast_1477_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1567_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp24_1564, dout => tmp25_1568, req => type_cast_1567_inst_req_0, ack => type_cast_1567_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1581_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp27_1578, dout => tmp28_1582, req => type_cast_1581_inst_req_0, ack => type_cast_1581_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1595_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp30_1592, dout => tmp31_1596, req => type_cast_1595_inst_req_0, ack => type_cast_1595_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1609_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp33_1606, dout => tmp34_1610, req => type_cast_1609_inst_req_0, ack => type_cast_1609_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1623_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp36_1620, dout => tmp37_1624, req => type_cast_1623_inst_req_0, ack => type_cast_1623_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1637_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp39_1634, dout => tmp40_1638, req => type_cast_1637_inst_req_0, ack => type_cast_1637_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1651_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp42_1648, dout => tmp43_1652, req => type_cast_1651_inst_req_0, ack => type_cast_1651_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1659_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp72_1352, dout => tmp45_1660, req => type_cast_1659_inst_req_0, ack => type_cast_1659_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1683_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp47_1680, dout => tmp48_1684, req => type_cast_1683_inst_req_0, ack => type_cast_1683_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1701_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp50_1698, dout => tmp51_1702, req => type_cast_1701_inst_req_0, ack => type_cast_1701_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1725_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp53_1722, dout => tmp54_1726, req => type_cast_1725_inst_req_0, ack => type_cast_1725_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1749_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp56_1746, dout => tmp57_1750, req => type_cast_1749_inst_req_0, ack => type_cast_1749_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1773_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp59_1770, dout => tmp60_1774, req => type_cast_1773_inst_req_0, ack => type_cast_1773_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1797_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp62_1794, dout => tmp63_1798, req => type_cast_1797_inst_req_0, ack => type_cast_1797_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1821_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp65_1818, dout => tmp66_1822, req => type_cast_1821_inst_req_0, ack => type_cast_1821_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1839_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => false ) 
      port map( din => tmp72_1352, dout => tmp68_1840, req => type_cast_1839_inst_req_0, ack => type_cast_1839_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1529_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1529_index_0_rename_ack_0 <= array_obj_ref_1529_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1528_resized;
      simple_obj_ref_1528_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1533_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1533_index_0_rename_ack_0 <= array_obj_ref_1533_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1532_resized;
      simple_obj_ref_1532_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1537_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1537_index_0_rename_ack_0 <= array_obj_ref_1537_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1536_resized;
      simple_obj_ref_1536_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1541_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1541_index_0_rename_ack_0 <= array_obj_ref_1541_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1540_resized;
      simple_obj_ref_1540_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1545_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1545_index_0_rename_ack_0 <= array_obj_ref_1545_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1544_resized;
      simple_obj_ref_1544_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1549_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1549_index_0_rename_ack_0 <= array_obj_ref_1549_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1548_resized;
      simple_obj_ref_1548_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1553_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1553_index_0_rename_ack_0 <= array_obj_ref_1553_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1552_resized;
      simple_obj_ref_1552_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1557_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1557_index_0_rename_ack_0 <= array_obj_ref_1557_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1556_resized;
      simple_obj_ref_1556_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1687_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1687_index_0_rename_ack_0 <= array_obj_ref_1687_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1686_resized;
      simple_obj_ref_1686_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1711_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1711_index_0_rename_ack_0 <= array_obj_ref_1711_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1710_resized;
      simple_obj_ref_1710_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1735_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1735_index_0_rename_ack_0 <= array_obj_ref_1735_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1734_resized;
      simple_obj_ref_1734_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1759_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1759_index_0_rename_ack_0 <= array_obj_ref_1759_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1758_resized;
      simple_obj_ref_1758_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1783_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1783_index_0_rename_ack_0 <= array_obj_ref_1783_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1782_resized;
      simple_obj_ref_1782_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1807_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1807_index_0_rename_ack_0 <= array_obj_ref_1807_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1806_resized;
      simple_obj_ref_1806_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1831_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1831_index_0_rename_ack_0 <= array_obj_ref_1831_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1830_resized;
      simple_obj_ref_1830_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_1849_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_1849_index_0_rename_ack_0 <= array_obj_ref_1849_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1848_resized;
      simple_obj_ref_1848_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1232_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1232_gather_scatter_ack_0 <= ptr_deref_1232_gather_scatter_req_0;
      aggregated_sig <= type_cast_1234_wire_constant;
      ptr_deref_1232_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1388_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1388_addr_0_ack_0 <= ptr_deref_1388_addr_0_req_0;
      aggregated_sig <= ptr_deref_1388_root_address;
      ptr_deref_1388_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1388_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1388_gather_scatter_ack_0 <= ptr_deref_1388_gather_scatter_req_0;
      aggregated_sig <= tmp2_1386;
      ptr_deref_1388_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1388_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1388_root_address_inst_ack_0 <= ptr_deref_1388_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1388_resized_base_address;
      ptr_deref_1388_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1402_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1402_addr_0_ack_0 <= ptr_deref_1402_addr_0_req_0;
      aggregated_sig <= ptr_deref_1402_root_address;
      ptr_deref_1402_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1402_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1402_gather_scatter_ack_0 <= ptr_deref_1402_gather_scatter_req_0;
      aggregated_sig <= tmp5_1400;
      ptr_deref_1402_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1402_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1402_root_address_inst_ack_0 <= ptr_deref_1402_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1402_resized_base_address;
      ptr_deref_1402_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1416_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1416_addr_0_ack_0 <= ptr_deref_1416_addr_0_req_0;
      aggregated_sig <= ptr_deref_1416_root_address;
      ptr_deref_1416_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1416_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1416_gather_scatter_ack_0 <= ptr_deref_1416_gather_scatter_req_0;
      aggregated_sig <= tmp8_1414;
      ptr_deref_1416_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1416_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1416_root_address_inst_ack_0 <= ptr_deref_1416_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1416_resized_base_address;
      ptr_deref_1416_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1430_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1430_addr_0_ack_0 <= ptr_deref_1430_addr_0_req_0;
      aggregated_sig <= ptr_deref_1430_root_address;
      ptr_deref_1430_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1430_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1430_gather_scatter_ack_0 <= ptr_deref_1430_gather_scatter_req_0;
      aggregated_sig <= tmp11_1428;
      ptr_deref_1430_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1430_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1430_root_address_inst_ack_0 <= ptr_deref_1430_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1430_resized_base_address;
      ptr_deref_1430_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1444_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1444_addr_0_ack_0 <= ptr_deref_1444_addr_0_req_0;
      aggregated_sig <= ptr_deref_1444_root_address;
      ptr_deref_1444_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1444_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1444_gather_scatter_ack_0 <= ptr_deref_1444_gather_scatter_req_0;
      aggregated_sig <= tmp14_1442;
      ptr_deref_1444_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1444_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1444_root_address_inst_ack_0 <= ptr_deref_1444_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1444_resized_base_address;
      ptr_deref_1444_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1458_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1458_addr_0_ack_0 <= ptr_deref_1458_addr_0_req_0;
      aggregated_sig <= ptr_deref_1458_root_address;
      ptr_deref_1458_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1458_gather_scatter_ack_0 <= ptr_deref_1458_gather_scatter_req_0;
      aggregated_sig <= tmp17_1456;
      ptr_deref_1458_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1458_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1458_root_address_inst_ack_0 <= ptr_deref_1458_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1458_resized_base_address;
      ptr_deref_1458_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1472_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1472_addr_0_ack_0 <= ptr_deref_1472_addr_0_req_0;
      aggregated_sig <= ptr_deref_1472_root_address;
      ptr_deref_1472_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1472_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1472_gather_scatter_ack_0 <= ptr_deref_1472_gather_scatter_req_0;
      aggregated_sig <= tmp20_1470;
      ptr_deref_1472_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1472_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1472_root_address_inst_ack_0 <= ptr_deref_1472_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1472_resized_base_address;
      ptr_deref_1472_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1480_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1480_addr_0_ack_0 <= ptr_deref_1480_addr_0_req_0;
      aggregated_sig <= ptr_deref_1480_root_address;
      ptr_deref_1480_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1480_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1480_gather_scatter_ack_0 <= ptr_deref_1480_gather_scatter_req_0;
      aggregated_sig <= tmp22_1478;
      ptr_deref_1480_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1480_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1480_root_address_inst_ack_0 <= ptr_deref_1480_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1480_resized_base_address;
      ptr_deref_1480_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1570_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1570_addr_0_ack_0 <= ptr_deref_1570_addr_0_req_0;
      aggregated_sig <= ptr_deref_1570_root_address;
      ptr_deref_1570_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1570_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1570_gather_scatter_ack_0 <= ptr_deref_1570_gather_scatter_req_0;
      aggregated_sig <= tmp25_1568;
      ptr_deref_1570_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1570_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1570_root_address_inst_ack_0 <= ptr_deref_1570_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1570_resized_base_address;
      ptr_deref_1570_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1584_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1584_addr_0_ack_0 <= ptr_deref_1584_addr_0_req_0;
      aggregated_sig <= ptr_deref_1584_root_address;
      ptr_deref_1584_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1584_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1584_gather_scatter_ack_0 <= ptr_deref_1584_gather_scatter_req_0;
      aggregated_sig <= tmp28_1582;
      ptr_deref_1584_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1584_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1584_root_address_inst_ack_0 <= ptr_deref_1584_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1584_resized_base_address;
      ptr_deref_1584_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1598_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1598_addr_0_ack_0 <= ptr_deref_1598_addr_0_req_0;
      aggregated_sig <= ptr_deref_1598_root_address;
      ptr_deref_1598_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1598_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1598_gather_scatter_ack_0 <= ptr_deref_1598_gather_scatter_req_0;
      aggregated_sig <= tmp31_1596;
      ptr_deref_1598_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1598_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1598_root_address_inst_ack_0 <= ptr_deref_1598_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1598_resized_base_address;
      ptr_deref_1598_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1612_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1612_addr_0_ack_0 <= ptr_deref_1612_addr_0_req_0;
      aggregated_sig <= ptr_deref_1612_root_address;
      ptr_deref_1612_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1612_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1612_gather_scatter_ack_0 <= ptr_deref_1612_gather_scatter_req_0;
      aggregated_sig <= tmp34_1610;
      ptr_deref_1612_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1612_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1612_root_address_inst_ack_0 <= ptr_deref_1612_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1612_resized_base_address;
      ptr_deref_1612_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1626_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1626_addr_0_ack_0 <= ptr_deref_1626_addr_0_req_0;
      aggregated_sig <= ptr_deref_1626_root_address;
      ptr_deref_1626_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1626_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1626_gather_scatter_ack_0 <= ptr_deref_1626_gather_scatter_req_0;
      aggregated_sig <= tmp37_1624;
      ptr_deref_1626_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1626_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1626_root_address_inst_ack_0 <= ptr_deref_1626_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1626_resized_base_address;
      ptr_deref_1626_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1640_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1640_addr_0_ack_0 <= ptr_deref_1640_addr_0_req_0;
      aggregated_sig <= ptr_deref_1640_root_address;
      ptr_deref_1640_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1640_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1640_gather_scatter_ack_0 <= ptr_deref_1640_gather_scatter_req_0;
      aggregated_sig <= tmp40_1638;
      ptr_deref_1640_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1640_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1640_root_address_inst_ack_0 <= ptr_deref_1640_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1640_resized_base_address;
      ptr_deref_1640_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1654_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1654_addr_0_ack_0 <= ptr_deref_1654_addr_0_req_0;
      aggregated_sig <= ptr_deref_1654_root_address;
      ptr_deref_1654_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1654_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1654_gather_scatter_ack_0 <= ptr_deref_1654_gather_scatter_req_0;
      aggregated_sig <= tmp43_1652;
      ptr_deref_1654_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1654_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1654_root_address_inst_ack_0 <= ptr_deref_1654_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1654_resized_base_address;
      ptr_deref_1654_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1662_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1662_addr_0_ack_0 <= ptr_deref_1662_addr_0_req_0;
      aggregated_sig <= ptr_deref_1662_root_address;
      ptr_deref_1662_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1662_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1662_gather_scatter_ack_0 <= ptr_deref_1662_gather_scatter_req_0;
      aggregated_sig <= tmp45_1660;
      ptr_deref_1662_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1662_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1662_root_address_inst_ack_0 <= ptr_deref_1662_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1662_resized_base_address;
      ptr_deref_1662_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1690_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1690_addr_0_ack_0 <= ptr_deref_1690_addr_0_req_0;
      aggregated_sig <= ptr_deref_1690_root_address;
      ptr_deref_1690_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1690_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1690_gather_scatter_ack_0 <= ptr_deref_1690_gather_scatter_req_0;
      aggregated_sig <= tmp48_1684;
      ptr_deref_1690_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1690_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1690_root_address_inst_ack_0 <= ptr_deref_1690_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1690_resized_base_address;
      ptr_deref_1690_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1714_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1714_addr_0_ack_0 <= ptr_deref_1714_addr_0_req_0;
      aggregated_sig <= ptr_deref_1714_root_address;
      ptr_deref_1714_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1714_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1714_gather_scatter_ack_0 <= ptr_deref_1714_gather_scatter_req_0;
      aggregated_sig <= tmp51_1702;
      ptr_deref_1714_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1714_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1714_root_address_inst_ack_0 <= ptr_deref_1714_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1714_resized_base_address;
      ptr_deref_1714_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1738_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1738_addr_0_ack_0 <= ptr_deref_1738_addr_0_req_0;
      aggregated_sig <= ptr_deref_1738_root_address;
      ptr_deref_1738_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1738_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1738_gather_scatter_ack_0 <= ptr_deref_1738_gather_scatter_req_0;
      aggregated_sig <= tmp54_1726;
      ptr_deref_1738_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1738_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1738_root_address_inst_ack_0 <= ptr_deref_1738_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1738_resized_base_address;
      ptr_deref_1738_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1762_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1762_addr_0_ack_0 <= ptr_deref_1762_addr_0_req_0;
      aggregated_sig <= ptr_deref_1762_root_address;
      ptr_deref_1762_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1762_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1762_gather_scatter_ack_0 <= ptr_deref_1762_gather_scatter_req_0;
      aggregated_sig <= tmp57_1750;
      ptr_deref_1762_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1762_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1762_root_address_inst_ack_0 <= ptr_deref_1762_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1762_resized_base_address;
      ptr_deref_1762_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1786_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1786_addr_0_ack_0 <= ptr_deref_1786_addr_0_req_0;
      aggregated_sig <= ptr_deref_1786_root_address;
      ptr_deref_1786_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1786_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1786_gather_scatter_ack_0 <= ptr_deref_1786_gather_scatter_req_0;
      aggregated_sig <= tmp60_1774;
      ptr_deref_1786_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1786_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1786_root_address_inst_ack_0 <= ptr_deref_1786_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1786_resized_base_address;
      ptr_deref_1786_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1810_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1810_addr_0_ack_0 <= ptr_deref_1810_addr_0_req_0;
      aggregated_sig <= ptr_deref_1810_root_address;
      ptr_deref_1810_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1810_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1810_gather_scatter_ack_0 <= ptr_deref_1810_gather_scatter_req_0;
      aggregated_sig <= tmp63_1798;
      ptr_deref_1810_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1810_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1810_root_address_inst_ack_0 <= ptr_deref_1810_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1810_resized_base_address;
      ptr_deref_1810_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1834_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1834_addr_0_ack_0 <= ptr_deref_1834_addr_0_req_0;
      aggregated_sig <= ptr_deref_1834_root_address;
      ptr_deref_1834_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1834_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1834_gather_scatter_ack_0 <= ptr_deref_1834_gather_scatter_req_0;
      aggregated_sig <= tmp66_1822;
      ptr_deref_1834_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1834_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1834_root_address_inst_ack_0 <= ptr_deref_1834_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1834_resized_base_address;
      ptr_deref_1834_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1852_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1852_addr_0_ack_0 <= ptr_deref_1852_addr_0_req_0;
      aggregated_sig <= ptr_deref_1852_root_address;
      ptr_deref_1852_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1852_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1852_gather_scatter_ack_0 <= ptr_deref_1852_gather_scatter_req_0;
      aggregated_sig <= tmp68_1840;
      ptr_deref_1852_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1852_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1852_root_address_inst_ack_0 <= ptr_deref_1852_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1852_resized_base_address;
      ptr_deref_1852_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_1263_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp2x_xi_1262;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1263_branch_req_0,
          ack0 => if_stmt_1263_branch_ack_0,
          ack1 => if_stmt_1263_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1366_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1368_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1366_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_1366_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1366_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_1371_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1366_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_1366_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_1366_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(1 downto 0);
      begin 
      condition_sig <= expr_1368_wire_constant_cmp & expr_1371_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 2)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_1366_branch_default_req_0,
          ack0 => switch_stmt_1366_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1292_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1292_resized_base_address;
      array_obj_ref_1292_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1292_root_address_inst_req_0,
          ackL => array_obj_ref_1292_root_address_inst_ack_0,
          reqR => array_obj_ref_1292_root_address_inst_req_1,
          ackR => array_obj_ref_1292_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1297_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1297_resized_base_address;
      array_obj_ref_1297_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1297_root_address_inst_req_0,
          ackL => array_obj_ref_1297_root_address_inst_ack_0,
          reqR => array_obj_ref_1297_root_address_inst_req_1,
          ackR => array_obj_ref_1297_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1302_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1302_resized_base_address;
      array_obj_ref_1302_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1302_root_address_inst_req_0,
          ackL => array_obj_ref_1302_root_address_inst_ack_0,
          reqR => array_obj_ref_1302_root_address_inst_req_1,
          ackR => array_obj_ref_1302_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1307_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1307_resized_base_address;
      array_obj_ref_1307_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1307_root_address_inst_req_0,
          ackL => array_obj_ref_1307_root_address_inst_ack_0,
          reqR => array_obj_ref_1307_root_address_inst_req_1,
          ackR => array_obj_ref_1307_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1316_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1316_resized_base_address;
      array_obj_ref_1316_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1316_root_address_inst_req_0,
          ackL => array_obj_ref_1316_root_address_inst_ack_0,
          reqR => array_obj_ref_1316_root_address_inst_req_1,
          ackR => array_obj_ref_1316_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1321_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1321_resized_base_address;
      array_obj_ref_1321_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1321_root_address_inst_req_0,
          ackL => array_obj_ref_1321_root_address_inst_ack_0,
          reqR => array_obj_ref_1321_root_address_inst_req_1,
          ackR => array_obj_ref_1321_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1326_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1326_resized_base_address;
      array_obj_ref_1326_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1326_root_address_inst_req_0,
          ackL => array_obj_ref_1326_root_address_inst_ack_0,
          reqR => array_obj_ref_1326_root_address_inst_req_1,
          ackR => array_obj_ref_1326_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1529_root_address_inst array_obj_ref_1687_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1529_final_offset & array_obj_ref_1529_resized_base_address & array_obj_ref_1687_final_offset & array_obj_ref_1687_resized_base_address;
      array_obj_ref_1529_root_address <= data_out(21 downto 11);
      array_obj_ref_1687_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1529_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1687_root_address_inst_req_0;
      array_obj_ref_1529_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1687_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1529_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1687_root_address_inst_req_1;
      array_obj_ref_1529_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1687_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1533_root_address_inst array_obj_ref_1711_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1533_final_offset & array_obj_ref_1533_resized_base_address & array_obj_ref_1711_final_offset & array_obj_ref_1711_resized_base_address;
      array_obj_ref_1533_root_address <= data_out(21 downto 11);
      array_obj_ref_1711_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1533_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1711_root_address_inst_req_0;
      array_obj_ref_1533_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1711_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1533_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1711_root_address_inst_req_1;
      array_obj_ref_1533_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1711_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1537_root_address_inst array_obj_ref_1735_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1537_final_offset & array_obj_ref_1537_resized_base_address & array_obj_ref_1735_final_offset & array_obj_ref_1735_resized_base_address;
      array_obj_ref_1537_root_address <= data_out(21 downto 11);
      array_obj_ref_1735_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1537_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1735_root_address_inst_req_0;
      array_obj_ref_1537_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1735_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1537_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1735_root_address_inst_req_1;
      array_obj_ref_1537_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1735_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1541_root_address_inst array_obj_ref_1759_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1541_final_offset & array_obj_ref_1541_resized_base_address & array_obj_ref_1759_final_offset & array_obj_ref_1759_resized_base_address;
      array_obj_ref_1541_root_address <= data_out(21 downto 11);
      array_obj_ref_1759_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1541_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1759_root_address_inst_req_0;
      array_obj_ref_1541_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1759_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1541_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1759_root_address_inst_req_1;
      array_obj_ref_1541_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1759_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1545_root_address_inst array_obj_ref_1783_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1545_final_offset & array_obj_ref_1545_resized_base_address & array_obj_ref_1783_final_offset & array_obj_ref_1783_resized_base_address;
      array_obj_ref_1545_root_address <= data_out(21 downto 11);
      array_obj_ref_1783_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1545_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1783_root_address_inst_req_0;
      array_obj_ref_1545_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1783_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1545_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1783_root_address_inst_req_1;
      array_obj_ref_1545_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1783_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1549_root_address_inst array_obj_ref_1807_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1549_final_offset & array_obj_ref_1549_resized_base_address & array_obj_ref_1807_final_offset & array_obj_ref_1807_resized_base_address;
      array_obj_ref_1549_root_address <= data_out(21 downto 11);
      array_obj_ref_1807_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1549_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1807_root_address_inst_req_0;
      array_obj_ref_1549_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1807_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1549_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1807_root_address_inst_req_1;
      array_obj_ref_1549_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1807_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_1553_root_address_inst array_obj_ref_1831_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1553_final_offset & array_obj_ref_1553_resized_base_address & array_obj_ref_1831_final_offset & array_obj_ref_1831_resized_base_address;
      array_obj_ref_1553_root_address <= data_out(21 downto 11);
      array_obj_ref_1831_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1553_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1831_root_address_inst_req_0;
      array_obj_ref_1553_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1831_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1553_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1831_root_address_inst_req_1;
      array_obj_ref_1553_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1831_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_1557_root_address_inst array_obj_ref_1849_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(43 downto 0);
      signal data_out: std_logic_vector(21 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1557_final_offset & array_obj_ref_1557_resized_base_address & array_obj_ref_1849_final_offset & array_obj_ref_1849_resized_base_address;
      array_obj_ref_1557_root_address <= data_out(21 downto 11);
      array_obj_ref_1849_root_address <= data_out(10 downto 0);
      reqL(1) <= array_obj_ref_1557_root_address_inst_req_0;
      reqL(0) <= array_obj_ref_1849_root_address_inst_req_0;
      array_obj_ref_1557_root_address_inst_ack_0 <= ackL(1);
      array_obj_ref_1849_root_address_inst_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1557_root_address_inst_req_1;
      reqR(0) <= array_obj_ref_1849_root_address_inst_req_1;
      array_obj_ref_1557_root_address_inst_ack_1 <= ackR(1);
      array_obj_ref_1849_root_address_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1261_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xi_1256;
      tmp2x_xi_1262 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1261_inst_req_0,
          ackL => binary_1261_inst_ack_0,
          reqR => binary_1261_inst_req_1,
          ackR => binary_1261_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1342_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_1330;
      tmp_1343 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1342_inst_req_0,
          ackL => binary_1342_inst_ack_0,
          reqR => binary_1342_inst_req_1,
          ackR => binary_1342_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1381_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp1_1382 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1381_inst_req_0,
          ackL => binary_1381_inst_ack_0,
          reqR => binary_1381_inst_req_1,
          ackR => binary_1381_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1395_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp4_1396 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1395_inst_req_0,
          ackL => binary_1395_inst_ack_0,
          reqR => binary_1395_inst_req_1,
          ackR => binary_1395_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1409_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp7_1410 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1409_inst_req_0,
          ackL => binary_1409_inst_ack_0,
          reqR => binary_1409_inst_req_1,
          ackR => binary_1409_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1423_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp10_1424 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1423_inst_req_0,
          ackL => binary_1423_inst_ack_0,
          reqR => binary_1423_inst_req_1,
          ackR => binary_1423_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1437_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp13_1438 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1437_inst_req_0,
          ackL => binary_1437_inst_ack_0,
          reqR => binary_1437_inst_req_1,
          ackR => binary_1437_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1451_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp16_1452 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1451_inst_req_0,
          ackL => binary_1451_inst_ack_0,
          reqR => binary_1451_inst_req_1,
          ackR => binary_1451_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1465_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp19_1466 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1465_inst_req_0,
          ackL => binary_1465_inst_ack_0,
          reqR => binary_1465_inst_req_1,
          ackR => binary_1465_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1489_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp142149_1490 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1489_inst_req_0,
          ackL => binary_1489_inst_ack_0,
          reqR => binary_1489_inst_req_1,
          ackR => binary_1489_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1495_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp141148_1496 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1495_inst_req_0,
          ackL => binary_1495_inst_ack_0,
          reqR => binary_1495_inst_req_1,
          ackR => binary_1495_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1501_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp140147_1502 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1501_inst_req_0,
          ackL => binary_1501_inst_ack_0,
          reqR => binary_1501_inst_req_1,
          ackR => binary_1501_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1507_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp139146_1508 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1507_inst_req_0,
          ackL => binary_1507_inst_ack_0,
          reqR => binary_1507_inst_req_1,
          ackR => binary_1507_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1513_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp138145_1514 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1513_inst_req_0,
          ackL => binary_1513_inst_ack_0,
          reqR => binary_1513_inst_req_1,
          ackR => binary_1513_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1519_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp137144_1520 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1519_inst_req_0,
          ackL => binary_1519_inst_ack_0,
          reqR => binary_1519_inst_req_1,
          ackR => binary_1519_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1525_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp136143_1526 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1525_inst_req_0,
          ackL => binary_1525_inst_ack_0,
          reqR => binary_1525_inst_req_1,
          ackR => binary_1525_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1563_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp24_1564 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1563_inst_req_0,
          ackL => binary_1563_inst_ack_0,
          reqR => binary_1563_inst_req_1,
          ackR => binary_1563_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1577_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp27_1578 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1577_inst_req_0,
          ackL => binary_1577_inst_ack_0,
          reqR => binary_1577_inst_req_1,
          ackR => binary_1577_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1591_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp30_1592 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1591_inst_req_0,
          ackL => binary_1591_inst_ack_0,
          reqR => binary_1591_inst_req_1,
          ackR => binary_1591_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1605_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp33_1606 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1605_inst_req_0,
          ackL => binary_1605_inst_ack_0,
          reqR => binary_1605_inst_req_1,
          ackR => binary_1605_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1619_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp36_1620 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1619_inst_req_0,
          ackL => binary_1619_inst_ack_0,
          reqR => binary_1619_inst_req_1,
          ackR => binary_1619_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1633_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp39_1634 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1633_inst_req_0,
          ackL => binary_1633_inst_ack_0,
          reqR => binary_1633_inst_req_1,
          ackR => binary_1633_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1647_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp42_1648 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1647_inst_req_0,
          ackL => binary_1647_inst_ack_0,
          reqR => binary_1647_inst_req_1,
          ackR => binary_1647_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_1671_inst binary_1859_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_9_1330 & iNsTr_9_1330;
      wordx_x0x_xbe_1672 <= data_out(63 downto 32);
      tmp134_1860 <= data_out(31 downto 0);
      reqL(1) <= binary_1671_inst_req_0;
      reqL(0) <= binary_1859_inst_req_0;
      binary_1671_inst_ack_0 <= ackL(1);
      binary_1859_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1671_inst_req_1;
      reqR(0) <= binary_1859_inst_req_1;
      binary_1671_inst_ack_1 <= ackR(1);
      binary_1859_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => true,
          min_clock_period => false,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_1679_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp47_1680 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1679_inst_req_0,
          ackL => binary_1679_inst_ack_0,
          reqR => binary_1679_inst_req_1,
          ackR => binary_1679_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_1697_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp50_1698 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1697_inst_req_0,
          ackL => binary_1697_inst_ack_0,
          reqR => binary_1697_inst_req_1,
          ackR => binary_1697_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_1707_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp114_1708 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1707_inst_req_0,
          ackL => binary_1707_inst_ack_0,
          reqR => binary_1707_inst_req_1,
          ackR => binary_1707_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_1721_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp53_1722 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1721_inst_req_0,
          ackL => binary_1721_inst_ack_0,
          reqR => binary_1721_inst_req_1,
          ackR => binary_1721_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_1731_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp117_1732 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1731_inst_req_0,
          ackL => binary_1731_inst_ack_0,
          reqR => binary_1731_inst_req_1,
          ackR => binary_1731_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_1745_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp56_1746 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1745_inst_req_0,
          ackL => binary_1745_inst_ack_0,
          reqR => binary_1745_inst_req_1,
          ackR => binary_1745_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_1755_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp120_1756 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1755_inst_req_0,
          ackL => binary_1755_inst_ack_0,
          reqR => binary_1755_inst_req_1,
          ackR => binary_1755_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_1769_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp59_1770 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1769_inst_req_0,
          ackL => binary_1769_inst_ack_0,
          reqR => binary_1769_inst_req_1,
          ackR => binary_1769_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_1779_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp123_1780 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1779_inst_req_0,
          ackL => binary_1779_inst_ack_0,
          reqR => binary_1779_inst_req_1,
          ackR => binary_1779_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_1793_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp62_1794 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1793_inst_req_0,
          ackL => binary_1793_inst_ack_0,
          reqR => binary_1793_inst_req_1,
          ackR => binary_1793_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_1803_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp126_1804 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1803_inst_req_0,
          ackL => binary_1803_inst_ack_0,
          reqR => binary_1803_inst_req_1,
          ackR => binary_1803_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_1817_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp72_1352;
      tmp65_1818 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1817_inst_req_0,
          ackL => binary_1817_inst_ack_0,
          reqR => binary_1817_inst_req_1,
          ackR => binary_1817_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_1827_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp129_1828 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1827_inst_req_0,
          ackL => binary_1827_inst_ack_0,
          reqR => binary_1827_inst_req_1,
          ackR => binary_1827_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_1845_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1343;
      tmp132_1846 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1845_inst_req_0,
          ackL => binary_1845_inst_ack_0,
          reqR => binary_1845_inst_req_1,
          ackR => binary_1845_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : switch_stmt_1366_select_expr_0 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1365;
      expr_1368_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000011111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1366_select_expr_0_req_0,
          ackL => switch_stmt_1366_select_expr_0_ack_0,
          reqR => switch_stmt_1366_select_expr_0_req_1,
          ackR => switch_stmt_1366_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : switch_stmt_1366_select_expr_1 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_1365;
      expr_1371_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_1366_select_expr_1_req_0,
          ackL => switch_stmt_1366_select_expr_1_ack_0,
          reqR => switch_stmt_1366_select_expr_1_req_1,
          ackR => switch_stmt_1366_select_expr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared store operator group (0) : ptr_deref_1232_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_1232_store_0_req_0;
      ptr_deref_1232_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_1232_store_0_req_1;
      ptr_deref_1232_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1232_word_address_0;
      data_in <= ptr_deref_1232_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 4,
        data_width => 8,
        num_reqs => 1,
        tag_length => 1,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(3 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(0 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared store operator group (1) : ptr_deref_1388_store_0 ptr_deref_1570_store_0 ptr_deref_1690_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1388_store_0_req_0;
      reqL(1) <= ptr_deref_1570_store_0_req_0;
      reqL(0) <= ptr_deref_1690_store_0_req_0;
      ptr_deref_1388_store_0_ack_0 <= ackL(2);
      ptr_deref_1570_store_0_ack_0 <= ackL(1);
      ptr_deref_1690_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1388_store_0_req_1;
      reqR(1) <= ptr_deref_1570_store_0_req_1;
      reqR(0) <= ptr_deref_1690_store_0_req_1;
      ptr_deref_1388_store_0_ack_1 <= ackR(2);
      ptr_deref_1570_store_0_ack_1 <= ackR(1);
      ptr_deref_1690_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1388_word_address_0 & ptr_deref_1570_word_address_0 & ptr_deref_1690_word_address_0;
      data_in <= ptr_deref_1388_data_0 & ptr_deref_1570_data_0 & ptr_deref_1690_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(7),
          mack => memory_space_3_sr_ack(7),
          maddr => memory_space_3_sr_addr(87 downto 77),
          mdata => memory_space_3_sr_data(63 downto 56),
          mtag => memory_space_3_sr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(7),
          mack => memory_space_3_sc_ack(7),
          mtag => memory_space_3_sc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared store operator group (2) : ptr_deref_1402_store_0 ptr_deref_1584_store_0 ptr_deref_1714_store_0 
    StoreGroup2: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1402_store_0_req_0;
      reqL(1) <= ptr_deref_1584_store_0_req_0;
      reqL(0) <= ptr_deref_1714_store_0_req_0;
      ptr_deref_1402_store_0_ack_0 <= ackL(2);
      ptr_deref_1584_store_0_ack_0 <= ackL(1);
      ptr_deref_1714_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1402_store_0_req_1;
      reqR(1) <= ptr_deref_1584_store_0_req_1;
      reqR(0) <= ptr_deref_1714_store_0_req_1;
      ptr_deref_1402_store_0_ack_1 <= ackR(2);
      ptr_deref_1584_store_0_ack_1 <= ackR(1);
      ptr_deref_1714_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1402_word_address_0 & ptr_deref_1584_word_address_0 & ptr_deref_1714_word_address_0;
      data_in <= ptr_deref_1402_data_0 & ptr_deref_1584_data_0 & ptr_deref_1714_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(6),
          mack => memory_space_3_sr_ack(6),
          maddr => memory_space_3_sr_addr(76 downto 66),
          mdata => memory_space_3_sr_data(55 downto 48),
          mtag => memory_space_3_sr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(6),
          mack => memory_space_3_sc_ack(6),
          mtag => memory_space_3_sc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 2
    -- shared store operator group (3) : ptr_deref_1416_store_0 ptr_deref_1598_store_0 ptr_deref_1738_store_0 
    StoreGroup3: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1416_store_0_req_0;
      reqL(1) <= ptr_deref_1598_store_0_req_0;
      reqL(0) <= ptr_deref_1738_store_0_req_0;
      ptr_deref_1416_store_0_ack_0 <= ackL(2);
      ptr_deref_1598_store_0_ack_0 <= ackL(1);
      ptr_deref_1738_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1416_store_0_req_1;
      reqR(1) <= ptr_deref_1598_store_0_req_1;
      reqR(0) <= ptr_deref_1738_store_0_req_1;
      ptr_deref_1416_store_0_ack_1 <= ackR(2);
      ptr_deref_1598_store_0_ack_1 <= ackR(1);
      ptr_deref_1738_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1416_word_address_0 & ptr_deref_1598_word_address_0 & ptr_deref_1738_word_address_0;
      data_in <= ptr_deref_1416_data_0 & ptr_deref_1598_data_0 & ptr_deref_1738_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(5),
          mack => memory_space_3_sr_ack(5),
          maddr => memory_space_3_sr_addr(65 downto 55),
          mdata => memory_space_3_sr_data(47 downto 40),
          mtag => memory_space_3_sr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(5),
          mack => memory_space_3_sc_ack(5),
          mtag => memory_space_3_sc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 3
    -- shared store operator group (4) : ptr_deref_1430_store_0 ptr_deref_1612_store_0 ptr_deref_1762_store_0 
    StoreGroup4: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1430_store_0_req_0;
      reqL(1) <= ptr_deref_1612_store_0_req_0;
      reqL(0) <= ptr_deref_1762_store_0_req_0;
      ptr_deref_1430_store_0_ack_0 <= ackL(2);
      ptr_deref_1612_store_0_ack_0 <= ackL(1);
      ptr_deref_1762_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1430_store_0_req_1;
      reqR(1) <= ptr_deref_1612_store_0_req_1;
      reqR(0) <= ptr_deref_1762_store_0_req_1;
      ptr_deref_1430_store_0_ack_1 <= ackR(2);
      ptr_deref_1612_store_0_ack_1 <= ackR(1);
      ptr_deref_1762_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1430_word_address_0 & ptr_deref_1612_word_address_0 & ptr_deref_1762_word_address_0;
      data_in <= ptr_deref_1430_data_0 & ptr_deref_1612_data_0 & ptr_deref_1762_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(4),
          mack => memory_space_3_sr_ack(4),
          maddr => memory_space_3_sr_addr(54 downto 44),
          mdata => memory_space_3_sr_data(39 downto 32),
          mtag => memory_space_3_sr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(4),
          mack => memory_space_3_sc_ack(4),
          mtag => memory_space_3_sc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 4
    -- shared store operator group (5) : ptr_deref_1444_store_0 ptr_deref_1626_store_0 ptr_deref_1786_store_0 
    StoreGroup5: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1444_store_0_req_0;
      reqL(1) <= ptr_deref_1626_store_0_req_0;
      reqL(0) <= ptr_deref_1786_store_0_req_0;
      ptr_deref_1444_store_0_ack_0 <= ackL(2);
      ptr_deref_1626_store_0_ack_0 <= ackL(1);
      ptr_deref_1786_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1444_store_0_req_1;
      reqR(1) <= ptr_deref_1626_store_0_req_1;
      reqR(0) <= ptr_deref_1786_store_0_req_1;
      ptr_deref_1444_store_0_ack_1 <= ackR(2);
      ptr_deref_1626_store_0_ack_1 <= ackR(1);
      ptr_deref_1786_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1444_word_address_0 & ptr_deref_1626_word_address_0 & ptr_deref_1786_word_address_0;
      data_in <= ptr_deref_1444_data_0 & ptr_deref_1626_data_0 & ptr_deref_1786_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(3),
          mack => memory_space_3_sr_ack(3),
          maddr => memory_space_3_sr_addr(43 downto 33),
          mdata => memory_space_3_sr_data(31 downto 24),
          mtag => memory_space_3_sr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(3),
          mack => memory_space_3_sc_ack(3),
          mtag => memory_space_3_sc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 5
    -- shared store operator group (6) : ptr_deref_1458_store_0 ptr_deref_1640_store_0 ptr_deref_1810_store_0 
    StoreGroup6: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1458_store_0_req_0;
      reqL(1) <= ptr_deref_1640_store_0_req_0;
      reqL(0) <= ptr_deref_1810_store_0_req_0;
      ptr_deref_1458_store_0_ack_0 <= ackL(2);
      ptr_deref_1640_store_0_ack_0 <= ackL(1);
      ptr_deref_1810_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1458_store_0_req_1;
      reqR(1) <= ptr_deref_1640_store_0_req_1;
      reqR(0) <= ptr_deref_1810_store_0_req_1;
      ptr_deref_1458_store_0_ack_1 <= ackR(2);
      ptr_deref_1640_store_0_ack_1 <= ackR(1);
      ptr_deref_1810_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1458_word_address_0 & ptr_deref_1640_word_address_0 & ptr_deref_1810_word_address_0;
      data_in <= ptr_deref_1458_data_0 & ptr_deref_1640_data_0 & ptr_deref_1810_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(2),
          mack => memory_space_3_sr_ack(2),
          maddr => memory_space_3_sr_addr(32 downto 22),
          mdata => memory_space_3_sr_data(23 downto 16),
          mtag => memory_space_3_sr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(2),
          mack => memory_space_3_sc_ack(2),
          mtag => memory_space_3_sc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 6
    -- shared store operator group (7) : ptr_deref_1472_store_0 ptr_deref_1654_store_0 ptr_deref_1834_store_0 
    StoreGroup7: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1472_store_0_req_0;
      reqL(1) <= ptr_deref_1654_store_0_req_0;
      reqL(0) <= ptr_deref_1834_store_0_req_0;
      ptr_deref_1472_store_0_ack_0 <= ackL(2);
      ptr_deref_1654_store_0_ack_0 <= ackL(1);
      ptr_deref_1834_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1472_store_0_req_1;
      reqR(1) <= ptr_deref_1654_store_0_req_1;
      reqR(0) <= ptr_deref_1834_store_0_req_1;
      ptr_deref_1472_store_0_ack_1 <= ackR(2);
      ptr_deref_1654_store_0_ack_1 <= ackR(1);
      ptr_deref_1834_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1472_word_address_0 & ptr_deref_1654_word_address_0 & ptr_deref_1834_word_address_0;
      data_in <= ptr_deref_1472_data_0 & ptr_deref_1654_data_0 & ptr_deref_1834_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(1),
          mack => memory_space_3_sr_ack(1),
          maddr => memory_space_3_sr_addr(21 downto 11),
          mdata => memory_space_3_sr_data(15 downto 8),
          mtag => memory_space_3_sr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(1),
          mack => memory_space_3_sc_ack(1),
          mtag => memory_space_3_sc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 7
    -- shared store operator group (8) : ptr_deref_1480_store_0 ptr_deref_1662_store_0 ptr_deref_1852_store_0 
    StoreGroup8: Block -- 
      signal addr_in: std_logic_vector(32 downto 0);
      signal data_in: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= ptr_deref_1480_store_0_req_0;
      reqL(1) <= ptr_deref_1662_store_0_req_0;
      reqL(0) <= ptr_deref_1852_store_0_req_0;
      ptr_deref_1480_store_0_ack_0 <= ackL(2);
      ptr_deref_1662_store_0_ack_0 <= ackL(1);
      ptr_deref_1852_store_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1480_store_0_req_1;
      reqR(1) <= ptr_deref_1662_store_0_req_1;
      reqR(0) <= ptr_deref_1852_store_0_req_1;
      ptr_deref_1480_store_0_ack_1 <= ackR(2);
      ptr_deref_1662_store_0_ack_1 <= ackR(1);
      ptr_deref_1852_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1480_word_address_0 & ptr_deref_1662_word_address_0 & ptr_deref_1852_word_address_0;
      data_in <= ptr_deref_1480_data_0 & ptr_deref_1662_data_0 & ptr_deref_1852_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 11,
        data_width => 8,
        num_reqs => 3,
        tag_length => 2,
        min_clock_period => false,
        no_arbitration => true)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(10 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 3,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 8
    -- shared inport operator group (0) : simple_obj_ref_1255_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1255_inst_req_0;
      simple_obj_ref_1255_inst_ack_0 <= ack(0);
      tmpx_xi_1256 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_ack_pipe_read_req(0),
          oack => free_queue_ack_pipe_read_ack(0),
          odata => free_queue_ack_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1277_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1277_inst_req_0;
      simple_obj_ref_1277_inst_ack_0 <= ack(0);
      tmp4x_xi_1278 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_get_pipe_read_req(0),
          oack => free_queue_get_pipe_read_ack(0),
          odata => free_queue_get_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_1351_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1351_inst_req_0;
      simple_obj_ref_1351_inst_ack_0 <= ack(0);
      tmp72_1352 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_1360_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1360_inst_req_0;
      simple_obj_ref_1360_inst_ack_0 <= ack(0);
      tmp73_1361 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_ctrl_pipe_read_req(0),
          oack => in_ctrl_pipe_read_ack(0),
          odata => in_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared outport operator group (0) : simple_obj_ref_1244_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1244_inst_req_0;
      simple_obj_ref_1244_inst_ack_0 <= ack(0);
      data_in <= type_cast_1246_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_1867_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1867_inst_req_0;
      simple_obj_ref_1867_inst_ack_0 <= ack(0);
      data_in <= tmp4x_xi_1278;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => midpipe_pipe_write_req(0),
          oack => midpipe_pipe_write_ack(0),
          odata => midpipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_1876_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1876_inst_req_0;
      simple_obj_ref_1876_inst_ack_0 <= ack(0);
      data_in <= tmp73_1361;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => last_ctrl_pipe_write_req(0),
          oack => last_ctrl_pipe_write_ack(0),
          odata => last_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_1885_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1885_inst_req_0;
      simple_obj_ref_1885_inst_ack_0 <= ack(0);
      data_in <= tmp134_1860;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => pkt_length_pipe_write_req(0),
          oack => pkt_length_pipe_write_ack(0),
          odata => pkt_length_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_3_lr_req : out  std_logic_vector(7 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(87 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(15 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(7 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(7 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(15 downto 0);
    midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    last_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    last_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    last_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    pkt_length_pipe_read_req : out  std_logic_vector(0 downto 0);
    pkt_length_pipe_read_ack : in   std_logic_vector(0 downto 0);
    pkt_length_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
    free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
    op_lut_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    op_lut_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    op_lut_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    op_lut_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    op_lut_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_output;
architecture Default of wrapper_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_output_CP_8674_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_1965_gather_scatter_req_0 : boolean;
  signal binary_2013_inst_ack_0 : boolean;
  signal ptr_deref_1965_base_resize_req_0 : boolean;
  signal array_obj_ref_2275_base_resize_ack_0 : boolean;
  signal binary_2013_inst_req_0 : boolean;
  signal ptr_deref_2003_addr_0_req_0 : boolean;
  signal array_obj_ref_1999_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2003_base_resize_req_0 : boolean;
  signal binary_2013_inst_req_1 : boolean;
  signal array_obj_ref_2018_base_resize_ack_0 : boolean;
  signal ptr_deref_2036_load_0_req_0 : boolean;
  signal binary_1975_inst_ack_1 : boolean;
  signal array_obj_ref_2051_root_address_inst_ack_1 : boolean;
  signal binary_2013_inst_ack_1 : boolean;
  signal ptr_deref_2022_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1980_base_resize_ack_0 : boolean;
  signal binary_2032_inst_ack_0 : boolean;
  signal array_obj_ref_2275_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2022_load_0_req_1 : boolean;
  signal array_obj_ref_2018_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2018_base_resize_req_0 : boolean;
  signal type_cast_2007_inst_req_0 : boolean;
  signal ptr_deref_2055_root_address_inst_ack_0 : boolean;
  signal binary_1994_inst_ack_0 : boolean;
  signal binary_1994_inst_ack_1 : boolean;
  signal ptr_deref_1965_base_resize_ack_0 : boolean;
  signal array_obj_ref_1999_base_resize_ack_0 : boolean;
  signal array_obj_ref_1999_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1999_root_address_inst_ack_1 : boolean;
  signal type_cast_2007_inst_ack_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1980_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1999_base_resize_req_0 : boolean;
  signal ptr_deref_1965_load_0_ack_1 : boolean;
  signal ptr_deref_2022_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2036_root_address_inst_req_0 : boolean;
  signal ptr_deref_2022_load_0_ack_1 : boolean;
  signal ptr_deref_1965_load_0_req_1 : boolean;
  signal binary_1975_inst_req_1 : boolean;
  signal array_obj_ref_1980_root_address_inst_req_1 : boolean;
  signal ptr_deref_2055_load_0_req_0 : boolean;
  signal type_cast_1988_inst_req_0 : boolean;
  signal array_obj_ref_2018_final_reg_req_0 : boolean;
  signal array_obj_ref_2203_base_resize_req_0 : boolean;
  signal ptr_deref_2022_base_resize_req_0 : boolean;
  signal ptr_deref_1965_addr_0_ack_0 : boolean;
  signal binary_2032_inst_req_1 : boolean;
  signal ptr_deref_1984_gather_scatter_req_0 : boolean;
  signal ptr_deref_1965_root_address_inst_req_0 : boolean;
  signal ptr_deref_1984_gather_scatter_ack_0 : boolean;
  signal binary_2046_inst_ack_1 : boolean;
  signal array_obj_ref_1961_root_address_inst_req_1 : boolean;
  signal ptr_deref_1965_load_0_req_0 : boolean;
  signal type_cast_1988_inst_ack_0 : boolean;
  signal ptr_deref_1965_load_0_ack_0 : boolean;
  signal ptr_deref_1984_load_0_ack_1 : boolean;
  signal type_cast_2026_inst_ack_0 : boolean;
  signal ptr_deref_2022_load_0_req_0 : boolean;
  signal ptr_deref_2036_addr_0_ack_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_ack_1 : boolean;
  signal binary_1994_inst_req_1 : boolean;
  signal array_obj_ref_2051_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1980_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1980_root_address_inst_req_0 : boolean;
  signal ptr_deref_1965_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2051_final_reg_ack_0 : boolean;
  signal ptr_deref_2036_base_resize_req_0 : boolean;
  signal ptr_deref_1965_addr_0_req_0 : boolean;
  signal ptr_deref_2003_gather_scatter_req_0 : boolean;
  signal ptr_deref_2022_load_0_ack_0 : boolean;
  signal binary_1994_inst_req_0 : boolean;
  signal type_cast_2026_inst_req_0 : boolean;
  signal ptr_deref_2279_addr_0_req_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_req_1 : boolean;
  signal binary_1975_inst_ack_0 : boolean;
  signal ptr_deref_2055_base_resize_req_0 : boolean;
  signal binary_2032_inst_ack_1 : boolean;
  signal array_obj_ref_2203_base_resize_ack_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_req_0 : boolean;
  signal binary_2046_inst_ack_0 : boolean;
  signal binary_2046_inst_req_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1984_load_0_req_1 : boolean;
  signal array_obj_ref_1961_final_reg_req_0 : boolean;
  signal ptr_deref_2055_load_0_ack_1 : boolean;
  signal binary_1975_inst_req_0 : boolean;
  signal array_obj_ref_1961_final_reg_ack_0 : boolean;
  signal array_obj_ref_2018_root_address_inst_req_0 : boolean;
  signal binary_2046_inst_req_1 : boolean;
  signal ptr_deref_2003_gather_scatter_ack_0 : boolean;
  signal binary_2032_inst_req_0 : boolean;
  signal binary_2217_inst_ack_0 : boolean;
  signal ptr_deref_2036_load_0_ack_0 : boolean;
  signal array_obj_ref_1961_base_resize_ack_0 : boolean;
  signal array_obj_ref_1961_base_resize_req_0 : boolean;
  signal ptr_deref_2036_addr_0_req_0 : boolean;
  signal ptr_deref_1984_load_0_ack_0 : boolean;
  signal ptr_deref_1984_load_0_req_0 : boolean;
  signal array_obj_ref_2051_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2003_load_0_ack_1 : boolean;
  signal ptr_deref_2003_load_0_req_1 : boolean;
  signal binary_2217_inst_req_0 : boolean;
  signal array_obj_ref_2051_root_address_inst_req_0 : boolean;
  signal ptr_deref_2279_load_0_req_0 : boolean;
  signal ptr_deref_2279_base_resize_ack_0 : boolean;
  signal ptr_deref_1984_addr_0_ack_0 : boolean;
  signal type_cast_2040_inst_ack_0 : boolean;
  signal type_cast_2040_inst_req_0 : boolean;
  signal ptr_deref_2055_addr_0_ack_0 : boolean;
  signal type_cast_2235_inst_req_0 : boolean;
  signal ptr_deref_1984_addr_0_req_0 : boolean;
  signal array_obj_ref_1999_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1980_final_reg_ack_0 : boolean;
  signal binary_1956_inst_ack_1 : boolean;
  signal binary_1956_inst_req_1 : boolean;
  signal ptr_deref_2055_load_0_ack_0 : boolean;
  signal ptr_deref_1984_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1984_root_address_inst_req_0 : boolean;
  signal binary_1956_inst_ack_0 : boolean;
  signal ptr_deref_2231_load_0_req_1 : boolean;
  signal ptr_deref_1984_base_resize_ack_0 : boolean;
  signal ptr_deref_1984_base_resize_req_0 : boolean;
  signal binary_1956_inst_req_0 : boolean;
  signal ptr_deref_2022_addr_0_ack_0 : boolean;
  signal ptr_deref_2003_load_0_ack_0 : boolean;
  signal ptr_deref_2003_load_0_req_0 : boolean;
  signal ptr_deref_2055_root_address_inst_req_0 : boolean;
  signal ptr_deref_2022_base_resize_ack_0 : boolean;
  signal ptr_deref_2022_addr_0_req_0 : boolean;
  signal ptr_deref_2036_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2036_gather_scatter_req_0 : boolean;
  signal array_obj_ref_2051_base_resize_ack_0 : boolean;
  signal binary_2271_inst_req_0 : boolean;
  signal ptr_deref_2036_load_0_ack_1 : boolean;
  signal array_obj_ref_2203_root_address_inst_ack_1 : boolean;
  signal binary_2289_inst_ack_1 : boolean;
  signal binary_2289_inst_req_1 : boolean;
  signal binary_2070_inst_req_0 : boolean;
  signal binary_2070_inst_ack_0 : boolean;
  signal type_cast_2259_inst_ack_0 : boolean;
  signal binary_2070_inst_req_1 : boolean;
  signal type_cast_2259_inst_req_0 : boolean;
  signal binary_2070_inst_ack_1 : boolean;
  signal ptr_deref_2231_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2231_root_address_inst_req_0 : boolean;
  signal binary_2289_inst_ack_0 : boolean;
  signal ptr_deref_2207_gather_scatter_ack_0 : boolean;
  signal binary_2295_inst_ack_1 : boolean;
  signal binary_2295_inst_req_1 : boolean;
  signal ptr_deref_2207_gather_scatter_req_0 : boolean;
  signal binary_2075_inst_req_0 : boolean;
  signal binary_2075_inst_ack_0 : boolean;
  signal binary_2075_inst_req_1 : boolean;
  signal binary_2075_inst_ack_1 : boolean;
  signal binary_2295_inst_ack_0 : boolean;
  signal ptr_deref_2207_load_0_ack_1 : boolean;
  signal ptr_deref_2255_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2231_base_resize_ack_0 : boolean;
  signal ptr_deref_2255_gather_scatter_req_0 : boolean;
  signal ptr_deref_2231_base_resize_req_0 : boolean;
  signal ptr_deref_2207_load_0_req_1 : boolean;
  signal binary_2289_inst_req_0 : boolean;
  signal binary_2295_inst_req_0 : boolean;
  signal ptr_deref_2255_load_0_ack_1 : boolean;
  signal binary_2080_inst_req_0 : boolean;
  signal ptr_deref_2255_load_0_req_1 : boolean;
  signal binary_2080_inst_ack_0 : boolean;
  signal binary_2080_inst_req_1 : boolean;
  signal array_obj_ref_2203_index_0_rename_ack_0 : boolean;
  signal binary_2080_inst_ack_1 : boolean;
  signal array_obj_ref_2275_final_reg_ack_0 : boolean;
  signal ptr_deref_2279_addr_0_ack_0 : boolean;
  signal array_obj_ref_2051_final_reg_req_0 : boolean;
  signal ptr_deref_2231_load_0_ack_0 : boolean;
  signal type_cast_2235_inst_ack_0 : boolean;
  signal array_obj_ref_2203_offset_inst_req_0 : boolean;
  signal binary_2065_inst_ack_1 : boolean;
  signal ptr_deref_2231_addr_0_ack_0 : boolean;
  signal ptr_deref_2231_addr_0_req_0 : boolean;
  signal ptr_deref_2279_base_resize_req_0 : boolean;
  signal binary_2265_inst_req_0 : boolean;
  signal binary_2065_inst_req_0 : boolean;
  signal binary_2065_inst_ack_0 : boolean;
  signal binary_2065_inst_req_1 : boolean;
  signal ptr_deref_1965_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2022_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1980_base_resize_req_0 : boolean;
  signal binary_2265_inst_req_1 : boolean;
  signal ptr_deref_2055_addr_0_req_0 : boolean;
  signal ptr_deref_2003_addr_0_ack_0 : boolean;
  signal type_cast_1969_inst_req_0 : boolean;
  signal ptr_deref_2003_root_address_inst_req_0 : boolean;
  signal ptr_deref_2036_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2003_base_resize_ack_0 : boolean;
  signal ptr_deref_2055_gather_scatter_ack_0 : boolean;
  signal type_cast_2211_inst_ack_0 : boolean;
  signal binary_2265_inst_ack_0 : boolean;
  signal ptr_deref_2022_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2003_root_address_inst_ack_0 : boolean;
  signal type_cast_2059_inst_req_0 : boolean;
  signal binary_2265_inst_ack_1 : boolean;
  signal type_cast_2059_inst_ack_0 : boolean;
  signal ptr_deref_2231_load_0_req_0 : boolean;
  signal array_obj_ref_2203_offset_inst_ack_0 : boolean;
  signal ptr_deref_2055_load_0_req_1 : boolean;
  signal type_cast_2211_inst_req_0 : boolean;
  signal ptr_deref_2055_gather_scatter_req_0 : boolean;
  signal type_cast_2283_inst_req_0 : boolean;
  signal type_cast_1969_inst_ack_0 : boolean;
  signal simple_obj_ref_1902_inst_req_0 : boolean;
  signal simple_obj_ref_1902_inst_ack_0 : boolean;
  signal type_cast_1906_inst_req_0 : boolean;
  signal type_cast_1906_inst_ack_0 : boolean;
  signal array_obj_ref_1980_final_reg_req_0 : boolean;
  signal simple_obj_ref_1915_inst_req_0 : boolean;
  signal simple_obj_ref_1915_inst_ack_0 : boolean;
  signal array_obj_ref_1999_final_reg_ack_0 : boolean;
  signal array_obj_ref_1999_final_reg_req_0 : boolean;
  signal simple_obj_ref_1924_inst_req_0 : boolean;
  signal simple_obj_ref_1924_inst_ack_0 : boolean;
  signal array_obj_ref_1929_base_resize_req_0 : boolean;
  signal array_obj_ref_1929_base_resize_ack_0 : boolean;
  signal array_obj_ref_1929_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1929_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1929_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1929_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1929_final_reg_req_0 : boolean;
  signal array_obj_ref_1929_final_reg_ack_0 : boolean;
  signal binary_2241_inst_ack_0 : boolean;
  signal ptr_deref_1933_base_resize_req_0 : boolean;
  signal ptr_deref_1933_base_resize_ack_0 : boolean;
  signal ptr_deref_1933_root_address_inst_req_0 : boolean;
  signal ptr_deref_1933_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1933_addr_0_req_0 : boolean;
  signal ptr_deref_1933_addr_0_ack_0 : boolean;
  signal ptr_deref_2055_base_resize_ack_0 : boolean;
  signal ptr_deref_1933_load_0_req_0 : boolean;
  signal ptr_deref_1933_load_0_ack_0 : boolean;
  signal ptr_deref_1933_load_0_req_1 : boolean;
  signal ptr_deref_1933_load_0_ack_1 : boolean;
  signal array_obj_ref_2051_base_resize_req_0 : boolean;
  signal ptr_deref_1933_gather_scatter_req_0 : boolean;
  signal ptr_deref_1933_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2036_load_0_req_1 : boolean;
  signal array_obj_ref_2018_final_reg_ack_0 : boolean;
  signal ptr_deref_2036_base_resize_ack_0 : boolean;
  signal ptr_deref_2231_load_0_ack_1 : boolean;
  signal type_cast_1937_inst_req_0 : boolean;
  signal binary_2271_inst_ack_0 : boolean;
  signal type_cast_1937_inst_ack_0 : boolean;
  signal binary_2241_inst_req_0 : boolean;
  signal binary_2271_inst_req_1 : boolean;
  signal binary_2271_inst_ack_1 : boolean;
  signal binary_2217_inst_req_1 : boolean;
  signal ptr_deref_2231_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1942_base_resize_req_0 : boolean;
  signal array_obj_ref_1942_base_resize_ack_0 : boolean;
  signal binary_2217_inst_ack_1 : boolean;
  signal ptr_deref_2231_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1942_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1942_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1942_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1942_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1942_final_reg_req_0 : boolean;
  signal binary_2241_inst_req_1 : boolean;
  signal array_obj_ref_1942_final_reg_ack_0 : boolean;
  signal array_obj_ref_2203_root_address_inst_req_0 : boolean;
  signal binary_2241_inst_ack_1 : boolean;
  signal ptr_deref_1946_base_resize_req_0 : boolean;
  signal array_obj_ref_2203_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1946_base_resize_ack_0 : boolean;
  signal array_obj_ref_2203_root_address_inst_req_1 : boolean;
  signal ptr_deref_1946_root_address_inst_req_0 : boolean;
  signal ptr_deref_1946_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1946_addr_0_req_0 : boolean;
  signal ptr_deref_1946_addr_0_ack_0 : boolean;
  signal ptr_deref_1946_load_0_req_0 : boolean;
  signal ptr_deref_1946_load_0_ack_0 : boolean;
  signal ptr_deref_1946_load_0_req_1 : boolean;
  signal ptr_deref_1946_load_0_ack_1 : boolean;
  signal ptr_deref_1946_gather_scatter_req_0 : boolean;
  signal ptr_deref_1946_gather_scatter_ack_0 : boolean;
  signal type_cast_1950_inst_req_0 : boolean;
  signal type_cast_1950_inst_ack_0 : boolean;
  signal binary_2085_inst_req_0 : boolean;
  signal binary_2085_inst_ack_0 : boolean;
  signal binary_2085_inst_req_1 : boolean;
  signal array_obj_ref_2203_index_0_rename_req_0 : boolean;
  signal binary_2085_inst_ack_1 : boolean;
  signal array_obj_ref_2299_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2207_load_0_ack_0 : boolean;
  signal ptr_deref_2255_load_0_ack_0 : boolean;
  signal ptr_deref_2255_load_0_req_0 : boolean;
  signal ptr_deref_2207_load_0_req_0 : boolean;
  signal array_obj_ref_2275_final_reg_req_0 : boolean;
  signal binary_2090_inst_req_0 : boolean;
  signal binary_2090_inst_ack_0 : boolean;
  signal binary_2090_inst_req_1 : boolean;
  signal binary_2090_inst_ack_1 : boolean;
  signal array_obj_ref_2299_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2227_final_reg_ack_0 : boolean;
  signal ptr_deref_2279_gather_scatter_ack_0 : boolean;
  signal binary_2095_inst_req_0 : boolean;
  signal ptr_deref_2255_addr_0_ack_0 : boolean;
  signal binary_2095_inst_ack_0 : boolean;
  signal array_obj_ref_2227_final_reg_req_0 : boolean;
  signal ptr_deref_2255_addr_0_req_0 : boolean;
  signal binary_2095_inst_req_1 : boolean;
  signal binary_2095_inst_ack_1 : boolean;
  signal ptr_deref_2207_addr_0_ack_0 : boolean;
  signal ptr_deref_2255_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2227_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2207_addr_0_req_0 : boolean;
  signal ptr_deref_2279_gather_scatter_req_0 : boolean;
  signal ptr_deref_2255_root_address_inst_req_0 : boolean;
  signal binary_2100_inst_req_0 : boolean;
  signal binary_2100_inst_ack_0 : boolean;
  signal array_obj_ref_2227_root_address_inst_req_1 : boolean;
  signal binary_2100_inst_req_1 : boolean;
  signal array_obj_ref_2203_index_0_resize_ack_0 : boolean;
  signal binary_2100_inst_ack_1 : boolean;
  signal array_obj_ref_2275_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2227_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2255_base_resize_ack_0 : boolean;
  signal ptr_deref_2255_base_resize_req_0 : boolean;
  signal array_obj_ref_2227_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2203_index_0_resize_req_0 : boolean;
  signal simple_obj_ref_2108_inst_req_0 : boolean;
  signal simple_obj_ref_2108_inst_ack_0 : boolean;
  signal array_obj_ref_2275_base_resize_req_0 : boolean;
  signal ptr_deref_2279_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2279_load_0_ack_1 : boolean;
  signal ptr_deref_2207_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2227_base_resize_ack_0 : boolean;
  signal simple_obj_ref_2118_inst_req_0 : boolean;
  signal simple_obj_ref_2118_inst_ack_0 : boolean;
  signal array_obj_ref_2227_base_resize_req_0 : boolean;
  signal ptr_deref_2279_root_address_inst_req_0 : boolean;
  signal ptr_deref_2279_load_0_req_1 : boolean;
  signal array_obj_ref_2275_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2207_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2251_final_reg_ack_0 : boolean;
  signal binary_2125_inst_req_0 : boolean;
  signal array_obj_ref_2251_final_reg_req_0 : boolean;
  signal binary_2125_inst_ack_0 : boolean;
  signal binary_2125_inst_req_1 : boolean;
  signal binary_2125_inst_ack_1 : boolean;
  signal array_obj_ref_2251_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2227_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2251_root_address_inst_req_1 : boolean;
  signal type_cast_2283_inst_ack_0 : boolean;
  signal array_obj_ref_2275_root_address_inst_req_1 : boolean;
  signal ptr_deref_2207_base_resize_ack_0 : boolean;
  signal array_obj_ref_2251_root_address_inst_ack_0 : boolean;
  signal type_cast_2140_inst_req_0 : boolean;
  signal array_obj_ref_2251_root_address_inst_req_0 : boolean;
  signal type_cast_2140_inst_ack_0 : boolean;
  signal ptr_deref_2207_base_resize_req_0 : boolean;
  signal array_obj_ref_2227_offset_inst_req_0 : boolean;
  signal array_obj_ref_2227_index_0_rename_ack_0 : boolean;
  signal binary_2145_inst_req_0 : boolean;
  signal array_obj_ref_2251_base_resize_ack_0 : boolean;
  signal binary_2145_inst_ack_0 : boolean;
  signal array_obj_ref_2227_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2251_base_resize_req_0 : boolean;
  signal binary_2145_inst_req_1 : boolean;
  signal binary_2145_inst_ack_1 : boolean;
  signal array_obj_ref_2227_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2227_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2251_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2251_offset_inst_req_0 : boolean;
  signal binary_2151_inst_req_0 : boolean;
  signal binary_2151_inst_ack_0 : boolean;
  signal binary_2151_inst_req_1 : boolean;
  signal binary_2151_inst_ack_1 : boolean;
  signal array_obj_ref_2275_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2275_offset_inst_req_0 : boolean;
  signal array_obj_ref_2251_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2251_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2275_index_0_rename_ack_0 : boolean;
  signal binary_2157_inst_req_0 : boolean;
  signal binary_2157_inst_ack_0 : boolean;
  signal array_obj_ref_2251_index_0_resize_ack_0 : boolean;
  signal binary_2157_inst_req_1 : boolean;
  signal array_obj_ref_2251_index_0_resize_req_0 : boolean;
  signal binary_2157_inst_ack_1 : boolean;
  signal array_obj_ref_2275_index_0_rename_req_0 : boolean;
  signal binary_2223_inst_ack_1 : boolean;
  signal binary_2223_inst_req_1 : boolean;
  signal binary_2223_inst_ack_0 : boolean;
  signal binary_2223_inst_req_0 : boolean;
  signal array_obj_ref_2275_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2275_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2161_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2161_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2299_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2203_final_reg_ack_0 : boolean;
  signal array_obj_ref_2161_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2161_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2299_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2203_final_reg_req_0 : boolean;
  signal array_obj_ref_2161_offset_inst_req_0 : boolean;
  signal array_obj_ref_2161_offset_inst_ack_0 : boolean;
  signal binary_2247_inst_ack_1 : boolean;
  signal binary_2247_inst_req_1 : boolean;
  signal array_obj_ref_2161_base_resize_req_0 : boolean;
  signal binary_2247_inst_ack_0 : boolean;
  signal array_obj_ref_2161_base_resize_ack_0 : boolean;
  signal binary_2247_inst_req_0 : boolean;
  signal ptr_deref_2279_load_0_ack_0 : boolean;
  signal array_obj_ref_2161_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2161_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2161_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2161_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2161_final_reg_req_0 : boolean;
  signal array_obj_ref_2161_final_reg_ack_0 : boolean;
  signal ptr_deref_2165_base_resize_req_0 : boolean;
  signal ptr_deref_2165_base_resize_ack_0 : boolean;
  signal ptr_deref_2165_root_address_inst_req_0 : boolean;
  signal ptr_deref_2165_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2165_addr_0_req_0 : boolean;
  signal ptr_deref_2165_addr_0_ack_0 : boolean;
  signal ptr_deref_2165_load_0_req_0 : boolean;
  signal ptr_deref_2165_load_0_ack_0 : boolean;
  signal ptr_deref_2165_load_0_req_1 : boolean;
  signal ptr_deref_2165_load_0_ack_1 : boolean;
  signal ptr_deref_2165_gather_scatter_req_0 : boolean;
  signal ptr_deref_2165_gather_scatter_ack_0 : boolean;
  signal type_cast_2169_inst_req_0 : boolean;
  signal type_cast_2169_inst_ack_0 : boolean;
  signal binary_2175_inst_req_0 : boolean;
  signal binary_2175_inst_ack_0 : boolean;
  signal binary_2175_inst_req_1 : boolean;
  signal binary_2175_inst_ack_1 : boolean;
  signal array_obj_ref_2179_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2179_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2179_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2179_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2179_offset_inst_req_0 : boolean;
  signal array_obj_ref_2179_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2179_base_resize_req_0 : boolean;
  signal array_obj_ref_2179_base_resize_ack_0 : boolean;
  signal array_obj_ref_2179_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2179_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2179_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2179_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2179_final_reg_req_0 : boolean;
  signal array_obj_ref_2179_final_reg_ack_0 : boolean;
  signal ptr_deref_2183_base_resize_req_0 : boolean;
  signal ptr_deref_2183_base_resize_ack_0 : boolean;
  signal ptr_deref_2183_root_address_inst_req_0 : boolean;
  signal ptr_deref_2183_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2183_addr_0_req_0 : boolean;
  signal ptr_deref_2183_addr_0_ack_0 : boolean;
  signal ptr_deref_2183_load_0_req_0 : boolean;
  signal ptr_deref_2183_load_0_ack_0 : boolean;
  signal ptr_deref_2183_load_0_req_1 : boolean;
  signal ptr_deref_2183_load_0_ack_1 : boolean;
  signal ptr_deref_2183_gather_scatter_req_0 : boolean;
  signal ptr_deref_2183_gather_scatter_ack_0 : boolean;
  signal type_cast_2187_inst_req_0 : boolean;
  signal type_cast_2187_inst_ack_0 : boolean;
  signal binary_2193_inst_req_0 : boolean;
  signal binary_2193_inst_ack_0 : boolean;
  signal binary_2193_inst_req_1 : boolean;
  signal binary_2193_inst_ack_1 : boolean;
  signal binary_2199_inst_req_0 : boolean;
  signal binary_2199_inst_ack_0 : boolean;
  signal binary_2199_inst_req_1 : boolean;
  signal binary_2199_inst_ack_1 : boolean;
  signal array_obj_ref_2299_offset_inst_req_0 : boolean;
  signal array_obj_ref_2299_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2299_base_resize_req_0 : boolean;
  signal array_obj_ref_2299_base_resize_ack_0 : boolean;
  signal array_obj_ref_2299_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2299_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2299_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2299_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2299_final_reg_req_0 : boolean;
  signal array_obj_ref_2299_final_reg_ack_0 : boolean;
  signal ptr_deref_2303_base_resize_req_0 : boolean;
  signal ptr_deref_2303_base_resize_ack_0 : boolean;
  signal ptr_deref_2303_root_address_inst_req_0 : boolean;
  signal ptr_deref_2303_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2303_addr_0_req_0 : boolean;
  signal ptr_deref_2303_addr_0_ack_0 : boolean;
  signal ptr_deref_2303_load_0_req_0 : boolean;
  signal ptr_deref_2303_load_0_ack_0 : boolean;
  signal ptr_deref_2303_load_0_req_1 : boolean;
  signal ptr_deref_2303_load_0_ack_1 : boolean;
  signal ptr_deref_2303_gather_scatter_req_0 : boolean;
  signal ptr_deref_2303_gather_scatter_ack_0 : boolean;
  signal type_cast_2307_inst_req_0 : boolean;
  signal type_cast_2307_inst_ack_0 : boolean;
  signal binary_2313_inst_req_0 : boolean;
  signal binary_2313_inst_ack_0 : boolean;
  signal binary_2313_inst_req_1 : boolean;
  signal binary_2313_inst_ack_1 : boolean;
  signal array_obj_ref_2317_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2317_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2317_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2317_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2317_offset_inst_req_0 : boolean;
  signal array_obj_ref_2317_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2317_base_resize_req_0 : boolean;
  signal array_obj_ref_2317_base_resize_ack_0 : boolean;
  signal array_obj_ref_2317_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2317_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2317_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2317_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2317_final_reg_req_0 : boolean;
  signal array_obj_ref_2317_final_reg_ack_0 : boolean;
  signal ptr_deref_2321_base_resize_req_0 : boolean;
  signal ptr_deref_2321_base_resize_ack_0 : boolean;
  signal ptr_deref_2321_root_address_inst_req_0 : boolean;
  signal ptr_deref_2321_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2321_addr_0_req_0 : boolean;
  signal ptr_deref_2321_addr_0_ack_0 : boolean;
  signal ptr_deref_2321_load_0_req_0 : boolean;
  signal ptr_deref_2321_load_0_ack_0 : boolean;
  signal ptr_deref_2321_load_0_req_1 : boolean;
  signal ptr_deref_2321_load_0_ack_1 : boolean;
  signal ptr_deref_2321_gather_scatter_req_0 : boolean;
  signal ptr_deref_2321_gather_scatter_ack_0 : boolean;
  signal type_cast_2325_inst_req_0 : boolean;
  signal type_cast_2325_inst_ack_0 : boolean;
  signal binary_2331_inst_req_0 : boolean;
  signal binary_2331_inst_ack_0 : boolean;
  signal binary_2331_inst_req_1 : boolean;
  signal binary_2331_inst_ack_1 : boolean;
  signal binary_2336_inst_req_0 : boolean;
  signal binary_2336_inst_ack_0 : boolean;
  signal binary_2336_inst_req_1 : boolean;
  signal binary_2336_inst_ack_1 : boolean;
  signal binary_2341_inst_req_0 : boolean;
  signal binary_2341_inst_ack_0 : boolean;
  signal binary_2341_inst_req_1 : boolean;
  signal binary_2341_inst_ack_1 : boolean;
  signal binary_2346_inst_req_0 : boolean;
  signal binary_2346_inst_ack_0 : boolean;
  signal binary_2346_inst_req_1 : boolean;
  signal binary_2346_inst_ack_1 : boolean;
  signal binary_2351_inst_req_0 : boolean;
  signal binary_2351_inst_ack_0 : boolean;
  signal binary_2351_inst_req_1 : boolean;
  signal binary_2351_inst_ack_1 : boolean;
  signal binary_2356_inst_req_0 : boolean;
  signal binary_2356_inst_ack_0 : boolean;
  signal binary_2356_inst_req_1 : boolean;
  signal binary_2356_inst_ack_1 : boolean;
  signal binary_2361_inst_req_0 : boolean;
  signal binary_2361_inst_ack_0 : boolean;
  signal binary_2361_inst_req_1 : boolean;
  signal binary_2361_inst_ack_1 : boolean;
  signal binary_2366_inst_req_0 : boolean;
  signal binary_2366_inst_ack_0 : boolean;
  signal binary_2366_inst_req_1 : boolean;
  signal binary_2366_inst_ack_1 : boolean;
  signal if_stmt_2374_branch_req_0 : boolean;
  signal if_stmt_2374_branch_ack_1 : boolean;
  signal if_stmt_2374_branch_ack_0 : boolean;
  signal simple_obj_ref_2381_inst_req_0 : boolean;
  signal simple_obj_ref_2381_inst_ack_0 : boolean;
  signal simple_obj_ref_2391_inst_req_0 : boolean;
  signal simple_obj_ref_2391_inst_ack_0 : boolean;
  signal binary_2398_inst_req_0 : boolean;
  signal binary_2398_inst_ack_0 : boolean;
  signal binary_2398_inst_req_1 : boolean;
  signal binary_2398_inst_ack_1 : boolean;
  signal simple_obj_ref_2402_inst_req_0 : boolean;
  signal simple_obj_ref_2402_inst_ack_0 : boolean;
  signal simple_obj_ref_2411_inst_req_0 : boolean;
  signal simple_obj_ref_2411_inst_ack_0 : boolean;
  signal simple_obj_ref_2420_inst_req_0 : boolean;
  signal simple_obj_ref_2420_inst_ack_0 : boolean;
  signal simple_obj_ref_2430_inst_req_0 : boolean;
  signal simple_obj_ref_2430_inst_ack_0 : boolean;
  signal phi_stmt_2129_req_1 : boolean;
  signal type_cast_2133_inst_req_0 : boolean;
  signal type_cast_2133_inst_ack_0 : boolean;
  signal phi_stmt_2129_req_0 : boolean;
  signal phi_stmt_2129_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 1 + 1) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_output_CP_8674: Block -- control-path 
    signal cp_elements: BooleanArray(528 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1);
    finAckJoin: join2 port map(pred0 => fin_req_symbol, pred1 => cp_elements(1), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= false; 
    cp_elements(2) <= cp_elements(499);
    cp_elements(3) <= OrReduce(cp_elements(506) & cp_elements(528));
    simple_obj_ref_2381_inst_req_0 <= cp_elements(3);
    cp_elements(4) <= simple_obj_ref_1902_inst_ack_0;
    cp_elements(5) <= cp_elements(4);
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(7) & cp_elements(8));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1906_inst_req_0 <= cp_elements(6);
    cp_elements(7) <= cp_elements(5);
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= type_cast_1906_inst_ack_0;
    simple_obj_ref_1915_inst_req_0 <= cp_elements(9);
    cp_elements(10) <= simple_obj_ref_1915_inst_ack_0;
    simple_obj_ref_1924_inst_req_0 <= cp_elements(10);
    cp_elements(11) <= simple_obj_ref_1924_inst_ack_0;
    cp_elements(12) <= cp_elements(11);
    cp_elements(13) <= cp_elements(12);
    cpelement_group_14 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(13) & cp_elements(18));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(14),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1929_final_reg_req_0 <= cp_elements(14);
    cp_elements(15) <= cp_elements(12);
    array_obj_ref_1929_base_resize_req_0 <= cp_elements(15);
    cp_elements(16) <= array_obj_ref_1929_base_resize_ack_0;
    array_obj_ref_1929_root_address_inst_req_0 <= cp_elements(16);
    cp_elements(17) <= array_obj_ref_1929_root_address_inst_ack_0;
    array_obj_ref_1929_root_address_inst_req_1 <= cp_elements(17);
    cp_elements(18) <= array_obj_ref_1929_root_address_inst_ack_1;
    cp_elements(19) <= array_obj_ref_1929_final_reg_ack_0;
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(24));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1933_load_0_req_0 <= cp_elements(20);
    cp_elements(21) <= cp_elements(19);
    ptr_deref_1933_base_resize_req_0 <= cp_elements(21);
    cp_elements(22) <= ptr_deref_1933_base_resize_ack_0;
    ptr_deref_1933_root_address_inst_req_0 <= cp_elements(22);
    cp_elements(23) <= ptr_deref_1933_root_address_inst_ack_0;
    ptr_deref_1933_addr_0_req_0 <= cp_elements(23);
    cp_elements(24) <= ptr_deref_1933_addr_0_ack_0;
    cp_elements(25) <= ptr_deref_1933_load_0_ack_0;
    ptr_deref_1933_load_0_req_1 <= cp_elements(25);
    cp_elements(26) <= ptr_deref_1933_load_0_ack_1;
    ptr_deref_1933_gather_scatter_req_0 <= cp_elements(26);
    cp_elements(27) <= ptr_deref_1933_gather_scatter_ack_0;
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1937_inst_req_0 <= cp_elements(28);
    cp_elements(29) <= cp_elements(12);
    cp_elements(30) <= type_cast_1937_inst_ack_0;
    cp_elements(31) <= cp_elements(12);
    cpelement_group_32 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(31) & cp_elements(36));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(32),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1942_final_reg_req_0 <= cp_elements(32);
    cp_elements(33) <= cp_elements(12);
    array_obj_ref_1942_base_resize_req_0 <= cp_elements(33);
    cp_elements(34) <= array_obj_ref_1942_base_resize_ack_0;
    array_obj_ref_1942_root_address_inst_req_0 <= cp_elements(34);
    cp_elements(35) <= array_obj_ref_1942_root_address_inst_ack_0;
    array_obj_ref_1942_root_address_inst_req_1 <= cp_elements(35);
    cp_elements(36) <= array_obj_ref_1942_root_address_inst_ack_1;
    cp_elements(37) <= array_obj_ref_1942_final_reg_ack_0;
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(37) & cp_elements(42));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1946_load_0_req_0 <= cp_elements(38);
    cp_elements(39) <= cp_elements(37);
    ptr_deref_1946_base_resize_req_0 <= cp_elements(39);
    cp_elements(40) <= ptr_deref_1946_base_resize_ack_0;
    ptr_deref_1946_root_address_inst_req_0 <= cp_elements(40);
    cp_elements(41) <= ptr_deref_1946_root_address_inst_ack_0;
    ptr_deref_1946_addr_0_req_0 <= cp_elements(41);
    cp_elements(42) <= ptr_deref_1946_addr_0_ack_0;
    cp_elements(43) <= ptr_deref_1946_load_0_ack_0;
    ptr_deref_1946_load_0_req_1 <= cp_elements(43);
    cp_elements(44) <= ptr_deref_1946_load_0_ack_1;
    ptr_deref_1946_gather_scatter_req_0 <= cp_elements(44);
    cp_elements(45) <= ptr_deref_1946_gather_scatter_ack_0;
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(47));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1950_inst_req_0 <= cp_elements(46);
    cp_elements(47) <= cp_elements(12);
    cp_elements(48) <= type_cast_1950_inst_ack_0;
    cpelement_group_49 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(49),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1956_inst_req_0 <= cp_elements(49);
    cp_elements(50) <= cp_elements(12);
    cp_elements(51) <= binary_1956_inst_ack_0;
    binary_1956_inst_req_1 <= cp_elements(51);
    cp_elements(52) <= binary_1956_inst_ack_1;
    cp_elements(53) <= cp_elements(12);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(58));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1961_final_reg_req_0 <= cp_elements(54);
    cp_elements(55) <= cp_elements(12);
    array_obj_ref_1961_base_resize_req_0 <= cp_elements(55);
    cp_elements(56) <= array_obj_ref_1961_base_resize_ack_0;
    array_obj_ref_1961_root_address_inst_req_0 <= cp_elements(56);
    cp_elements(57) <= array_obj_ref_1961_root_address_inst_ack_0;
    array_obj_ref_1961_root_address_inst_req_1 <= cp_elements(57);
    cp_elements(58) <= array_obj_ref_1961_root_address_inst_ack_1;
    cp_elements(59) <= array_obj_ref_1961_final_reg_ack_0;
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(59) & cp_elements(64));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1965_load_0_req_0 <= cp_elements(60);
    cp_elements(61) <= cp_elements(59);
    ptr_deref_1965_base_resize_req_0 <= cp_elements(61);
    cp_elements(62) <= ptr_deref_1965_base_resize_ack_0;
    ptr_deref_1965_root_address_inst_req_0 <= cp_elements(62);
    cp_elements(63) <= ptr_deref_1965_root_address_inst_ack_0;
    ptr_deref_1965_addr_0_req_0 <= cp_elements(63);
    cp_elements(64) <= ptr_deref_1965_addr_0_ack_0;
    cp_elements(65) <= ptr_deref_1965_load_0_ack_0;
    ptr_deref_1965_load_0_req_1 <= cp_elements(65);
    cp_elements(66) <= ptr_deref_1965_load_0_ack_1;
    ptr_deref_1965_gather_scatter_req_0 <= cp_elements(66);
    cp_elements(67) <= ptr_deref_1965_gather_scatter_ack_0;
    cpelement_group_68 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(67) & cp_elements(69));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(68),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1969_inst_req_0 <= cp_elements(68);
    cp_elements(69) <= cp_elements(12);
    cp_elements(70) <= type_cast_1969_inst_ack_0;
    cpelement_group_71 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(70) & cp_elements(72));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(71),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1975_inst_req_0 <= cp_elements(71);
    cp_elements(72) <= cp_elements(12);
    cp_elements(73) <= binary_1975_inst_ack_0;
    binary_1975_inst_req_1 <= cp_elements(73);
    cp_elements(74) <= binary_1975_inst_ack_1;
    cp_elements(75) <= cp_elements(12);
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(80));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1980_final_reg_req_0 <= cp_elements(76);
    cp_elements(77) <= cp_elements(12);
    array_obj_ref_1980_base_resize_req_0 <= cp_elements(77);
    cp_elements(78) <= array_obj_ref_1980_base_resize_ack_0;
    array_obj_ref_1980_root_address_inst_req_0 <= cp_elements(78);
    cp_elements(79) <= array_obj_ref_1980_root_address_inst_ack_0;
    array_obj_ref_1980_root_address_inst_req_1 <= cp_elements(79);
    cp_elements(80) <= array_obj_ref_1980_root_address_inst_ack_1;
    cp_elements(81) <= array_obj_ref_1980_final_reg_ack_0;
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(86));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_1984_load_0_req_0 <= cp_elements(82);
    cp_elements(83) <= cp_elements(81);
    ptr_deref_1984_base_resize_req_0 <= cp_elements(83);
    cp_elements(84) <= ptr_deref_1984_base_resize_ack_0;
    ptr_deref_1984_root_address_inst_req_0 <= cp_elements(84);
    cp_elements(85) <= ptr_deref_1984_root_address_inst_ack_0;
    ptr_deref_1984_addr_0_req_0 <= cp_elements(85);
    cp_elements(86) <= ptr_deref_1984_addr_0_ack_0;
    cp_elements(87) <= ptr_deref_1984_load_0_ack_0;
    ptr_deref_1984_load_0_req_1 <= cp_elements(87);
    cp_elements(88) <= ptr_deref_1984_load_0_ack_1;
    ptr_deref_1984_gather_scatter_req_0 <= cp_elements(88);
    cp_elements(89) <= ptr_deref_1984_gather_scatter_ack_0;
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(91));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_1988_inst_req_0 <= cp_elements(90);
    cp_elements(91) <= cp_elements(12);
    cp_elements(92) <= type_cast_1988_inst_ack_0;
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(92) & cp_elements(94));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_1994_inst_req_0 <= cp_elements(93);
    cp_elements(94) <= cp_elements(12);
    cp_elements(95) <= binary_1994_inst_ack_0;
    binary_1994_inst_req_1 <= cp_elements(95);
    cp_elements(96) <= binary_1994_inst_ack_1;
    cp_elements(97) <= cp_elements(12);
    cpelement_group_98 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(97) & cp_elements(102));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(98),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_1999_final_reg_req_0 <= cp_elements(98);
    cp_elements(99) <= cp_elements(12);
    array_obj_ref_1999_base_resize_req_0 <= cp_elements(99);
    cp_elements(100) <= array_obj_ref_1999_base_resize_ack_0;
    array_obj_ref_1999_root_address_inst_req_0 <= cp_elements(100);
    cp_elements(101) <= array_obj_ref_1999_root_address_inst_ack_0;
    array_obj_ref_1999_root_address_inst_req_1 <= cp_elements(101);
    cp_elements(102) <= array_obj_ref_1999_root_address_inst_ack_1;
    cp_elements(103) <= array_obj_ref_1999_final_reg_ack_0;
    cpelement_group_104 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(103) & cp_elements(108));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(104),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2003_load_0_req_0 <= cp_elements(104);
    cp_elements(105) <= cp_elements(103);
    ptr_deref_2003_base_resize_req_0 <= cp_elements(105);
    cp_elements(106) <= ptr_deref_2003_base_resize_ack_0;
    ptr_deref_2003_root_address_inst_req_0 <= cp_elements(106);
    cp_elements(107) <= ptr_deref_2003_root_address_inst_ack_0;
    ptr_deref_2003_addr_0_req_0 <= cp_elements(107);
    cp_elements(108) <= ptr_deref_2003_addr_0_ack_0;
    cp_elements(109) <= ptr_deref_2003_load_0_ack_0;
    ptr_deref_2003_load_0_req_1 <= cp_elements(109);
    cp_elements(110) <= ptr_deref_2003_load_0_ack_1;
    ptr_deref_2003_gather_scatter_req_0 <= cp_elements(110);
    cp_elements(111) <= ptr_deref_2003_gather_scatter_ack_0;
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(111) & cp_elements(113));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2007_inst_req_0 <= cp_elements(112);
    cp_elements(113) <= cp_elements(12);
    cp_elements(114) <= type_cast_2007_inst_ack_0;
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(116));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2013_inst_req_0 <= cp_elements(115);
    cp_elements(116) <= cp_elements(12);
    cp_elements(117) <= binary_2013_inst_ack_0;
    binary_2013_inst_req_1 <= cp_elements(117);
    cp_elements(118) <= binary_2013_inst_ack_1;
    cp_elements(119) <= cp_elements(12);
    cpelement_group_120 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(119) & cp_elements(124));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(120),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2018_final_reg_req_0 <= cp_elements(120);
    cp_elements(121) <= cp_elements(12);
    array_obj_ref_2018_base_resize_req_0 <= cp_elements(121);
    cp_elements(122) <= array_obj_ref_2018_base_resize_ack_0;
    array_obj_ref_2018_root_address_inst_req_0 <= cp_elements(122);
    cp_elements(123) <= array_obj_ref_2018_root_address_inst_ack_0;
    array_obj_ref_2018_root_address_inst_req_1 <= cp_elements(123);
    cp_elements(124) <= array_obj_ref_2018_root_address_inst_ack_1;
    cp_elements(125) <= array_obj_ref_2018_final_reg_ack_0;
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(130));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2022_load_0_req_0 <= cp_elements(126);
    cp_elements(127) <= cp_elements(125);
    ptr_deref_2022_base_resize_req_0 <= cp_elements(127);
    cp_elements(128) <= ptr_deref_2022_base_resize_ack_0;
    ptr_deref_2022_root_address_inst_req_0 <= cp_elements(128);
    cp_elements(129) <= ptr_deref_2022_root_address_inst_ack_0;
    ptr_deref_2022_addr_0_req_0 <= cp_elements(129);
    cp_elements(130) <= ptr_deref_2022_addr_0_ack_0;
    cp_elements(131) <= ptr_deref_2022_load_0_ack_0;
    ptr_deref_2022_load_0_req_1 <= cp_elements(131);
    cp_elements(132) <= ptr_deref_2022_load_0_ack_1;
    ptr_deref_2022_gather_scatter_req_0 <= cp_elements(132);
    cp_elements(133) <= ptr_deref_2022_gather_scatter_ack_0;
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(135));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2026_inst_req_0 <= cp_elements(134);
    cp_elements(135) <= cp_elements(12);
    cp_elements(136) <= type_cast_2026_inst_ack_0;
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(136) & cp_elements(138));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2032_inst_req_0 <= cp_elements(137);
    cp_elements(138) <= cp_elements(12);
    cp_elements(139) <= binary_2032_inst_ack_0;
    binary_2032_inst_req_1 <= cp_elements(139);
    cp_elements(140) <= binary_2032_inst_ack_1;
    cpelement_group_141 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(142) & cp_elements(146));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(141),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2036_load_0_req_0 <= cp_elements(141);
    cp_elements(142) <= cp_elements(12);
    cp_elements(143) <= cp_elements(142);
    ptr_deref_2036_base_resize_req_0 <= cp_elements(143);
    cp_elements(144) <= ptr_deref_2036_base_resize_ack_0;
    ptr_deref_2036_root_address_inst_req_0 <= cp_elements(144);
    cp_elements(145) <= ptr_deref_2036_root_address_inst_ack_0;
    ptr_deref_2036_addr_0_req_0 <= cp_elements(145);
    cp_elements(146) <= ptr_deref_2036_addr_0_ack_0;
    cp_elements(147) <= ptr_deref_2036_load_0_ack_0;
    ptr_deref_2036_load_0_req_1 <= cp_elements(147);
    cp_elements(148) <= ptr_deref_2036_load_0_ack_1;
    ptr_deref_2036_gather_scatter_req_0 <= cp_elements(148);
    cp_elements(149) <= ptr_deref_2036_gather_scatter_ack_0;
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(151));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2040_inst_req_0 <= cp_elements(150);
    cp_elements(151) <= cp_elements(12);
    cp_elements(152) <= type_cast_2040_inst_ack_0;
    cpelement_group_153 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(153),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2046_inst_req_0 <= cp_elements(153);
    cp_elements(154) <= cp_elements(12);
    cp_elements(155) <= binary_2046_inst_ack_0;
    binary_2046_inst_req_1 <= cp_elements(155);
    cp_elements(156) <= binary_2046_inst_ack_1;
    cp_elements(157) <= cp_elements(12);
    cpelement_group_158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(157) & cp_elements(162));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2051_final_reg_req_0 <= cp_elements(158);
    cp_elements(159) <= cp_elements(12);
    array_obj_ref_2051_base_resize_req_0 <= cp_elements(159);
    cp_elements(160) <= array_obj_ref_2051_base_resize_ack_0;
    array_obj_ref_2051_root_address_inst_req_0 <= cp_elements(160);
    cp_elements(161) <= array_obj_ref_2051_root_address_inst_ack_0;
    array_obj_ref_2051_root_address_inst_req_1 <= cp_elements(161);
    cp_elements(162) <= array_obj_ref_2051_root_address_inst_ack_1;
    cp_elements(163) <= array_obj_ref_2051_final_reg_ack_0;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(163) & cp_elements(168));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2055_load_0_req_0 <= cp_elements(164);
    cp_elements(165) <= cp_elements(163);
    ptr_deref_2055_base_resize_req_0 <= cp_elements(165);
    cp_elements(166) <= ptr_deref_2055_base_resize_ack_0;
    ptr_deref_2055_root_address_inst_req_0 <= cp_elements(166);
    cp_elements(167) <= ptr_deref_2055_root_address_inst_ack_0;
    ptr_deref_2055_addr_0_req_0 <= cp_elements(167);
    cp_elements(168) <= ptr_deref_2055_addr_0_ack_0;
    cp_elements(169) <= ptr_deref_2055_load_0_ack_0;
    ptr_deref_2055_load_0_req_1 <= cp_elements(169);
    cp_elements(170) <= ptr_deref_2055_load_0_ack_1;
    ptr_deref_2055_gather_scatter_req_0 <= cp_elements(170);
    cp_elements(171) <= ptr_deref_2055_gather_scatter_ack_0;
    cpelement_group_172 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(171) & cp_elements(173));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(172),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2059_inst_req_0 <= cp_elements(172);
    cp_elements(173) <= cp_elements(12);
    cp_elements(174) <= type_cast_2059_inst_ack_0;
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(174) & cp_elements(176));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2065_inst_req_0 <= cp_elements(175);
    cp_elements(176) <= cp_elements(12);
    cp_elements(177) <= binary_2065_inst_ack_0;
    binary_2065_inst_req_1 <= cp_elements(177);
    cp_elements(178) <= binary_2065_inst_ack_1;
    cpelement_group_179 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(52) & cp_elements(180));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(179),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2070_inst_req_0 <= cp_elements(179);
    cp_elements(180) <= cp_elements(12);
    cp_elements(181) <= binary_2070_inst_ack_0;
    binary_2070_inst_req_1 <= cp_elements(181);
    cp_elements(182) <= binary_2070_inst_ack_1;
    cpelement_group_183 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(182) & cp_elements(184));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(183),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2075_inst_req_0 <= cp_elements(183);
    cp_elements(184) <= cp_elements(12);
    cp_elements(185) <= binary_2075_inst_ack_0;
    binary_2075_inst_req_1 <= cp_elements(185);
    cp_elements(186) <= binary_2075_inst_ack_1;
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(96) & cp_elements(186) & cp_elements(188));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2080_inst_req_0 <= cp_elements(187);
    cp_elements(188) <= cp_elements(12);
    cp_elements(189) <= binary_2080_inst_ack_0;
    binary_2080_inst_req_1 <= cp_elements(189);
    cp_elements(190) <= binary_2080_inst_ack_1;
    cpelement_group_191 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(190) & cp_elements(192));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(191),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2085_inst_req_0 <= cp_elements(191);
    cp_elements(192) <= cp_elements(12);
    cp_elements(193) <= binary_2085_inst_ack_0;
    binary_2085_inst_req_1 <= cp_elements(193);
    cp_elements(194) <= binary_2085_inst_ack_1;
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(140) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2090_inst_req_0 <= cp_elements(195);
    cp_elements(196) <= cp_elements(12);
    cp_elements(197) <= binary_2090_inst_ack_0;
    binary_2090_inst_req_1 <= cp_elements(197);
    cp_elements(198) <= binary_2090_inst_ack_1;
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(198) & cp_elements(200));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2095_inst_req_0 <= cp_elements(199);
    cp_elements(200) <= cp_elements(12);
    cp_elements(201) <= binary_2095_inst_ack_0;
    binary_2095_inst_req_1 <= cp_elements(201);
    cp_elements(202) <= binary_2095_inst_ack_1;
    cpelement_group_203 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(202) & cp_elements(204));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(203),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2100_inst_req_0 <= cp_elements(203);
    cp_elements(204) <= cp_elements(12);
    cp_elements(205) <= binary_2100_inst_ack_0;
    binary_2100_inst_req_1 <= cp_elements(205);
    cp_elements(206) <= binary_2100_inst_ack_1;
    simple_obj_ref_2108_inst_req_0 <= cp_elements(206);
    cp_elements(207) <= simple_obj_ref_2108_inst_ack_0;
    simple_obj_ref_2118_inst_req_0 <= cp_elements(207);
    cp_elements(208) <= simple_obj_ref_2118_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    cpelement_group_210 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(212));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(210),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2125_inst_req_0 <= cp_elements(210);
    cp_elements(211) <= cp_elements(209);
    cp_elements(212) <= cp_elements(209);
    cp_elements(213) <= binary_2125_inst_ack_0;
    binary_2125_inst_req_1 <= cp_elements(213);
    cp_elements(214) <= binary_2125_inst_ack_1;
    phi_stmt_2129_req_1 <= cp_elements(214);
    cp_elements(215) <= cp_elements(526);
    cpelement_group_216 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(217) & cp_elements(218));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(216),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2140_inst_req_0 <= cp_elements(216);
    cp_elements(217) <= cp_elements(215);
    cp_elements(218) <= cp_elements(215);
    cp_elements(219) <= type_cast_2140_inst_ack_0;
    cpelement_group_220 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(221) & cp_elements(222) & cp_elements(223));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(220),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2145_inst_req_0 <= cp_elements(220);
    cp_elements(221) <= cp_elements(215);
    cp_elements(222) <= cp_elements(219);
    cp_elements(223) <= cp_elements(215);
    cp_elements(224) <= binary_2145_inst_ack_0;
    binary_2145_inst_req_1 <= cp_elements(224);
    cp_elements(225) <= binary_2145_inst_ack_1;
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(227) & cp_elements(228));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2151_inst_req_0 <= cp_elements(226);
    cp_elements(227) <= cp_elements(215);
    cp_elements(228) <= cp_elements(219);
    cp_elements(229) <= binary_2151_inst_ack_0;
    binary_2151_inst_req_1 <= cp_elements(229);
    cp_elements(230) <= binary_2151_inst_ack_1;
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(232) & cp_elements(233));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2157_inst_req_0 <= cp_elements(231);
    cp_elements(232) <= cp_elements(215);
    cp_elements(233) <= cp_elements(230);
    cp_elements(234) <= binary_2157_inst_ack_0;
    binary_2157_inst_req_1 <= cp_elements(234);
    cp_elements(235) <= binary_2157_inst_ack_1;
    array_obj_ref_2161_index_0_resize_req_0 <= cp_elements(235);
    cp_elements(236) <= cp_elements(215);
    cpelement_group_237 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(236) & cp_elements(245));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(237),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2161_final_reg_req_0 <= cp_elements(237);
    cp_elements(238) <= cp_elements(215);
    array_obj_ref_2161_base_resize_req_0 <= cp_elements(238);
    cp_elements(239) <= array_obj_ref_2161_index_0_resize_ack_0;
    array_obj_ref_2161_index_0_rename_req_0 <= cp_elements(239);
    cp_elements(240) <= array_obj_ref_2161_index_0_rename_ack_0;
    array_obj_ref_2161_offset_inst_req_0 <= cp_elements(240);
    cp_elements(241) <= array_obj_ref_2161_offset_inst_ack_0;
    cp_elements(242) <= array_obj_ref_2161_base_resize_ack_0;
    cpelement_group_243 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(241) & cp_elements(242));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(243),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2161_root_address_inst_req_0 <= cp_elements(243);
    cp_elements(244) <= array_obj_ref_2161_root_address_inst_ack_0;
    array_obj_ref_2161_root_address_inst_req_1 <= cp_elements(244);
    cp_elements(245) <= array_obj_ref_2161_root_address_inst_ack_1;
    cp_elements(246) <= array_obj_ref_2161_final_reg_ack_0;
    cpelement_group_247 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(246) & cp_elements(251));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(247),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2165_load_0_req_0 <= cp_elements(247);
    cp_elements(248) <= cp_elements(246);
    ptr_deref_2165_base_resize_req_0 <= cp_elements(248);
    cp_elements(249) <= ptr_deref_2165_base_resize_ack_0;
    ptr_deref_2165_root_address_inst_req_0 <= cp_elements(249);
    cp_elements(250) <= ptr_deref_2165_root_address_inst_ack_0;
    ptr_deref_2165_addr_0_req_0 <= cp_elements(250);
    cp_elements(251) <= ptr_deref_2165_addr_0_ack_0;
    cp_elements(252) <= ptr_deref_2165_load_0_ack_0;
    ptr_deref_2165_load_0_req_1 <= cp_elements(252);
    cp_elements(253) <= ptr_deref_2165_load_0_ack_1;
    ptr_deref_2165_gather_scatter_req_0 <= cp_elements(253);
    cp_elements(254) <= ptr_deref_2165_gather_scatter_ack_0;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(256));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2169_inst_req_0 <= cp_elements(255);
    cp_elements(256) <= cp_elements(215);
    cp_elements(257) <= type_cast_2169_inst_ack_0;
    cpelement_group_258 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(259) & cp_elements(260));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(258),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2175_inst_req_0 <= cp_elements(258);
    cp_elements(259) <= cp_elements(215);
    cp_elements(260) <= cp_elements(230);
    cp_elements(261) <= binary_2175_inst_ack_0;
    binary_2175_inst_req_1 <= cp_elements(261);
    cp_elements(262) <= binary_2175_inst_ack_1;
    array_obj_ref_2179_index_0_resize_req_0 <= cp_elements(262);
    cp_elements(263) <= cp_elements(215);
    cpelement_group_264 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(263) & cp_elements(272));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(264),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2179_final_reg_req_0 <= cp_elements(264);
    cp_elements(265) <= cp_elements(215);
    array_obj_ref_2179_base_resize_req_0 <= cp_elements(265);
    cp_elements(266) <= array_obj_ref_2179_index_0_resize_ack_0;
    array_obj_ref_2179_index_0_rename_req_0 <= cp_elements(266);
    cp_elements(267) <= array_obj_ref_2179_index_0_rename_ack_0;
    array_obj_ref_2179_offset_inst_req_0 <= cp_elements(267);
    cp_elements(268) <= array_obj_ref_2179_offset_inst_ack_0;
    cp_elements(269) <= array_obj_ref_2179_base_resize_ack_0;
    cpelement_group_270 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(268) & cp_elements(269));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(270),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2179_root_address_inst_req_0 <= cp_elements(270);
    cp_elements(271) <= array_obj_ref_2179_root_address_inst_ack_0;
    array_obj_ref_2179_root_address_inst_req_1 <= cp_elements(271);
    cp_elements(272) <= array_obj_ref_2179_root_address_inst_ack_1;
    cp_elements(273) <= array_obj_ref_2179_final_reg_ack_0;
    cpelement_group_274 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(273) & cp_elements(278));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(274),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2183_load_0_req_0 <= cp_elements(274);
    cp_elements(275) <= cp_elements(273);
    ptr_deref_2183_base_resize_req_0 <= cp_elements(275);
    cp_elements(276) <= ptr_deref_2183_base_resize_ack_0;
    ptr_deref_2183_root_address_inst_req_0 <= cp_elements(276);
    cp_elements(277) <= ptr_deref_2183_root_address_inst_ack_0;
    ptr_deref_2183_addr_0_req_0 <= cp_elements(277);
    cp_elements(278) <= ptr_deref_2183_addr_0_ack_0;
    cp_elements(279) <= ptr_deref_2183_load_0_ack_0;
    ptr_deref_2183_load_0_req_1 <= cp_elements(279);
    cp_elements(280) <= ptr_deref_2183_load_0_ack_1;
    ptr_deref_2183_gather_scatter_req_0 <= cp_elements(280);
    cp_elements(281) <= ptr_deref_2183_gather_scatter_ack_0;
    cpelement_group_282 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(281) & cp_elements(283));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(282),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2187_inst_req_0 <= cp_elements(282);
    cp_elements(283) <= cp_elements(215);
    cp_elements(284) <= type_cast_2187_inst_ack_0;
    cpelement_group_285 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(284) & cp_elements(286));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(285),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2193_inst_req_0 <= cp_elements(285);
    cp_elements(286) <= cp_elements(215);
    cp_elements(287) <= binary_2193_inst_ack_0;
    binary_2193_inst_req_1 <= cp_elements(287);
    cp_elements(288) <= binary_2193_inst_ack_1;
    cpelement_group_289 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(290) & cp_elements(291));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(289),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2199_inst_req_0 <= cp_elements(289);
    cp_elements(290) <= cp_elements(215);
    cp_elements(291) <= cp_elements(230);
    cp_elements(292) <= binary_2199_inst_ack_0;
    binary_2199_inst_req_1 <= cp_elements(292);
    cp_elements(293) <= binary_2199_inst_ack_1;
    array_obj_ref_2203_index_0_resize_req_0 <= cp_elements(293);
    cp_elements(294) <= cp_elements(215);
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(294) & cp_elements(303));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2203_final_reg_req_0 <= cp_elements(295);
    cp_elements(296) <= cp_elements(215);
    array_obj_ref_2203_base_resize_req_0 <= cp_elements(296);
    cp_elements(297) <= array_obj_ref_2203_index_0_resize_ack_0;
    array_obj_ref_2203_index_0_rename_req_0 <= cp_elements(297);
    cp_elements(298) <= array_obj_ref_2203_index_0_rename_ack_0;
    array_obj_ref_2203_offset_inst_req_0 <= cp_elements(298);
    cp_elements(299) <= array_obj_ref_2203_offset_inst_ack_0;
    cp_elements(300) <= array_obj_ref_2203_base_resize_ack_0;
    cpelement_group_301 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(301),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2203_root_address_inst_req_0 <= cp_elements(301);
    cp_elements(302) <= array_obj_ref_2203_root_address_inst_ack_0;
    array_obj_ref_2203_root_address_inst_req_1 <= cp_elements(302);
    cp_elements(303) <= array_obj_ref_2203_root_address_inst_ack_1;
    cp_elements(304) <= array_obj_ref_2203_final_reg_ack_0;
    cpelement_group_305 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(304) & cp_elements(309));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(305),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2207_load_0_req_0 <= cp_elements(305);
    cp_elements(306) <= cp_elements(304);
    ptr_deref_2207_base_resize_req_0 <= cp_elements(306);
    cp_elements(307) <= ptr_deref_2207_base_resize_ack_0;
    ptr_deref_2207_root_address_inst_req_0 <= cp_elements(307);
    cp_elements(308) <= ptr_deref_2207_root_address_inst_ack_0;
    ptr_deref_2207_addr_0_req_0 <= cp_elements(308);
    cp_elements(309) <= ptr_deref_2207_addr_0_ack_0;
    cp_elements(310) <= ptr_deref_2207_load_0_ack_0;
    ptr_deref_2207_load_0_req_1 <= cp_elements(310);
    cp_elements(311) <= ptr_deref_2207_load_0_ack_1;
    ptr_deref_2207_gather_scatter_req_0 <= cp_elements(311);
    cp_elements(312) <= ptr_deref_2207_gather_scatter_ack_0;
    cpelement_group_313 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(312) & cp_elements(314));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(313),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2211_inst_req_0 <= cp_elements(313);
    cp_elements(314) <= cp_elements(215);
    cp_elements(315) <= type_cast_2211_inst_ack_0;
    cpelement_group_316 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(315) & cp_elements(317));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(316),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2217_inst_req_0 <= cp_elements(316);
    cp_elements(317) <= cp_elements(215);
    cp_elements(318) <= binary_2217_inst_ack_0;
    binary_2217_inst_req_1 <= cp_elements(318);
    cp_elements(319) <= binary_2217_inst_ack_1;
    cpelement_group_320 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(321) & cp_elements(322));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(320),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2223_inst_req_0 <= cp_elements(320);
    cp_elements(321) <= cp_elements(215);
    cp_elements(322) <= cp_elements(230);
    cp_elements(323) <= binary_2223_inst_ack_0;
    binary_2223_inst_req_1 <= cp_elements(323);
    cp_elements(324) <= binary_2223_inst_ack_1;
    array_obj_ref_2227_index_0_resize_req_0 <= cp_elements(324);
    cp_elements(325) <= cp_elements(215);
    cpelement_group_326 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(325) & cp_elements(334));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(326),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2227_final_reg_req_0 <= cp_elements(326);
    cp_elements(327) <= cp_elements(215);
    array_obj_ref_2227_base_resize_req_0 <= cp_elements(327);
    cp_elements(328) <= array_obj_ref_2227_index_0_resize_ack_0;
    array_obj_ref_2227_index_0_rename_req_0 <= cp_elements(328);
    cp_elements(329) <= array_obj_ref_2227_index_0_rename_ack_0;
    array_obj_ref_2227_offset_inst_req_0 <= cp_elements(329);
    cp_elements(330) <= array_obj_ref_2227_offset_inst_ack_0;
    cp_elements(331) <= array_obj_ref_2227_base_resize_ack_0;
    cpelement_group_332 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(330) & cp_elements(331));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(332),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2227_root_address_inst_req_0 <= cp_elements(332);
    cp_elements(333) <= array_obj_ref_2227_root_address_inst_ack_0;
    array_obj_ref_2227_root_address_inst_req_1 <= cp_elements(333);
    cp_elements(334) <= array_obj_ref_2227_root_address_inst_ack_1;
    cp_elements(335) <= array_obj_ref_2227_final_reg_ack_0;
    cpelement_group_336 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(335) & cp_elements(340));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(336),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2231_load_0_req_0 <= cp_elements(336);
    cp_elements(337) <= cp_elements(335);
    ptr_deref_2231_base_resize_req_0 <= cp_elements(337);
    cp_elements(338) <= ptr_deref_2231_base_resize_ack_0;
    ptr_deref_2231_root_address_inst_req_0 <= cp_elements(338);
    cp_elements(339) <= ptr_deref_2231_root_address_inst_ack_0;
    ptr_deref_2231_addr_0_req_0 <= cp_elements(339);
    cp_elements(340) <= ptr_deref_2231_addr_0_ack_0;
    cp_elements(341) <= ptr_deref_2231_load_0_ack_0;
    ptr_deref_2231_load_0_req_1 <= cp_elements(341);
    cp_elements(342) <= ptr_deref_2231_load_0_ack_1;
    ptr_deref_2231_gather_scatter_req_0 <= cp_elements(342);
    cp_elements(343) <= ptr_deref_2231_gather_scatter_ack_0;
    cpelement_group_344 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(343) & cp_elements(345));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2235_inst_req_0 <= cp_elements(344);
    cp_elements(345) <= cp_elements(215);
    cp_elements(346) <= type_cast_2235_inst_ack_0;
    cpelement_group_347 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(346) & cp_elements(348));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(347),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2241_inst_req_0 <= cp_elements(347);
    cp_elements(348) <= cp_elements(215);
    cp_elements(349) <= binary_2241_inst_ack_0;
    binary_2241_inst_req_1 <= cp_elements(349);
    cp_elements(350) <= binary_2241_inst_ack_1;
    cpelement_group_351 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(352) & cp_elements(353));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(351),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2247_inst_req_0 <= cp_elements(351);
    cp_elements(352) <= cp_elements(215);
    cp_elements(353) <= cp_elements(230);
    cp_elements(354) <= binary_2247_inst_ack_0;
    binary_2247_inst_req_1 <= cp_elements(354);
    cp_elements(355) <= binary_2247_inst_ack_1;
    array_obj_ref_2251_index_0_resize_req_0 <= cp_elements(355);
    cp_elements(356) <= cp_elements(215);
    cpelement_group_357 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(356) & cp_elements(365));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(357),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2251_final_reg_req_0 <= cp_elements(357);
    cp_elements(358) <= cp_elements(215);
    array_obj_ref_2251_base_resize_req_0 <= cp_elements(358);
    cp_elements(359) <= array_obj_ref_2251_index_0_resize_ack_0;
    array_obj_ref_2251_index_0_rename_req_0 <= cp_elements(359);
    cp_elements(360) <= array_obj_ref_2251_index_0_rename_ack_0;
    array_obj_ref_2251_offset_inst_req_0 <= cp_elements(360);
    cp_elements(361) <= array_obj_ref_2251_offset_inst_ack_0;
    cp_elements(362) <= array_obj_ref_2251_base_resize_ack_0;
    cpelement_group_363 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(362));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2251_root_address_inst_req_0 <= cp_elements(363);
    cp_elements(364) <= array_obj_ref_2251_root_address_inst_ack_0;
    array_obj_ref_2251_root_address_inst_req_1 <= cp_elements(364);
    cp_elements(365) <= array_obj_ref_2251_root_address_inst_ack_1;
    cp_elements(366) <= array_obj_ref_2251_final_reg_ack_0;
    cpelement_group_367 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(366) & cp_elements(371));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(367),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2255_load_0_req_0 <= cp_elements(367);
    cp_elements(368) <= cp_elements(366);
    ptr_deref_2255_base_resize_req_0 <= cp_elements(368);
    cp_elements(369) <= ptr_deref_2255_base_resize_ack_0;
    ptr_deref_2255_root_address_inst_req_0 <= cp_elements(369);
    cp_elements(370) <= ptr_deref_2255_root_address_inst_ack_0;
    ptr_deref_2255_addr_0_req_0 <= cp_elements(370);
    cp_elements(371) <= ptr_deref_2255_addr_0_ack_0;
    cp_elements(372) <= ptr_deref_2255_load_0_ack_0;
    ptr_deref_2255_load_0_req_1 <= cp_elements(372);
    cp_elements(373) <= ptr_deref_2255_load_0_ack_1;
    ptr_deref_2255_gather_scatter_req_0 <= cp_elements(373);
    cp_elements(374) <= ptr_deref_2255_gather_scatter_ack_0;
    cpelement_group_375 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(374) & cp_elements(376));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(375),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2259_inst_req_0 <= cp_elements(375);
    cp_elements(376) <= cp_elements(215);
    cp_elements(377) <= type_cast_2259_inst_ack_0;
    cpelement_group_378 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(377) & cp_elements(379));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(378),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2265_inst_req_0 <= cp_elements(378);
    cp_elements(379) <= cp_elements(215);
    cp_elements(380) <= binary_2265_inst_ack_0;
    binary_2265_inst_req_1 <= cp_elements(380);
    cp_elements(381) <= binary_2265_inst_ack_1;
    cpelement_group_382 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(383) & cp_elements(384));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(382),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2271_inst_req_0 <= cp_elements(382);
    cp_elements(383) <= cp_elements(215);
    cp_elements(384) <= cp_elements(230);
    cp_elements(385) <= binary_2271_inst_ack_0;
    binary_2271_inst_req_1 <= cp_elements(385);
    cp_elements(386) <= binary_2271_inst_ack_1;
    array_obj_ref_2275_index_0_resize_req_0 <= cp_elements(386);
    cp_elements(387) <= cp_elements(215);
    cpelement_group_388 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(387) & cp_elements(396));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(388),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2275_final_reg_req_0 <= cp_elements(388);
    cp_elements(389) <= cp_elements(215);
    array_obj_ref_2275_base_resize_req_0 <= cp_elements(389);
    cp_elements(390) <= array_obj_ref_2275_index_0_resize_ack_0;
    array_obj_ref_2275_index_0_rename_req_0 <= cp_elements(390);
    cp_elements(391) <= array_obj_ref_2275_index_0_rename_ack_0;
    array_obj_ref_2275_offset_inst_req_0 <= cp_elements(391);
    cp_elements(392) <= array_obj_ref_2275_offset_inst_ack_0;
    cp_elements(393) <= array_obj_ref_2275_base_resize_ack_0;
    cpelement_group_394 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(392) & cp_elements(393));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(394),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2275_root_address_inst_req_0 <= cp_elements(394);
    cp_elements(395) <= array_obj_ref_2275_root_address_inst_ack_0;
    array_obj_ref_2275_root_address_inst_req_1 <= cp_elements(395);
    cp_elements(396) <= array_obj_ref_2275_root_address_inst_ack_1;
    cp_elements(397) <= array_obj_ref_2275_final_reg_ack_0;
    cpelement_group_398 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(397) & cp_elements(402));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(398),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2279_load_0_req_0 <= cp_elements(398);
    cp_elements(399) <= cp_elements(397);
    ptr_deref_2279_base_resize_req_0 <= cp_elements(399);
    cp_elements(400) <= ptr_deref_2279_base_resize_ack_0;
    ptr_deref_2279_root_address_inst_req_0 <= cp_elements(400);
    cp_elements(401) <= ptr_deref_2279_root_address_inst_ack_0;
    ptr_deref_2279_addr_0_req_0 <= cp_elements(401);
    cp_elements(402) <= ptr_deref_2279_addr_0_ack_0;
    cp_elements(403) <= ptr_deref_2279_load_0_ack_0;
    ptr_deref_2279_load_0_req_1 <= cp_elements(403);
    cp_elements(404) <= ptr_deref_2279_load_0_ack_1;
    ptr_deref_2279_gather_scatter_req_0 <= cp_elements(404);
    cp_elements(405) <= ptr_deref_2279_gather_scatter_ack_0;
    cpelement_group_406 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(405) & cp_elements(407));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(406),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2283_inst_req_0 <= cp_elements(406);
    cp_elements(407) <= cp_elements(215);
    cp_elements(408) <= type_cast_2283_inst_ack_0;
    cpelement_group_409 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(408) & cp_elements(410));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(409),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2289_inst_req_0 <= cp_elements(409);
    cp_elements(410) <= cp_elements(215);
    cp_elements(411) <= binary_2289_inst_ack_0;
    binary_2289_inst_req_1 <= cp_elements(411);
    cp_elements(412) <= binary_2289_inst_ack_1;
    cpelement_group_413 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(414) & cp_elements(415));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(413),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2295_inst_req_0 <= cp_elements(413);
    cp_elements(414) <= cp_elements(215);
    cp_elements(415) <= cp_elements(230);
    cp_elements(416) <= binary_2295_inst_ack_0;
    binary_2295_inst_req_1 <= cp_elements(416);
    cp_elements(417) <= binary_2295_inst_ack_1;
    array_obj_ref_2299_index_0_resize_req_0 <= cp_elements(417);
    cp_elements(418) <= cp_elements(215);
    cpelement_group_419 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(418) & cp_elements(427));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(419),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2299_final_reg_req_0 <= cp_elements(419);
    cp_elements(420) <= cp_elements(215);
    array_obj_ref_2299_base_resize_req_0 <= cp_elements(420);
    cp_elements(421) <= array_obj_ref_2299_index_0_resize_ack_0;
    array_obj_ref_2299_index_0_rename_req_0 <= cp_elements(421);
    cp_elements(422) <= array_obj_ref_2299_index_0_rename_ack_0;
    array_obj_ref_2299_offset_inst_req_0 <= cp_elements(422);
    cp_elements(423) <= array_obj_ref_2299_offset_inst_ack_0;
    cp_elements(424) <= array_obj_ref_2299_base_resize_ack_0;
    cpelement_group_425 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(423) & cp_elements(424));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(425),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2299_root_address_inst_req_0 <= cp_elements(425);
    cp_elements(426) <= array_obj_ref_2299_root_address_inst_ack_0;
    array_obj_ref_2299_root_address_inst_req_1 <= cp_elements(426);
    cp_elements(427) <= array_obj_ref_2299_root_address_inst_ack_1;
    cp_elements(428) <= array_obj_ref_2299_final_reg_ack_0;
    cpelement_group_429 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(428) & cp_elements(433));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(429),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2303_load_0_req_0 <= cp_elements(429);
    cp_elements(430) <= cp_elements(428);
    ptr_deref_2303_base_resize_req_0 <= cp_elements(430);
    cp_elements(431) <= ptr_deref_2303_base_resize_ack_0;
    ptr_deref_2303_root_address_inst_req_0 <= cp_elements(431);
    cp_elements(432) <= ptr_deref_2303_root_address_inst_ack_0;
    ptr_deref_2303_addr_0_req_0 <= cp_elements(432);
    cp_elements(433) <= ptr_deref_2303_addr_0_ack_0;
    cp_elements(434) <= ptr_deref_2303_load_0_ack_0;
    ptr_deref_2303_load_0_req_1 <= cp_elements(434);
    cp_elements(435) <= ptr_deref_2303_load_0_ack_1;
    ptr_deref_2303_gather_scatter_req_0 <= cp_elements(435);
    cp_elements(436) <= ptr_deref_2303_gather_scatter_ack_0;
    cpelement_group_437 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(436) & cp_elements(438));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(437),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2307_inst_req_0 <= cp_elements(437);
    cp_elements(438) <= cp_elements(215);
    cp_elements(439) <= type_cast_2307_inst_ack_0;
    cpelement_group_440 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(439) & cp_elements(441));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(440),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2313_inst_req_0 <= cp_elements(440);
    cp_elements(441) <= cp_elements(215);
    cp_elements(442) <= binary_2313_inst_ack_0;
    binary_2313_inst_req_1 <= cp_elements(442);
    cp_elements(443) <= binary_2313_inst_ack_1;
    cp_elements(444) <= cp_elements(215);
    cpelement_group_445 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(444) & cp_elements(454));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(445),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2317_final_reg_req_0 <= cp_elements(445);
    cp_elements(446) <= cp_elements(215);
    array_obj_ref_2317_base_resize_req_0 <= cp_elements(446);
    cp_elements(447) <= cp_elements(230);
    array_obj_ref_2317_index_0_resize_req_0 <= cp_elements(447);
    cp_elements(448) <= array_obj_ref_2317_index_0_resize_ack_0;
    array_obj_ref_2317_index_0_rename_req_0 <= cp_elements(448);
    cp_elements(449) <= array_obj_ref_2317_index_0_rename_ack_0;
    array_obj_ref_2317_offset_inst_req_0 <= cp_elements(449);
    cp_elements(450) <= array_obj_ref_2317_offset_inst_ack_0;
    cp_elements(451) <= array_obj_ref_2317_base_resize_ack_0;
    cpelement_group_452 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(450) & cp_elements(451));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(452),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    array_obj_ref_2317_root_address_inst_req_0 <= cp_elements(452);
    cp_elements(453) <= array_obj_ref_2317_root_address_inst_ack_0;
    array_obj_ref_2317_root_address_inst_req_1 <= cp_elements(453);
    cp_elements(454) <= array_obj_ref_2317_root_address_inst_ack_1;
    cp_elements(455) <= array_obj_ref_2317_final_reg_ack_0;
    cpelement_group_456 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(455) & cp_elements(460));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(456),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    ptr_deref_2321_load_0_req_0 <= cp_elements(456);
    cp_elements(457) <= cp_elements(455);
    ptr_deref_2321_base_resize_req_0 <= cp_elements(457);
    cp_elements(458) <= ptr_deref_2321_base_resize_ack_0;
    ptr_deref_2321_root_address_inst_req_0 <= cp_elements(458);
    cp_elements(459) <= ptr_deref_2321_root_address_inst_ack_0;
    ptr_deref_2321_addr_0_req_0 <= cp_elements(459);
    cp_elements(460) <= ptr_deref_2321_addr_0_ack_0;
    cp_elements(461) <= ptr_deref_2321_load_0_ack_0;
    ptr_deref_2321_load_0_req_1 <= cp_elements(461);
    cp_elements(462) <= ptr_deref_2321_load_0_ack_1;
    ptr_deref_2321_gather_scatter_req_0 <= cp_elements(462);
    cp_elements(463) <= ptr_deref_2321_gather_scatter_ack_0;
    cpelement_group_464 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(463) & cp_elements(465));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(464),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    type_cast_2325_inst_req_0 <= cp_elements(464);
    cp_elements(465) <= cp_elements(215);
    cp_elements(466) <= type_cast_2325_inst_ack_0;
    cpelement_group_467 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(466) & cp_elements(468));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(467),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2331_inst_req_0 <= cp_elements(467);
    cp_elements(468) <= cp_elements(215);
    cp_elements(469) <= binary_2331_inst_ack_0;
    binary_2331_inst_req_1 <= cp_elements(469);
    cp_elements(470) <= binary_2331_inst_ack_1;
    cpelement_group_471 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(257) & cp_elements(288) & cp_elements(472));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(471),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2336_inst_req_0 <= cp_elements(471);
    cp_elements(472) <= cp_elements(215);
    cp_elements(473) <= binary_2336_inst_ack_0;
    binary_2336_inst_req_1 <= cp_elements(473);
    cp_elements(474) <= binary_2336_inst_ack_1;
    cpelement_group_475 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(474) & cp_elements(476));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(475),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2341_inst_req_0 <= cp_elements(475);
    cp_elements(476) <= cp_elements(215);
    cp_elements(477) <= binary_2341_inst_ack_0;
    binary_2341_inst_req_1 <= cp_elements(477);
    cp_elements(478) <= binary_2341_inst_ack_1;
    cpelement_group_479 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(350) & cp_elements(478) & cp_elements(480));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(479),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2346_inst_req_0 <= cp_elements(479);
    cp_elements(480) <= cp_elements(215);
    cp_elements(481) <= binary_2346_inst_ack_0;
    binary_2346_inst_req_1 <= cp_elements(481);
    cp_elements(482) <= binary_2346_inst_ack_1;
    cpelement_group_483 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(381) & cp_elements(482) & cp_elements(484));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(483),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2351_inst_req_0 <= cp_elements(483);
    cp_elements(484) <= cp_elements(215);
    cp_elements(485) <= binary_2351_inst_ack_0;
    binary_2351_inst_req_1 <= cp_elements(485);
    cp_elements(486) <= binary_2351_inst_ack_1;
    cpelement_group_487 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(412) & cp_elements(486) & cp_elements(488));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(487),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2356_inst_req_0 <= cp_elements(487);
    cp_elements(488) <= cp_elements(215);
    cp_elements(489) <= binary_2356_inst_ack_0;
    binary_2356_inst_req_1 <= cp_elements(489);
    cp_elements(490) <= binary_2356_inst_ack_1;
    cpelement_group_491 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(443) & cp_elements(490) & cp_elements(492));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(491),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2361_inst_req_0 <= cp_elements(491);
    cp_elements(492) <= cp_elements(215);
    cp_elements(493) <= binary_2361_inst_ack_0;
    binary_2361_inst_req_1 <= cp_elements(493);
    cp_elements(494) <= binary_2361_inst_ack_1;
    cpelement_group_495 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(470) & cp_elements(494) & cp_elements(496));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(495),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2366_inst_req_0 <= cp_elements(495);
    cp_elements(496) <= cp_elements(215);
    cp_elements(497) <= binary_2366_inst_ack_0;
    binary_2366_inst_req_1 <= cp_elements(497);
    cp_elements(498) <= binary_2366_inst_ack_1;
    cpelement_group_499 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(225) & cp_elements(498));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(499),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(500) <= cp_elements(2);
    cp_elements(501) <= false;
    cp_elements(502) <= cp_elements(501);
    cp_elements(503) <= cp_elements(2);
    if_stmt_2374_branch_req_0 <= cp_elements(503);
    cp_elements(504) <= cp_elements(503);
    cp_elements(505) <= cp_elements(504);
    cp_elements(506) <= if_stmt_2374_branch_ack_1;
    cp_elements(507) <= cp_elements(504);
    cp_elements(508) <= if_stmt_2374_branch_ack_0;
    simple_obj_ref_2402_inst_req_0 <= cp_elements(508);
    cp_elements(509) <= simple_obj_ref_2381_inst_ack_0;
    simple_obj_ref_2391_inst_req_0 <= cp_elements(509);
    cp_elements(510) <= simple_obj_ref_2391_inst_ack_0;
    cp_elements(511) <= cp_elements(510);
    cpelement_group_512 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(513) & cp_elements(514));
      jNoI: join -- 
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(512),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    binary_2398_inst_req_0 <= cp_elements(512);
    cp_elements(513) <= cp_elements(511);
    cp_elements(514) <= cp_elements(511);
    cp_elements(515) <= binary_2398_inst_ack_0;
    binary_2398_inst_req_1 <= cp_elements(515);
    cp_elements(516) <= binary_2398_inst_ack_1;
    type_cast_2133_inst_req_0 <= cp_elements(516);
    cp_elements(517) <= simple_obj_ref_2402_inst_ack_0;
    simple_obj_ref_2411_inst_req_0 <= cp_elements(517);
    cp_elements(518) <= simple_obj_ref_2411_inst_ack_0;
    simple_obj_ref_2420_inst_req_0 <= cp_elements(518);
    cp_elements(519) <= simple_obj_ref_2420_inst_ack_0;
    simple_obj_ref_2430_inst_req_0 <= cp_elements(519);
    cp_elements(520) <= simple_obj_ref_2430_inst_ack_0;
    cp_elements(521) <= OrReduce(cp_elements(0) & cp_elements(520));
    cp_elements(522) <= cp_elements(521);
    simple_obj_ref_1902_inst_req_0 <= cp_elements(522);
    cp_elements(523) <= type_cast_2133_inst_ack_0;
    phi_stmt_2129_req_0 <= cp_elements(523);
    cp_elements(524) <= OrReduce(cp_elements(214) & cp_elements(523));
    cp_elements(525) <= cp_elements(524);
    cp_elements(526) <= phi_stmt_2129_ack_0;
    cp_elements(527) <= false;
    cp_elements(528) <= cp_elements(527);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1929_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1929_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1929_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1942_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1942_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1942_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1961_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1961_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1961_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1980_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1980_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1980_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1999_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_1999_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_1999_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2018_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2051_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2051_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2051_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2161_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2161_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2161_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2161_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2179_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2179_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2179_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2179_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2203_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2203_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2203_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2203_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2227_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2227_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2227_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2227_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2251_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2251_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2251_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2251_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2275_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2275_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2275_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2275_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2299_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2299_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2299_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2299_root_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2317_final_offset : std_logic_vector(10 downto 0);
    signal array_obj_ref_2317_offset_scale_factor_0 : std_logic_vector(10 downto 0);
    signal array_obj_ref_2317_resized_base_address : std_logic_vector(10 downto 0);
    signal array_obj_ref_2317_root_address : std_logic_vector(10 downto 0);
    signal iNsTr_12_2390 : std_logic_vector(31 downto 0);
    signal iNsTr_16_2410 : std_logic_vector(31 downto 0);
    signal iNsTr_18_2419 : std_logic_vector(31 downto 0);
    signal iNsTr_1_1900 : std_logic_vector(31 downto 0);
    signal iNsTr_20_2429 : std_logic_vector(31 downto 0);
    signal iNsTr_2_1913 : std_logic_vector(31 downto 0);
    signal iNsTr_3_1922 : std_logic_vector(31 downto 0);
    signal iNsTr_4_2107 : std_logic_vector(31 downto 0);
    signal iNsTr_6_2117 : std_logic_vector(31 downto 0);
    signal iNsTr_9_2373 : std_logic_vector(31 downto 0);
    signal indvar_2129 : std_logic_vector(15 downto 0);
    signal ins38_2101 : std_logic_vector(63 downto 0);
    signal ins77_2367 : std_logic_vector(63 downto 0);
    signal mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2071 : std_logic_vector(63 downto 0);
    signal mask17x_xmaskedx_xmaskedx_xmasked_2076 : std_logic_vector(63 downto 0);
    signal mask22x_xmaskedx_xmaskedx_xmasked_2081 : std_logic_vector(63 downto 0);
    signal mask27x_xmaskedx_xmasked_2086 : std_logic_vector(63 downto 0);
    signal mask32x_xmasked_2091 : std_logic_vector(63 downto 0);
    signal mask37_2096 : std_logic_vector(63 downto 0);
    signal mask51_2337 : std_logic_vector(63 downto 0);
    signal mask56_2342 : std_logic_vector(63 downto 0);
    signal mask61x_xmaskedx_xmasked_2347 : std_logic_vector(63 downto 0);
    signal mask66x_xmaskedx_xmasked_2352 : std_logic_vector(63 downto 0);
    signal mask71x_xmasked_2357 : std_logic_vector(63 downto 0);
    signal mask76_2362 : std_logic_vector(63 downto 0);
    signal phitmp_2399 : std_logic_vector(15 downto 0);
    signal ptr_deref_1933_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1933_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1933_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1933_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1933_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1946_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1946_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1946_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1946_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1946_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1965_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1965_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1965_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1965_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1965_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1984_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1984_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1984_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_1984_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_1984_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2003_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2003_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2003_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2003_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2003_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2022_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2022_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2022_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2022_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2022_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2036_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2036_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2036_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2036_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2036_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2055_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2055_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2055_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2055_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2055_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2165_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2165_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2183_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2183_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2207_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2207_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2207_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2207_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2207_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2231_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2231_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2231_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2231_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2231_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2255_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2255_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2255_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2255_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2255_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2279_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2279_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2279_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2279_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2279_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2303_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2303_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2303_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2303_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2303_word_offset_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2321_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2321_resized_base_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2321_root_address : std_logic_vector(10 downto 0);
    signal ptr_deref_2321_word_address_0 : std_logic_vector(10 downto 0);
    signal ptr_deref_2321_word_offset_0 : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2160_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2160_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2178_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2178_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2202_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2202_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2226_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2226_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2250_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2250_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2274_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2274_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2298_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2298_scaled : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2316_resized : std_logic_vector(10 downto 0);
    signal simple_obj_ref_2316_scaled : std_logic_vector(10 downto 0);
    signal tmp10_1970 : std_logic_vector(63 downto 0);
    signal tmp11_1976 : std_logic_vector(63 downto 0);
    signal tmp124_1907 : std_logic_vector(31 downto 0);
    signal tmp125_1916 : std_logic_vector(31 downto 0);
    signal tmp126_1925 : std_logic_vector(7 downto 0);
    signal tmp127_1930 : std_logic_vector(31 downto 0);
    signal tmp128_1934 : std_logic_vector(7 downto 0);
    signal tmp129_1943 : std_logic_vector(31 downto 0);
    signal tmp130_1947 : std_logic_vector(7 downto 0);
    signal tmp131_1962 : std_logic_vector(31 downto 0);
    signal tmp132_1966 : std_logic_vector(7 downto 0);
    signal tmp133_1981 : std_logic_vector(31 downto 0);
    signal tmp134_1985 : std_logic_vector(7 downto 0);
    signal tmp135_2000 : std_logic_vector(31 downto 0);
    signal tmp136_2004 : std_logic_vector(7 downto 0);
    signal tmp137_2019 : std_logic_vector(31 downto 0);
    signal tmp138_2023 : std_logic_vector(7 downto 0);
    signal tmp139_2037 : std_logic_vector(7 downto 0);
    signal tmp140_2052 : std_logic_vector(31 downto 0);
    signal tmp141_2056 : std_logic_vector(7 downto 0);
    signal tmp143_2141 : std_logic_vector(31 downto 0);
    signal tmp144_2126 : std_logic_vector(31 downto 0);
    signal tmp145_2146 : std_logic_vector(0 downto 0);
    signal tmp148_2152 : std_logic_vector(31 downto 0);
    signal tmp149_2158 : std_logic_vector(31 downto 0);
    signal tmp150_2162 : std_logic_vector(31 downto 0);
    signal tmp151_2166 : std_logic_vector(7 downto 0);
    signal tmp154_2176 : std_logic_vector(31 downto 0);
    signal tmp155_2180 : std_logic_vector(31 downto 0);
    signal tmp156_2184 : std_logic_vector(7 downto 0);
    signal tmp159_2200 : std_logic_vector(31 downto 0);
    signal tmp15_1989 : std_logic_vector(63 downto 0);
    signal tmp160_2204 : std_logic_vector(31 downto 0);
    signal tmp161_2208 : std_logic_vector(7 downto 0);
    signal tmp164_2224 : std_logic_vector(31 downto 0);
    signal tmp165_2228 : std_logic_vector(31 downto 0);
    signal tmp166_2232 : std_logic_vector(7 downto 0);
    signal tmp169_2248 : std_logic_vector(31 downto 0);
    signal tmp16_1995 : std_logic_vector(63 downto 0);
    signal tmp170_2252 : std_logic_vector(31 downto 0);
    signal tmp171_2256 : std_logic_vector(7 downto 0);
    signal tmp174_2272 : std_logic_vector(31 downto 0);
    signal tmp175_2276 : std_logic_vector(31 downto 0);
    signal tmp176_2280 : std_logic_vector(7 downto 0);
    signal tmp179_2296 : std_logic_vector(31 downto 0);
    signal tmp180_2300 : std_logic_vector(31 downto 0);
    signal tmp181_2304 : std_logic_vector(7 downto 0);
    signal tmp184_2318 : std_logic_vector(31 downto 0);
    signal tmp185_2322 : std_logic_vector(7 downto 0);
    signal tmp20_2008 : std_logic_vector(63 downto 0);
    signal tmp21_2014 : std_logic_vector(63 downto 0);
    signal tmp25_2027 : std_logic_vector(63 downto 0);
    signal tmp26_2033 : std_logic_vector(63 downto 0);
    signal tmp30_2041 : std_logic_vector(63 downto 0);
    signal tmp31_2047 : std_logic_vector(63 downto 0);
    signal tmp35_2060 : std_logic_vector(63 downto 0);
    signal tmp36_2066 : std_logic_vector(63 downto 0);
    signal tmp3_1938 : std_logic_vector(63 downto 0);
    signal tmp40_2170 : std_logic_vector(63 downto 0);
    signal tmp44_2188 : std_logic_vector(63 downto 0);
    signal tmp45_2194 : std_logic_vector(63 downto 0);
    signal tmp49_2212 : std_logic_vector(63 downto 0);
    signal tmp50_2218 : std_logic_vector(63 downto 0);
    signal tmp54_2236 : std_logic_vector(63 downto 0);
    signal tmp55_2242 : std_logic_vector(63 downto 0);
    signal tmp59_2260 : std_logic_vector(63 downto 0);
    signal tmp5_1951 : std_logic_vector(63 downto 0);
    signal tmp60_2266 : std_logic_vector(63 downto 0);
    signal tmp64_2284 : std_logic_vector(63 downto 0);
    signal tmp65_2290 : std_logic_vector(63 downto 0);
    signal tmp69_2308 : std_logic_vector(63 downto 0);
    signal tmp6_1957 : std_logic_vector(63 downto 0);
    signal tmp70_2314 : std_logic_vector(63 downto 0);
    signal tmp74_2326 : std_logic_vector(63 downto 0);
    signal tmp75_2332 : std_logic_vector(63 downto 0);
    signal tmp_1903 : std_logic_vector(31 downto 0);
    signal type_cast_1955_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1993_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2012_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2031_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2045_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2064_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2110_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2124_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2133_wire : std_logic_vector(15 downto 0);
    signal type_cast_2136_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2150_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2156_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2174_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2192_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2198_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2216_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2222_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2240_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2246_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2264_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2270_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2288_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2294_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2312_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2330_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_2383_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2397_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2422_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_1929_final_offset <= "00000000111";
    array_obj_ref_1942_final_offset <= "00000000110";
    array_obj_ref_1961_final_offset <= "00000000101";
    array_obj_ref_1980_final_offset <= "00000000100";
    array_obj_ref_1999_final_offset <= "00000000011";
    array_obj_ref_2018_final_offset <= "00000000010";
    array_obj_ref_2051_final_offset <= "00000000001";
    array_obj_ref_2161_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2179_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2203_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2227_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2251_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2275_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2299_offset_scale_factor_0 <= "00000000001";
    array_obj_ref_2317_offset_scale_factor_0 <= "00000000001";
    iNsTr_12_2390 <= "00000000000000000000000000000000";
    iNsTr_16_2410 <= "00000000000000000000000000000000";
    iNsTr_18_2419 <= "00000000000000000000000000000000";
    iNsTr_1_1900 <= "00000000000000000000000000000000";
    iNsTr_20_2429 <= "00000000000000000000000000000000";
    iNsTr_2_1913 <= "00000000000000000000000000000000";
    iNsTr_3_1922 <= "00000000000000000000000000000000";
    iNsTr_4_2107 <= "00000000000000000000000000000000";
    iNsTr_6_2117 <= "00000000000000000000000000000000";
    iNsTr_9_2373 <= "00000000000000000000000000000000";
    ptr_deref_1933_word_offset_0 <= "00000000000";
    ptr_deref_1946_word_offset_0 <= "00000000000";
    ptr_deref_1965_word_offset_0 <= "00000000000";
    ptr_deref_1984_word_offset_0 <= "00000000000";
    ptr_deref_2003_word_offset_0 <= "00000000000";
    ptr_deref_2022_word_offset_0 <= "00000000000";
    ptr_deref_2036_word_offset_0 <= "00000000000";
    ptr_deref_2055_word_offset_0 <= "00000000000";
    ptr_deref_2165_word_offset_0 <= "00000000000";
    ptr_deref_2183_word_offset_0 <= "00000000000";
    ptr_deref_2207_word_offset_0 <= "00000000000";
    ptr_deref_2231_word_offset_0 <= "00000000000";
    ptr_deref_2255_word_offset_0 <= "00000000000";
    ptr_deref_2279_word_offset_0 <= "00000000000";
    ptr_deref_2303_word_offset_0 <= "00000000000";
    ptr_deref_2321_word_offset_0 <= "00000000000";
    type_cast_1955_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_1974_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_1993_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2012_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2031_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2045_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2064_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2110_wire_constant <= "11111111";
    type_cast_2124_wire_constant <= "11111111111111111111111111111111";
    type_cast_2136_wire_constant <= "0000000000000001";
    type_cast_2150_wire_constant <= "00000000000000000000000000000011";
    type_cast_2156_wire_constant <= "00000000000000000000000000000111";
    type_cast_2174_wire_constant <= "00000000000000000000000000000110";
    type_cast_2192_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    type_cast_2198_wire_constant <= "00000000000000000000000000000101";
    type_cast_2216_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    type_cast_2222_wire_constant <= "00000000000000000000000000000100";
    type_cast_2240_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    type_cast_2246_wire_constant <= "00000000000000000000000000000011";
    type_cast_2264_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    type_cast_2270_wire_constant <= "00000000000000000000000000000010";
    type_cast_2288_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    type_cast_2294_wire_constant <= "00000000000000000000000000000001";
    type_cast_2312_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    type_cast_2330_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    type_cast_2383_wire_constant <= "00000000";
    type_cast_2397_wire_constant <= "0000000000000001";
    type_cast_2422_wire_constant <= "00000001";
    phi_stmt_2129: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2133_wire & type_cast_2136_wire_constant;
      req <= phi_stmt_2129_req_0 & phi_stmt_2129_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2129_ack_0,
          idata => idata,
          odata => indvar_2129,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2129
    array_obj_ref_1929_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_1929_resized_base_address, req => array_obj_ref_1929_base_resize_req_0, ack => array_obj_ref_1929_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1929_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1929_root_address, dout => tmp127_1930, req => array_obj_ref_1929_final_reg_req_0, ack => array_obj_ref_1929_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1942_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_1942_resized_base_address, req => array_obj_ref_1942_base_resize_req_0, ack => array_obj_ref_1942_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1942_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1942_root_address, dout => tmp129_1943, req => array_obj_ref_1942_final_reg_req_0, ack => array_obj_ref_1942_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1961_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_1961_resized_base_address, req => array_obj_ref_1961_base_resize_req_0, ack => array_obj_ref_1961_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1961_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1961_root_address, dout => tmp131_1962, req => array_obj_ref_1961_final_reg_req_0, ack => array_obj_ref_1961_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1980_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_1980_resized_base_address, req => array_obj_ref_1980_base_resize_req_0, ack => array_obj_ref_1980_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1980_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1980_root_address, dout => tmp133_1981, req => array_obj_ref_1980_final_reg_req_0, ack => array_obj_ref_1980_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1999_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_1999_resized_base_address, req => array_obj_ref_1999_base_resize_req_0, ack => array_obj_ref_1999_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1999_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1999_root_address, dout => tmp135_2000, req => array_obj_ref_1999_final_reg_req_0, ack => array_obj_ref_1999_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2018_resized_base_address, req => array_obj_ref_2018_base_resize_req_0, ack => array_obj_ref_2018_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2018_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2018_root_address, dout => tmp137_2019, req => array_obj_ref_2018_final_reg_req_0, ack => array_obj_ref_2018_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2051_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2051_resized_base_address, req => array_obj_ref_2051_base_resize_req_0, ack => array_obj_ref_2051_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2051_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2051_root_address, dout => tmp140_2052, req => array_obj_ref_2051_final_reg_req_0, ack => array_obj_ref_2051_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2161_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2161_resized_base_address, req => array_obj_ref_2161_base_resize_req_0, ack => array_obj_ref_2161_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2161_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2161_root_address, dout => tmp150_2162, req => array_obj_ref_2161_final_reg_req_0, ack => array_obj_ref_2161_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2161_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp149_2158, dout => simple_obj_ref_2160_resized, req => array_obj_ref_2161_index_0_resize_req_0, ack => array_obj_ref_2161_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2161_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2160_scaled, dout => array_obj_ref_2161_final_offset, req => array_obj_ref_2161_offset_inst_req_0, ack => array_obj_ref_2161_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2179_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2179_resized_base_address, req => array_obj_ref_2179_base_resize_req_0, ack => array_obj_ref_2179_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2179_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2179_root_address, dout => tmp155_2180, req => array_obj_ref_2179_final_reg_req_0, ack => array_obj_ref_2179_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2179_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp154_2176, dout => simple_obj_ref_2178_resized, req => array_obj_ref_2179_index_0_resize_req_0, ack => array_obj_ref_2179_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2179_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2178_scaled, dout => array_obj_ref_2179_final_offset, req => array_obj_ref_2179_offset_inst_req_0, ack => array_obj_ref_2179_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2203_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2203_resized_base_address, req => array_obj_ref_2203_base_resize_req_0, ack => array_obj_ref_2203_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2203_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2203_root_address, dout => tmp160_2204, req => array_obj_ref_2203_final_reg_req_0, ack => array_obj_ref_2203_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2203_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp159_2200, dout => simple_obj_ref_2202_resized, req => array_obj_ref_2203_index_0_resize_req_0, ack => array_obj_ref_2203_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2203_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2202_scaled, dout => array_obj_ref_2203_final_offset, req => array_obj_ref_2203_offset_inst_req_0, ack => array_obj_ref_2203_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2227_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2227_resized_base_address, req => array_obj_ref_2227_base_resize_req_0, ack => array_obj_ref_2227_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2227_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2227_root_address, dout => tmp165_2228, req => array_obj_ref_2227_final_reg_req_0, ack => array_obj_ref_2227_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2227_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp164_2224, dout => simple_obj_ref_2226_resized, req => array_obj_ref_2227_index_0_resize_req_0, ack => array_obj_ref_2227_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2227_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2226_scaled, dout => array_obj_ref_2227_final_offset, req => array_obj_ref_2227_offset_inst_req_0, ack => array_obj_ref_2227_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2251_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2251_resized_base_address, req => array_obj_ref_2251_base_resize_req_0, ack => array_obj_ref_2251_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2251_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2251_root_address, dout => tmp170_2252, req => array_obj_ref_2251_final_reg_req_0, ack => array_obj_ref_2251_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2251_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp169_2248, dout => simple_obj_ref_2250_resized, req => array_obj_ref_2251_index_0_resize_req_0, ack => array_obj_ref_2251_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2251_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2250_scaled, dout => array_obj_ref_2251_final_offset, req => array_obj_ref_2251_offset_inst_req_0, ack => array_obj_ref_2251_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2275_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2275_resized_base_address, req => array_obj_ref_2275_base_resize_req_0, ack => array_obj_ref_2275_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2275_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2275_root_address, dout => tmp175_2276, req => array_obj_ref_2275_final_reg_req_0, ack => array_obj_ref_2275_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2275_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp174_2272, dout => simple_obj_ref_2274_resized, req => array_obj_ref_2275_index_0_resize_req_0, ack => array_obj_ref_2275_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2275_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2274_scaled, dout => array_obj_ref_2275_final_offset, req => array_obj_ref_2275_offset_inst_req_0, ack => array_obj_ref_2275_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2299_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2299_resized_base_address, req => array_obj_ref_2299_base_resize_req_0, ack => array_obj_ref_2299_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2299_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2299_root_address, dout => tmp180_2300, req => array_obj_ref_2299_final_reg_req_0, ack => array_obj_ref_2299_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2299_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp179_2296, dout => simple_obj_ref_2298_resized, req => array_obj_ref_2299_index_0_resize_req_0, ack => array_obj_ref_2299_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2299_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2298_scaled, dout => array_obj_ref_2299_final_offset, req => array_obj_ref_2299_offset_inst_req_0, ack => array_obj_ref_2299_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2317_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => array_obj_ref_2317_resized_base_address, req => array_obj_ref_2317_base_resize_req_0, ack => array_obj_ref_2317_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2317_final_reg: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2317_root_address, dout => tmp184_2318, req => array_obj_ref_2317_final_reg_req_0, ack => array_obj_ref_2317_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2317_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp148_2152, dout => simple_obj_ref_2316_resized, req => array_obj_ref_2317_index_0_resize_req_0, ack => array_obj_ref_2317_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2317_offset_inst: RegisterBase --
      generic map(in_data_width => 11,out_data_width => 11, flow_through => true ) 
      port map( din => simple_obj_ref_2316_scaled, dout => array_obj_ref_2317_final_offset, req => array_obj_ref_2317_offset_inst_req_0, ack => array_obj_ref_2317_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1933_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp127_1930, dout => ptr_deref_1933_resized_base_address, req => ptr_deref_1933_base_resize_req_0, ack => ptr_deref_1933_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1946_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp129_1943, dout => ptr_deref_1946_resized_base_address, req => ptr_deref_1946_base_resize_req_0, ack => ptr_deref_1946_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1965_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp131_1962, dout => ptr_deref_1965_resized_base_address, req => ptr_deref_1965_base_resize_req_0, ack => ptr_deref_1965_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1984_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp133_1981, dout => ptr_deref_1984_resized_base_address, req => ptr_deref_1984_base_resize_req_0, ack => ptr_deref_1984_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2003_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp135_2000, dout => ptr_deref_2003_resized_base_address, req => ptr_deref_2003_base_resize_req_0, ack => ptr_deref_2003_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2022_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp137_2019, dout => ptr_deref_2022_resized_base_address, req => ptr_deref_2022_base_resize_req_0, ack => ptr_deref_2022_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2036_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp124_1907, dout => ptr_deref_2036_resized_base_address, req => ptr_deref_2036_base_resize_req_0, ack => ptr_deref_2036_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2055_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp140_2052, dout => ptr_deref_2055_resized_base_address, req => ptr_deref_2055_base_resize_req_0, ack => ptr_deref_2055_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2165_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp150_2162, dout => ptr_deref_2165_resized_base_address, req => ptr_deref_2165_base_resize_req_0, ack => ptr_deref_2165_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2183_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp155_2180, dout => ptr_deref_2183_resized_base_address, req => ptr_deref_2183_base_resize_req_0, ack => ptr_deref_2183_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2207_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp160_2204, dout => ptr_deref_2207_resized_base_address, req => ptr_deref_2207_base_resize_req_0, ack => ptr_deref_2207_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2231_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp165_2228, dout => ptr_deref_2231_resized_base_address, req => ptr_deref_2231_base_resize_req_0, ack => ptr_deref_2231_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2255_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp170_2252, dout => ptr_deref_2255_resized_base_address, req => ptr_deref_2255_base_resize_req_0, ack => ptr_deref_2255_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2279_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp175_2276, dout => ptr_deref_2279_resized_base_address, req => ptr_deref_2279_base_resize_req_0, ack => ptr_deref_2279_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2303_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp180_2300, dout => ptr_deref_2303_resized_base_address, req => ptr_deref_2303_base_resize_req_0, ack => ptr_deref_2303_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2321_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 11, flow_through => true ) 
      port map( din => tmp184_2318, dout => ptr_deref_2321_resized_base_address, req => ptr_deref_2321_base_resize_req_0, ack => ptr_deref_2321_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1906_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1903, dout => tmp124_1907, req => type_cast_1906_inst_req_0, ack => type_cast_1906_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1937_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp128_1934, dout => tmp3_1938, req => type_cast_1937_inst_req_0, ack => type_cast_1937_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1950_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp130_1947, dout => tmp5_1951, req => type_cast_1950_inst_req_0, ack => type_cast_1950_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1969_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp132_1966, dout => tmp10_1970, req => type_cast_1969_inst_req_0, ack => type_cast_1969_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1988_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp134_1985, dout => tmp15_1989, req => type_cast_1988_inst_req_0, ack => type_cast_1988_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2007_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp136_2004, dout => tmp20_2008, req => type_cast_2007_inst_req_0, ack => type_cast_2007_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2026_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp138_2023, dout => tmp25_2027, req => type_cast_2026_inst_req_0, ack => type_cast_2026_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2040_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp139_2037, dout => tmp30_2041, req => type_cast_2040_inst_req_0, ack => type_cast_2040_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2059_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp141_2056, dout => tmp35_2060, req => type_cast_2059_inst_req_0, ack => type_cast_2059_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2133_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => phitmp_2399, dout => type_cast_2133_wire, req => type_cast_2133_inst_req_0, ack => type_cast_2133_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2140_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => indvar_2129, dout => tmp143_2141, req => type_cast_2140_inst_req_0, ack => type_cast_2140_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2169_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp151_2166, dout => tmp40_2170, req => type_cast_2169_inst_req_0, ack => type_cast_2169_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2187_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp156_2184, dout => tmp44_2188, req => type_cast_2187_inst_req_0, ack => type_cast_2187_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2211_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp161_2208, dout => tmp49_2212, req => type_cast_2211_inst_req_0, ack => type_cast_2211_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2235_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp166_2232, dout => tmp54_2236, req => type_cast_2235_inst_req_0, ack => type_cast_2235_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2259_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp171_2256, dout => tmp59_2260, req => type_cast_2259_inst_req_0, ack => type_cast_2259_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2283_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp176_2280, dout => tmp64_2284, req => type_cast_2283_inst_req_0, ack => type_cast_2283_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2307_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp181_2304, dout => tmp69_2308, req => type_cast_2307_inst_req_0, ack => type_cast_2307_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2325_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 64, flow_through => false ) 
      port map( din => tmp185_2322, dout => tmp74_2326, req => type_cast_2325_inst_req_0, ack => type_cast_2325_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2161_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2161_index_0_rename_ack_0 <= array_obj_ref_2161_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2160_resized;
      simple_obj_ref_2160_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2179_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2179_index_0_rename_ack_0 <= array_obj_ref_2179_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2178_resized;
      simple_obj_ref_2178_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2203_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2203_index_0_rename_ack_0 <= array_obj_ref_2203_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2202_resized;
      simple_obj_ref_2202_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2227_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2227_index_0_rename_ack_0 <= array_obj_ref_2227_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2226_resized;
      simple_obj_ref_2226_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2251_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2251_index_0_rename_ack_0 <= array_obj_ref_2251_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2250_resized;
      simple_obj_ref_2250_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2275_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2275_index_0_rename_ack_0 <= array_obj_ref_2275_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2274_resized;
      simple_obj_ref_2274_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2299_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2299_index_0_rename_ack_0 <= array_obj_ref_2299_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2298_resized;
      simple_obj_ref_2298_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    array_obj_ref_2317_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      array_obj_ref_2317_index_0_rename_ack_0 <= array_obj_ref_2317_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2316_resized;
      simple_obj_ref_2316_scaled <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1933_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1933_addr_0_ack_0 <= ptr_deref_1933_addr_0_req_0;
      aggregated_sig <= ptr_deref_1933_root_address;
      ptr_deref_1933_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1933_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1933_gather_scatter_ack_0 <= ptr_deref_1933_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1933_data_0;
      tmp128_1934 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1933_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1933_root_address_inst_ack_0 <= ptr_deref_1933_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1933_resized_base_address;
      ptr_deref_1933_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1946_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1946_addr_0_ack_0 <= ptr_deref_1946_addr_0_req_0;
      aggregated_sig <= ptr_deref_1946_root_address;
      ptr_deref_1946_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1946_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1946_gather_scatter_ack_0 <= ptr_deref_1946_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1946_data_0;
      tmp130_1947 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1946_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1946_root_address_inst_ack_0 <= ptr_deref_1946_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1946_resized_base_address;
      ptr_deref_1946_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1965_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1965_addr_0_ack_0 <= ptr_deref_1965_addr_0_req_0;
      aggregated_sig <= ptr_deref_1965_root_address;
      ptr_deref_1965_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1965_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1965_gather_scatter_ack_0 <= ptr_deref_1965_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1965_data_0;
      tmp132_1966 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1965_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1965_root_address_inst_ack_0 <= ptr_deref_1965_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1965_resized_base_address;
      ptr_deref_1965_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1984_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1984_addr_0_ack_0 <= ptr_deref_1984_addr_0_req_0;
      aggregated_sig <= ptr_deref_1984_root_address;
      ptr_deref_1984_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_1984_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1984_gather_scatter_ack_0 <= ptr_deref_1984_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1984_data_0;
      tmp134_1985 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1984_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_1984_root_address_inst_ack_0 <= ptr_deref_1984_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1984_resized_base_address;
      ptr_deref_1984_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2003_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2003_addr_0_ack_0 <= ptr_deref_2003_addr_0_req_0;
      aggregated_sig <= ptr_deref_2003_root_address;
      ptr_deref_2003_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2003_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2003_gather_scatter_ack_0 <= ptr_deref_2003_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2003_data_0;
      tmp136_2004 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2003_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2003_root_address_inst_ack_0 <= ptr_deref_2003_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2003_resized_base_address;
      ptr_deref_2003_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2022_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2022_addr_0_ack_0 <= ptr_deref_2022_addr_0_req_0;
      aggregated_sig <= ptr_deref_2022_root_address;
      ptr_deref_2022_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2022_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2022_gather_scatter_ack_0 <= ptr_deref_2022_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2022_data_0;
      tmp138_2023 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2022_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2022_root_address_inst_ack_0 <= ptr_deref_2022_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2022_resized_base_address;
      ptr_deref_2022_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2036_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2036_addr_0_ack_0 <= ptr_deref_2036_addr_0_req_0;
      aggregated_sig <= ptr_deref_2036_root_address;
      ptr_deref_2036_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2036_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2036_gather_scatter_ack_0 <= ptr_deref_2036_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2036_data_0;
      tmp139_2037 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2036_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2036_root_address_inst_ack_0 <= ptr_deref_2036_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2036_resized_base_address;
      ptr_deref_2036_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2055_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2055_addr_0_ack_0 <= ptr_deref_2055_addr_0_req_0;
      aggregated_sig <= ptr_deref_2055_root_address;
      ptr_deref_2055_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2055_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2055_gather_scatter_ack_0 <= ptr_deref_2055_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2055_data_0;
      tmp141_2056 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2055_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2055_root_address_inst_ack_0 <= ptr_deref_2055_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2055_resized_base_address;
      ptr_deref_2055_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2165_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2165_addr_0_ack_0 <= ptr_deref_2165_addr_0_req_0;
      aggregated_sig <= ptr_deref_2165_root_address;
      ptr_deref_2165_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2165_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2165_gather_scatter_ack_0 <= ptr_deref_2165_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2165_data_0;
      tmp151_2166 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2165_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2165_root_address_inst_ack_0 <= ptr_deref_2165_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2165_resized_base_address;
      ptr_deref_2165_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2183_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2183_addr_0_ack_0 <= ptr_deref_2183_addr_0_req_0;
      aggregated_sig <= ptr_deref_2183_root_address;
      ptr_deref_2183_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2183_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2183_gather_scatter_ack_0 <= ptr_deref_2183_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2183_data_0;
      tmp156_2184 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2183_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2183_root_address_inst_ack_0 <= ptr_deref_2183_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2183_resized_base_address;
      ptr_deref_2183_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2207_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2207_addr_0_ack_0 <= ptr_deref_2207_addr_0_req_0;
      aggregated_sig <= ptr_deref_2207_root_address;
      ptr_deref_2207_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2207_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2207_gather_scatter_ack_0 <= ptr_deref_2207_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2207_data_0;
      tmp161_2208 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2207_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2207_root_address_inst_ack_0 <= ptr_deref_2207_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2207_resized_base_address;
      ptr_deref_2207_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2231_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2231_addr_0_ack_0 <= ptr_deref_2231_addr_0_req_0;
      aggregated_sig <= ptr_deref_2231_root_address;
      ptr_deref_2231_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2231_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2231_gather_scatter_ack_0 <= ptr_deref_2231_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2231_data_0;
      tmp166_2232 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2231_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2231_root_address_inst_ack_0 <= ptr_deref_2231_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2231_resized_base_address;
      ptr_deref_2231_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2255_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2255_addr_0_ack_0 <= ptr_deref_2255_addr_0_req_0;
      aggregated_sig <= ptr_deref_2255_root_address;
      ptr_deref_2255_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2255_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2255_gather_scatter_ack_0 <= ptr_deref_2255_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2255_data_0;
      tmp171_2256 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2255_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2255_root_address_inst_ack_0 <= ptr_deref_2255_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2255_resized_base_address;
      ptr_deref_2255_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2279_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2279_addr_0_ack_0 <= ptr_deref_2279_addr_0_req_0;
      aggregated_sig <= ptr_deref_2279_root_address;
      ptr_deref_2279_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2279_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2279_gather_scatter_ack_0 <= ptr_deref_2279_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2279_data_0;
      tmp176_2280 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2279_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2279_root_address_inst_ack_0 <= ptr_deref_2279_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2279_resized_base_address;
      ptr_deref_2279_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2303_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2303_addr_0_ack_0 <= ptr_deref_2303_addr_0_req_0;
      aggregated_sig <= ptr_deref_2303_root_address;
      ptr_deref_2303_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2303_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2303_gather_scatter_ack_0 <= ptr_deref_2303_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2303_data_0;
      tmp181_2304 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2303_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2303_root_address_inst_ack_0 <= ptr_deref_2303_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2303_resized_base_address;
      ptr_deref_2303_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2321_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2321_addr_0_ack_0 <= ptr_deref_2321_addr_0_req_0;
      aggregated_sig <= ptr_deref_2321_root_address;
      ptr_deref_2321_word_address_0 <= aggregated_sig(10 downto 0);
      --
    end Block;
    ptr_deref_2321_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2321_gather_scatter_ack_0 <= ptr_deref_2321_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2321_data_0;
      tmp185_2322 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2321_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(10 downto 0); --
    begin -- 
      ptr_deref_2321_root_address_inst_ack_0 <= ptr_deref_2321_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2321_resized_base_address;
      ptr_deref_2321_root_address <= aggregated_sig(10 downto 0);
      --
    end Block;
    if_stmt_2374_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp145_2146;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2374_branch_req_0,
          ack0 => if_stmt_2374_branch_ack_0,
          ack1 => if_stmt_2374_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1929_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1929_resized_base_address;
      array_obj_ref_1929_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000111",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1929_root_address_inst_req_0,
          ackL => array_obj_ref_1929_root_address_inst_ack_0,
          reqR => array_obj_ref_1929_root_address_inst_req_1,
          ackR => array_obj_ref_1929_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1942_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1942_resized_base_address;
      array_obj_ref_1942_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000110",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1942_root_address_inst_req_0,
          ackL => array_obj_ref_1942_root_address_inst_ack_0,
          reqR => array_obj_ref_1942_root_address_inst_req_1,
          ackR => array_obj_ref_1942_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1961_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1961_resized_base_address;
      array_obj_ref_1961_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000101",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1961_root_address_inst_req_0,
          ackL => array_obj_ref_1961_root_address_inst_ack_0,
          reqR => array_obj_ref_1961_root_address_inst_req_1,
          ackR => array_obj_ref_1961_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1980_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1980_resized_base_address;
      array_obj_ref_1980_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000100",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1980_root_address_inst_req_0,
          ackL => array_obj_ref_1980_root_address_inst_ack_0,
          reqR => array_obj_ref_1980_root_address_inst_req_1,
          ackR => array_obj_ref_1980_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1999_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1999_resized_base_address;
      array_obj_ref_1999_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000011",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1999_root_address_inst_req_0,
          ackL => array_obj_ref_1999_root_address_inst_ack_0,
          reqR => array_obj_ref_1999_root_address_inst_req_1,
          ackR => array_obj_ref_1999_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_2018_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2018_resized_base_address;
      array_obj_ref_2018_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000010",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2018_root_address_inst_req_0,
          ackL => array_obj_ref_2018_root_address_inst_ack_0,
          reqR => array_obj_ref_2018_root_address_inst_req_1,
          ackR => array_obj_ref_2018_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_2051_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2051_resized_base_address;
      array_obj_ref_2051_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000000001",
          constant_width => 11,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2051_root_address_inst_req_0,
          ackL => array_obj_ref_2051_root_address_inst_ack_0,
          reqR => array_obj_ref_2051_root_address_inst_req_1,
          ackR => array_obj_ref_2051_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_2161_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2161_final_offset & array_obj_ref_2161_resized_base_address;
      array_obj_ref_2161_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2161_root_address_inst_req_0,
          ackL => array_obj_ref_2161_root_address_inst_ack_0,
          reqR => array_obj_ref_2161_root_address_inst_req_1,
          ackR => array_obj_ref_2161_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_2179_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2179_final_offset & array_obj_ref_2179_resized_base_address;
      array_obj_ref_2179_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2179_root_address_inst_req_0,
          ackL => array_obj_ref_2179_root_address_inst_ack_0,
          reqR => array_obj_ref_2179_root_address_inst_req_1,
          ackR => array_obj_ref_2179_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_2203_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2203_final_offset & array_obj_ref_2203_resized_base_address;
      array_obj_ref_2203_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2203_root_address_inst_req_0,
          ackL => array_obj_ref_2203_root_address_inst_ack_0,
          reqR => array_obj_ref_2203_root_address_inst_req_1,
          ackR => array_obj_ref_2203_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_2227_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2227_final_offset & array_obj_ref_2227_resized_base_address;
      array_obj_ref_2227_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2227_root_address_inst_req_0,
          ackL => array_obj_ref_2227_root_address_inst_ack_0,
          reqR => array_obj_ref_2227_root_address_inst_req_1,
          ackR => array_obj_ref_2227_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_2251_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2251_final_offset & array_obj_ref_2251_resized_base_address;
      array_obj_ref_2251_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2251_root_address_inst_req_0,
          ackL => array_obj_ref_2251_root_address_inst_ack_0,
          reqR => array_obj_ref_2251_root_address_inst_req_1,
          ackR => array_obj_ref_2251_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_2275_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2275_final_offset & array_obj_ref_2275_resized_base_address;
      array_obj_ref_2275_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2275_root_address_inst_req_0,
          ackL => array_obj_ref_2275_root_address_inst_ack_0,
          reqR => array_obj_ref_2275_root_address_inst_req_1,
          ackR => array_obj_ref_2275_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_2299_root_address_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2299_final_offset & array_obj_ref_2299_resized_base_address;
      array_obj_ref_2299_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2299_root_address_inst_req_0,
          ackL => array_obj_ref_2299_root_address_inst_ack_0,
          reqR => array_obj_ref_2299_root_address_inst_req_1,
          ackR => array_obj_ref_2299_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_2317_root_address_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2317_final_offset & array_obj_ref_2317_resized_base_address;
      array_obj_ref_2317_root_address <= data_out(10 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2317_root_address_inst_req_0,
          ackL => array_obj_ref_2317_root_address_inst_ack_0,
          reqR => array_obj_ref_2317_root_address_inst_req_1,
          ackR => array_obj_ref_2317_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1956_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_1951;
      tmp6_1957 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1956_inst_req_0,
          ackL => binary_1956_inst_ack_0,
          reqR => binary_1956_inst_req_1,
          ackR => binary_1956_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1975_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp10_1970;
      tmp11_1976 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1975_inst_req_0,
          ackL => binary_1975_inst_ack_0,
          reqR => binary_1975_inst_req_1,
          ackR => binary_1975_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1994_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_1989;
      tmp16_1995 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1994_inst_req_0,
          ackL => binary_1994_inst_ack_0,
          reqR => binary_1994_inst_req_1,
          ackR => binary_1994_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_2013_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_2008;
      tmp21_2014 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2013_inst_req_0,
          ackL => binary_2013_inst_ack_0,
          reqR => binary_2013_inst_req_1,
          ackR => binary_2013_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_2032_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp25_2027;
      tmp26_2033 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2032_inst_req_0,
          ackL => binary_2032_inst_ack_0,
          reqR => binary_2032_inst_req_1,
          ackR => binary_2032_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_2046_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_2041;
      tmp31_2047 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2046_inst_req_0,
          ackL => binary_2046_inst_ack_0,
          reqR => binary_2046_inst_req_1,
          ackR => binary_2046_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_2065_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp35_2060;
      tmp36_2066 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2065_inst_req_0,
          ackL => binary_2065_inst_ack_0,
          reqR => binary_2065_inst_req_1,
          ackR => binary_2065_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_2070_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp6_1957 & tmp3_1938;
      mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2071 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2070_inst_req_0,
          ackL => binary_2070_inst_ack_0,
          reqR => binary_2070_inst_req_1,
          ackR => binary_2070_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_2075_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask12x_xmaskedx_xmaskedx_xmaskedx_xmasked_2071 & tmp11_1976;
      mask17x_xmaskedx_xmaskedx_xmasked_2076 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2075_inst_req_0,
          ackL => binary_2075_inst_ack_0,
          reqR => binary_2075_inst_req_1,
          ackR => binary_2075_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_2080_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask17x_xmaskedx_xmaskedx_xmasked_2076 & tmp16_1995;
      mask22x_xmaskedx_xmaskedx_xmasked_2081 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2080_inst_req_0,
          ackL => binary_2080_inst_ack_0,
          reqR => binary_2080_inst_req_1,
          ackR => binary_2080_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_2085_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask22x_xmaskedx_xmaskedx_xmasked_2081 & tmp21_2014;
      mask27x_xmaskedx_xmasked_2086 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2085_inst_req_0,
          ackL => binary_2085_inst_ack_0,
          reqR => binary_2085_inst_req_1,
          ackR => binary_2085_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_2090_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask27x_xmaskedx_xmasked_2086 & tmp26_2033;
      mask32x_xmasked_2091 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2090_inst_req_0,
          ackL => binary_2090_inst_ack_0,
          reqR => binary_2090_inst_req_1,
          ackR => binary_2090_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_2095_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask32x_xmasked_2091 & tmp31_2047;
      mask37_2096 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2095_inst_req_0,
          ackL => binary_2095_inst_ack_0,
          reqR => binary_2095_inst_req_1,
          ackR => binary_2095_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_2100_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask37_2096 & tmp36_2066;
      ins38_2101 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2100_inst_req_0,
          ackL => binary_2100_inst_ack_0,
          reqR => binary_2100_inst_req_1,
          ackR => binary_2100_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_2125_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp125_1916;
      tmp144_2126 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2125_inst_req_0,
          ackL => binary_2125_inst_ack_0,
          reqR => binary_2125_inst_req_1,
          ackR => binary_2125_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_2145_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp143_2141 & tmp144_2126;
      tmp145_2146 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2145_inst_req_0,
          ackL => binary_2145_inst_ack_0,
          reqR => binary_2145_inst_req_1,
          ackR => binary_2145_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_2151_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp143_2141;
      tmp148_2152 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2151_inst_req_0,
          ackL => binary_2151_inst_ack_0,
          reqR => binary_2151_inst_req_1,
          ackR => binary_2151_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_2157_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp149_2158 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2157_inst_req_0,
          ackL => binary_2157_inst_ack_0,
          reqR => binary_2157_inst_req_1,
          ackR => binary_2157_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_2175_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp154_2176 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2175_inst_req_0,
          ackL => binary_2175_inst_ack_0,
          reqR => binary_2175_inst_req_1,
          ackR => binary_2175_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_2193_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_2188;
      tmp45_2194 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2193_inst_req_0,
          ackL => binary_2193_inst_ack_0,
          reqR => binary_2193_inst_req_1,
          ackR => binary_2193_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_2199_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp159_2200 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2199_inst_req_0,
          ackL => binary_2199_inst_ack_0,
          reqR => binary_2199_inst_req_1,
          ackR => binary_2199_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_2217_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_2212;
      tmp50_2218 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2217_inst_req_0,
          ackL => binary_2217_inst_ack_0,
          reqR => binary_2217_inst_req_1,
          ackR => binary_2217_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_2223_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp164_2224 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2223_inst_req_0,
          ackL => binary_2223_inst_ack_0,
          reqR => binary_2223_inst_req_1,
          ackR => binary_2223_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_2241_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp54_2236;
      tmp55_2242 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2241_inst_req_0,
          ackL => binary_2241_inst_ack_0,
          reqR => binary_2241_inst_req_1,
          ackR => binary_2241_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_2247_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp169_2248 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2247_inst_req_0,
          ackL => binary_2247_inst_ack_0,
          reqR => binary_2247_inst_req_1,
          ackR => binary_2247_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_2265_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp59_2260;
      tmp60_2266 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2265_inst_req_0,
          ackL => binary_2265_inst_ack_0,
          reqR => binary_2265_inst_req_1,
          ackR => binary_2265_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_2271_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp174_2272 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2271_inst_req_0,
          ackL => binary_2271_inst_ack_0,
          reqR => binary_2271_inst_req_1,
          ackR => binary_2271_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_2289_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp64_2284;
      tmp65_2290 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2289_inst_req_0,
          ackL => binary_2289_inst_ack_0,
          reqR => binary_2289_inst_req_1,
          ackR => binary_2289_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_2295_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp148_2152;
      tmp179_2296 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2295_inst_req_0,
          ackL => binary_2295_inst_ack_0,
          reqR => binary_2295_inst_req_1,
          ackR => binary_2295_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_2313_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp69_2308;
      tmp70_2314 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2313_inst_req_0,
          ackL => binary_2313_inst_ack_0,
          reqR => binary_2313_inst_req_1,
          ackR => binary_2313_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_2331_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp74_2326;
      tmp75_2332 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2331_inst_req_0,
          ackL => binary_2331_inst_ack_0,
          reqR => binary_2331_inst_req_1,
          ackR => binary_2331_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_2336_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp45_2194 & tmp40_2170;
      mask51_2337 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2336_inst_req_0,
          ackL => binary_2336_inst_ack_0,
          reqR => binary_2336_inst_req_1,
          ackR => binary_2336_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_2341_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask51_2337 & tmp50_2218;
      mask56_2342 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2341_inst_req_0,
          ackL => binary_2341_inst_ack_0,
          reqR => binary_2341_inst_req_1,
          ackR => binary_2341_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_2346_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask56_2342 & tmp55_2242;
      mask61x_xmaskedx_xmasked_2347 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2346_inst_req_0,
          ackL => binary_2346_inst_ack_0,
          reqR => binary_2346_inst_req_1,
          ackR => binary_2346_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_2351_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask61x_xmaskedx_xmasked_2347 & tmp60_2266;
      mask66x_xmaskedx_xmasked_2352 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2351_inst_req_0,
          ackL => binary_2351_inst_ack_0,
          reqR => binary_2351_inst_req_1,
          ackR => binary_2351_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_2356_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask66x_xmaskedx_xmasked_2352 & tmp65_2290;
      mask71x_xmasked_2357 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2356_inst_req_0,
          ackL => binary_2356_inst_ack_0,
          reqR => binary_2356_inst_req_1,
          ackR => binary_2356_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_2361_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask71x_xmasked_2357 & tmp70_2314;
      mask76_2362 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2361_inst_req_0,
          ackL => binary_2361_inst_ack_0,
          reqR => binary_2361_inst_req_1,
          ackR => binary_2361_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : binary_2366_inst 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= mask76_2362 & tmp75_2332;
      ins77_2367 <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 64, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2366_inst_req_0,
          ackL => binary_2366_inst_ack_0,
          reqR => binary_2366_inst_req_1,
          ackR => binary_2366_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : binary_2398_inst 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_2129;
      phitmp_2399 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2398_inst_req_0,
          ackL => binary_2398_inst_ack_0,
          reqR => binary_2398_inst_req_1,
          ackR => binary_2398_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared load operator group (0) : ptr_deref_1933_load_0 ptr_deref_2165_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1933_load_0_req_0;
      reqL(0) <= ptr_deref_2165_load_0_req_0;
      ptr_deref_1933_load_0_ack_0 <= ackL(1);
      ptr_deref_2165_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1933_load_0_req_1;
      reqR(0) <= ptr_deref_2165_load_0_req_1;
      ptr_deref_1933_load_0_ack_1 <= ackR(1);
      ptr_deref_2165_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1933_word_address_0 & ptr_deref_2165_word_address_0;
      ptr_deref_1933_data_0 <= data_out(15 downto 8);
      ptr_deref_2165_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(7),
          mack => memory_space_3_lr_ack(7),
          maddr => memory_space_3_lr_addr(87 downto 77),
          mtag => memory_space_3_lr_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(7),
          mack => memory_space_3_lc_ack(7),
          mdata => memory_space_3_lc_data(63 downto 56),
          mtag => memory_space_3_lc_tag(15 downto 14),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1946_load_0 ptr_deref_2183_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1946_load_0_req_0;
      reqL(0) <= ptr_deref_2183_load_0_req_0;
      ptr_deref_1946_load_0_ack_0 <= ackL(1);
      ptr_deref_2183_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1946_load_0_req_1;
      reqR(0) <= ptr_deref_2183_load_0_req_1;
      ptr_deref_1946_load_0_ack_1 <= ackR(1);
      ptr_deref_2183_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1946_word_address_0 & ptr_deref_2183_word_address_0;
      ptr_deref_1946_data_0 <= data_out(15 downto 8);
      ptr_deref_2183_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(6),
          mack => memory_space_3_lr_ack(6),
          maddr => memory_space_3_lr_addr(76 downto 66),
          mtag => memory_space_3_lr_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(6),
          mack => memory_space_3_lc_ack(6),
          mdata => memory_space_3_lc_data(55 downto 48),
          mtag => memory_space_3_lc_tag(13 downto 12),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_2207_load_0 ptr_deref_1965_load_0 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2207_load_0_req_0;
      reqL(0) <= ptr_deref_1965_load_0_req_0;
      ptr_deref_2207_load_0_ack_0 <= ackL(1);
      ptr_deref_1965_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2207_load_0_req_1;
      reqR(0) <= ptr_deref_1965_load_0_req_1;
      ptr_deref_2207_load_0_ack_1 <= ackR(1);
      ptr_deref_1965_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2207_word_address_0 & ptr_deref_1965_word_address_0;
      ptr_deref_2207_data_0 <= data_out(15 downto 8);
      ptr_deref_1965_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(5),
          mack => memory_space_3_lr_ack(5),
          maddr => memory_space_3_lr_addr(65 downto 55),
          mtag => memory_space_3_lr_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(5),
          mack => memory_space_3_lc_ack(5),
          mdata => memory_space_3_lc_data(47 downto 40),
          mtag => memory_space_3_lc_tag(11 downto 10),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_1984_load_0 ptr_deref_2231_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_1984_load_0_req_0;
      reqL(0) <= ptr_deref_2231_load_0_req_0;
      ptr_deref_1984_load_0_ack_0 <= ackL(1);
      ptr_deref_2231_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_1984_load_0_req_1;
      reqR(0) <= ptr_deref_2231_load_0_req_1;
      ptr_deref_1984_load_0_ack_1 <= ackR(1);
      ptr_deref_2231_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1984_word_address_0 & ptr_deref_2231_word_address_0;
      ptr_deref_1984_data_0 <= data_out(15 downto 8);
      ptr_deref_2231_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(4),
          mack => memory_space_3_lr_ack(4),
          maddr => memory_space_3_lr_addr(54 downto 44),
          mtag => memory_space_3_lr_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(4),
          mack => memory_space_3_lc_ack(4),
          mdata => memory_space_3_lc_data(39 downto 32),
          mtag => memory_space_3_lc_tag(9 downto 8),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : ptr_deref_2003_load_0 ptr_deref_2255_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2003_load_0_req_0;
      reqL(0) <= ptr_deref_2255_load_0_req_0;
      ptr_deref_2003_load_0_ack_0 <= ackL(1);
      ptr_deref_2255_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2003_load_0_req_1;
      reqR(0) <= ptr_deref_2255_load_0_req_1;
      ptr_deref_2003_load_0_ack_1 <= ackR(1);
      ptr_deref_2255_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2003_word_address_0 & ptr_deref_2255_word_address_0;
      ptr_deref_2003_data_0 <= data_out(15 downto 8);
      ptr_deref_2255_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(3),
          mack => memory_space_3_lr_ack(3),
          maddr => memory_space_3_lr_addr(43 downto 33),
          mtag => memory_space_3_lr_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(3),
          mack => memory_space_3_lc_ack(3),
          mdata => memory_space_3_lc_data(31 downto 24),
          mtag => memory_space_3_lc_tag(7 downto 6),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- shared load operator group (5) : ptr_deref_2022_load_0 ptr_deref_2279_load_0 
    LoadGroup5: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2022_load_0_req_0;
      reqL(0) <= ptr_deref_2279_load_0_req_0;
      ptr_deref_2022_load_0_ack_0 <= ackL(1);
      ptr_deref_2279_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2022_load_0_req_1;
      reqR(0) <= ptr_deref_2279_load_0_req_1;
      ptr_deref_2022_load_0_ack_1 <= ackR(1);
      ptr_deref_2279_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2022_word_address_0 & ptr_deref_2279_word_address_0;
      ptr_deref_2022_data_0 <= data_out(15 downto 8);
      ptr_deref_2279_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(2),
          mack => memory_space_3_lr_ack(2),
          maddr => memory_space_3_lr_addr(32 downto 22),
          mtag => memory_space_3_lr_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(2),
          mack => memory_space_3_lc_ack(2),
          mdata => memory_space_3_lc_data(23 downto 16),
          mtag => memory_space_3_lc_tag(5 downto 4),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 5
    -- shared load operator group (6) : ptr_deref_2036_load_0 ptr_deref_2303_load_0 
    LoadGroup6: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2036_load_0_req_0;
      reqL(0) <= ptr_deref_2303_load_0_req_0;
      ptr_deref_2036_load_0_ack_0 <= ackL(1);
      ptr_deref_2303_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2036_load_0_req_1;
      reqR(0) <= ptr_deref_2303_load_0_req_1;
      ptr_deref_2036_load_0_ack_1 <= ackR(1);
      ptr_deref_2303_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2036_word_address_0 & ptr_deref_2303_word_address_0;
      ptr_deref_2036_data_0 <= data_out(15 downto 8);
      ptr_deref_2303_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(1),
          mack => memory_space_3_lr_ack(1),
          maddr => memory_space_3_lr_addr(21 downto 11),
          mtag => memory_space_3_lr_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(1),
          mack => memory_space_3_lc_ack(1),
          mdata => memory_space_3_lc_data(15 downto 8),
          mtag => memory_space_3_lc_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 6
    -- shared load operator group (7) : ptr_deref_2055_load_0 ptr_deref_2321_load_0 
    LoadGroup7: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_2055_load_0_req_0;
      reqL(0) <= ptr_deref_2321_load_0_req_0;
      ptr_deref_2055_load_0_ack_0 <= ackL(1);
      ptr_deref_2321_load_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2055_load_0_req_1;
      reqR(0) <= ptr_deref_2321_load_0_req_1;
      ptr_deref_2055_load_0_ack_1 <= ackR(1);
      ptr_deref_2321_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2055_word_address_0 & ptr_deref_2321_word_address_0;
      ptr_deref_2055_data_0 <= data_out(15 downto 8);
      ptr_deref_2321_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 11,  num_reqs => 2,  tag_length => 2, min_clock_period => false,
        no_arbitration => true)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(10 downto 0),
          mtag => memory_space_3_lr_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 2,  no_arbitration => true)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 7
    -- shared inport operator group (0) : simple_obj_ref_1902_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1902_inst_req_0;
      simple_obj_ref_1902_inst_ack_0 <= ack(0);
      tmp_1903 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => midpipe_pipe_read_req(0),
          oack => midpipe_pipe_read_ack(0),
          odata => midpipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_1915_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1915_inst_req_0;
      simple_obj_ref_1915_inst_ack_0 <= ack(0);
      tmp125_1916 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => pkt_length_pipe_read_req(0),
          oack => pkt_length_pipe_read_ack(0),
          odata => pkt_length_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_1924_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1924_inst_req_0;
      simple_obj_ref_1924_inst_ack_0 <= ack(0);
      tmp126_1925 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => last_ctrl_pipe_read_req(0),
          oack => last_ctrl_pipe_read_ack(0),
          odata => last_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : simple_obj_ref_2108_inst simple_obj_ref_2381_inst simple_obj_ref_2402_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_2108_inst_req_0;
      req(1) <= simple_obj_ref_2381_inst_req_0;
      req(0) <= simple_obj_ref_2402_inst_req_0;
      simple_obj_ref_2108_inst_ack_0 <= ack(2);
      simple_obj_ref_2381_inst_ack_0 <= ack(1);
      simple_obj_ref_2402_inst_ack_0 <= ack(0);
      data_in <= type_cast_2110_wire_constant & type_cast_2383_wire_constant & tmp126_1925;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => op_lut_ctrl_pipe_write_req(0),
          oack => op_lut_ctrl_pipe_write_ack(0),
          odata => op_lut_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : simple_obj_ref_2118_inst simple_obj_ref_2391_inst simple_obj_ref_2411_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_2118_inst_req_0;
      req(1) <= simple_obj_ref_2391_inst_req_0;
      req(0) <= simple_obj_ref_2411_inst_req_0;
      simple_obj_ref_2118_inst_ack_0 <= ack(2);
      simple_obj_ref_2391_inst_ack_0 <= ack(1);
      simple_obj_ref_2411_inst_ack_0 <= ack(0);
      data_in <= ins38_2101 & ins77_2367 & ins77_2367;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 3,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => op_lut_data_pipe_write_req(0),
          oack => op_lut_data_pipe_write_ack(0),
          odata => op_lut_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : simple_obj_ref_2420_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2420_inst_req_0;
      simple_obj_ref_2420_inst_ack_0 <= ack(0);
      data_in <= type_cast_2422_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_request_pipe_write_req(0),
          oack => free_queue_request_pipe_write_ack(0),
          odata => free_queue_request_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : simple_obj_ref_2430_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2430_inst_req_0;
      simple_obj_ref_2430_inst_ack_0 <= ack(0);
      data_in <= tmp_1903;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => true)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_put_pipe_write_req(0),
          oack => free_queue_put_pipe_write_ack(0),
          odata => free_queue_put_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
    in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
    in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
    out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(3 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_10
  -- interface signals to connect to memory space memory_space_11
  -- interface signals to connect to memory space memory_space_12
  -- interface signals to connect to memory space memory_space_13
  -- interface signals to connect to memory space memory_space_14
  -- interface signals to connect to memory space memory_space_15
  -- interface signals to connect to memory space memory_space_16
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(2 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(3 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(11 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(3 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(3 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(7 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(7 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(7 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(87 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(15 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(15 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(7 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(87 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(15 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(7 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(15 downto 0);
  -- interface signals to connect to memory space memory_space_4
  -- interface signals to connect to memory space memory_space_5
  -- interface signals to connect to memory space memory_space_6
  -- interface signals to connect to memory space memory_space_7
  -- interface signals to connect to memory space memory_space_8
  -- interface signals to connect to memory space memory_space_9
  -- declarations related to module free_queue_manager
  component free_queue_manager is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(2 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(1 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(1 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(11 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(3 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(3 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(7 downto 0);
      free_queue_request_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_put_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_get_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_manager
  signal free_queue_manager_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal free_queue_manager_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_manager_start_req : std_logic;
  signal free_queue_manager_start_ack : std_logic;
  signal free_queue_manager_fin_req   : std_logic;
  signal free_queue_manager_fin_ack : std_logic;
  -- declarations related to module output_port_lookup
  component output_port_lookup is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      op_lut_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      op_lut_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      op_lut_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      op_lut_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module output_port_lookup
  signal output_port_lookup_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal output_port_lookup_tag_out   : std_logic_vector(0 downto 0);
  signal output_port_lookup_start_req : std_logic;
  signal output_port_lookup_start_ack : std_logic;
  signal output_port_lookup_fin_req   : std_logic;
  signal output_port_lookup_fin_ack : std_logic;
  -- declarations related to module wrapper_input
  component wrapper_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_3_sr_req : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(87 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(63 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(7 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(15 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(3 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(0 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_ack_pipe_read_data : in   std_logic_vector(7 downto 0);
      free_queue_get_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_get_pipe_read_data : in   std_logic_vector(31 downto 0);
      in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      midpipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      last_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      last_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      last_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      pkt_length_pipe_write_req : out  std_logic_vector(0 downto 0);
      pkt_length_pipe_write_ack : in   std_logic_vector(0 downto 0);
      pkt_length_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_input
  signal wrapper_input_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_input_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic;
  signal wrapper_input_start_ack : std_logic;
  signal wrapper_input_fin_req   : std_logic;
  signal wrapper_input_fin_ack : std_logic;
  -- declarations related to module wrapper_output
  component wrapper_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_3_lr_req : out  std_logic_vector(7 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(87 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(15 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(7 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(7 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(63 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(15 downto 0);
      midpipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      midpipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      midpipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      last_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      last_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      last_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      pkt_length_pipe_read_req : out  std_logic_vector(0 downto 0);
      pkt_length_pipe_read_ack : in   std_logic_vector(0 downto 0);
      pkt_length_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_request_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_request_pipe_write_data : out  std_logic_vector(7 downto 0);
      free_queue_put_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_put_pipe_write_data : out  std_logic_vector(31 downto 0);
      op_lut_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      op_lut_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      op_lut_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      op_lut_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      op_lut_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_output
  signal wrapper_output_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_output_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic;
  signal wrapper_output_start_ack : std_logic;
  signal wrapper_output_fin_req   : std_logic;
  signal wrapper_output_fin_ack : std_logic;
  -- aggregate signals for write to pipe free_queue_ack
  signal free_queue_ack_pipe_write_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_ack
  signal free_queue_ack_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_ack_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_ack_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_get
  signal free_queue_get_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_get
  signal free_queue_get_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_get_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_get_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_put
  signal free_queue_put_pipe_write_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_write_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe free_queue_put
  signal free_queue_put_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_put_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_put_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe free_queue_request
  signal free_queue_request_pipe_write_data: std_logic_vector(15 downto 0);
  signal free_queue_request_pipe_write_req: std_logic_vector(1 downto 0);
  signal free_queue_request_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe free_queue_request
  signal free_queue_request_pipe_read_data: std_logic_vector(7 downto 0);
  signal free_queue_request_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_request_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_ctrl
  signal in_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe last_ctrl
  signal last_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal last_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal last_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe last_ctrl
  signal last_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal last_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal last_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe midpipe
  signal midpipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe midpipe
  signal midpipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal midpipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal midpipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe op_lut_ctrl
  signal op_lut_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal op_lut_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal op_lut_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe op_lut_ctrl
  signal op_lut_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal op_lut_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal op_lut_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe op_lut_data
  signal op_lut_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal op_lut_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal op_lut_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe op_lut_data
  signal op_lut_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal op_lut_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal op_lut_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_ctrl
  signal out_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe pkt_length
  signal pkt_length_pipe_write_data: std_logic_vector(31 downto 0);
  signal pkt_length_pipe_write_req: std_logic_vector(0 downto 0);
  signal pkt_length_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe pkt_length
  signal pkt_length_pipe_read_data: std_logic_vector(31 downto 0);
  signal pkt_length_pipe_read_req: std_logic_vector(0 downto 0);
  signal pkt_length_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module free_queue_manager
  free_queue_manager_instance:free_queue_manager-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => free_queue_manager_start_req,
      start_ack => free_queue_manager_start_ack,
      fin_req => free_queue_manager_fin_req,
      fin_ack => free_queue_manager_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(2 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(1 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(7 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(1 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(3 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(3 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(11 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(7 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(3 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(3 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(7 downto 0),
      free_queue_request_pipe_read_req => free_queue_request_pipe_read_req(0 downto 0),
      free_queue_request_pipe_read_ack => free_queue_request_pipe_read_ack(0 downto 0),
      free_queue_request_pipe_read_data => free_queue_request_pipe_read_data(7 downto 0),
      free_queue_put_pipe_read_req => free_queue_put_pipe_read_req(0 downto 0),
      free_queue_put_pipe_read_ack => free_queue_put_pipe_read_ack(0 downto 0),
      free_queue_put_pipe_read_data => free_queue_put_pipe_read_data(31 downto 0),
      free_queue_ack_pipe_write_req => free_queue_ack_pipe_write_req(0 downto 0),
      free_queue_ack_pipe_write_ack => free_queue_ack_pipe_write_ack(0 downto 0),
      free_queue_ack_pipe_write_data => free_queue_ack_pipe_write_data(7 downto 0),
      free_queue_get_pipe_write_req => free_queue_get_pipe_write_req(0 downto 0),
      free_queue_get_pipe_write_ack => free_queue_get_pipe_write_ack(0 downto 0),
      free_queue_get_pipe_write_data => free_queue_get_pipe_write_data(31 downto 0),
      tag_in => free_queue_manager_tag_in,
      tag_out => free_queue_manager_tag_out-- 
    ); -- 
  -- module will be run forever 
  free_queue_manager_tag_in <= (others => '0');
  free_queue_manager_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => free_queue_manager_start_req, start_ack => free_queue_manager_start_ack,  fin_req => free_queue_manager_fin_req,  fin_ack => free_queue_manager_fin_ack);
  -- module output_port_lookup
  output_port_lookup_instance:output_port_lookup-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => output_port_lookup_start_req,
      start_ack => output_port_lookup_start_ack,
      fin_req => output_port_lookup_fin_req,
      fin_ack => output_port_lookup_fin_ack,
      clk => clk,
      reset => reset,
      op_lut_ctrl_pipe_read_req => op_lut_ctrl_pipe_read_req(0 downto 0),
      op_lut_ctrl_pipe_read_ack => op_lut_ctrl_pipe_read_ack(0 downto 0),
      op_lut_ctrl_pipe_read_data => op_lut_ctrl_pipe_read_data(7 downto 0),
      op_lut_data_pipe_read_req => op_lut_data_pipe_read_req(0 downto 0),
      op_lut_data_pipe_read_ack => op_lut_data_pipe_read_ack(0 downto 0),
      op_lut_data_pipe_read_data => op_lut_data_pipe_read_data(63 downto 0),
      out_ctrl_pipe_write_req => out_ctrl_pipe_write_req(0 downto 0),
      out_ctrl_pipe_write_ack => out_ctrl_pipe_write_ack(0 downto 0),
      out_ctrl_pipe_write_data => out_ctrl_pipe_write_data(7 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      tag_in => output_port_lookup_tag_in,
      tag_out => output_port_lookup_tag_out-- 
    ); -- 
  -- module will be run forever 
  output_port_lookup_tag_in <= (others => '0');
  output_port_lookup_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => output_port_lookup_start_req, start_ack => output_port_lookup_start_ack,  fin_req => output_port_lookup_fin_req,  fin_ack => output_port_lookup_fin_ack);
  -- module wrapper_input
  wrapper_input_instance:wrapper_input-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_input_start_req,
      start_ack => wrapper_input_start_ack,
      fin_req => wrapper_input_fin_req,
      fin_ack => wrapper_input_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(3 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(0 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(0 downto 0),
      memory_space_3_sr_req => memory_space_3_sr_req(7 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(7 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(87 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(63 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(15 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(7 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(7 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(15 downto 0),
      free_queue_ack_pipe_read_req => free_queue_ack_pipe_read_req(0 downto 0),
      free_queue_ack_pipe_read_ack => free_queue_ack_pipe_read_ack(0 downto 0),
      free_queue_ack_pipe_read_data => free_queue_ack_pipe_read_data(7 downto 0),
      free_queue_get_pipe_read_req => free_queue_get_pipe_read_req(0 downto 0),
      free_queue_get_pipe_read_ack => free_queue_get_pipe_read_ack(0 downto 0),
      free_queue_get_pipe_read_data => free_queue_get_pipe_read_data(31 downto 0),
      in_ctrl_pipe_read_req => in_ctrl_pipe_read_req(0 downto 0),
      in_ctrl_pipe_read_ack => in_ctrl_pipe_read_ack(0 downto 0),
      in_ctrl_pipe_read_data => in_ctrl_pipe_read_data(7 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(1 downto 1),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(1 downto 1),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(15 downto 8),
      midpipe_pipe_write_req => midpipe_pipe_write_req(0 downto 0),
      midpipe_pipe_write_ack => midpipe_pipe_write_ack(0 downto 0),
      midpipe_pipe_write_data => midpipe_pipe_write_data(31 downto 0),
      last_ctrl_pipe_write_req => last_ctrl_pipe_write_req(0 downto 0),
      last_ctrl_pipe_write_ack => last_ctrl_pipe_write_ack(0 downto 0),
      last_ctrl_pipe_write_data => last_ctrl_pipe_write_data(7 downto 0),
      pkt_length_pipe_write_req => pkt_length_pipe_write_req(0 downto 0),
      pkt_length_pipe_write_ack => pkt_length_pipe_write_ack(0 downto 0),
      pkt_length_pipe_write_data => pkt_length_pipe_write_data(31 downto 0),
      tag_in => wrapper_input_tag_in,
      tag_out => wrapper_input_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_input_tag_in <= (others => '0');
  wrapper_input_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_input_start_req, start_ack => wrapper_input_start_ack,  fin_req => wrapper_input_fin_req,  fin_ack => wrapper_input_fin_ack);
  -- module wrapper_output
  wrapper_output_instance:wrapper_output-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_output_start_req,
      start_ack => wrapper_output_start_ack,
      fin_req => wrapper_output_fin_req,
      fin_ack => wrapper_output_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_3_lr_req => memory_space_3_lr_req(7 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(7 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(87 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(15 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(7 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(7 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(63 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(15 downto 0),
      midpipe_pipe_read_req => midpipe_pipe_read_req(0 downto 0),
      midpipe_pipe_read_ack => midpipe_pipe_read_ack(0 downto 0),
      midpipe_pipe_read_data => midpipe_pipe_read_data(31 downto 0),
      last_ctrl_pipe_read_req => last_ctrl_pipe_read_req(0 downto 0),
      last_ctrl_pipe_read_ack => last_ctrl_pipe_read_ack(0 downto 0),
      last_ctrl_pipe_read_data => last_ctrl_pipe_read_data(7 downto 0),
      pkt_length_pipe_read_req => pkt_length_pipe_read_req(0 downto 0),
      pkt_length_pipe_read_ack => pkt_length_pipe_read_ack(0 downto 0),
      pkt_length_pipe_read_data => pkt_length_pipe_read_data(31 downto 0),
      free_queue_request_pipe_write_req => free_queue_request_pipe_write_req(0 downto 0),
      free_queue_request_pipe_write_ack => free_queue_request_pipe_write_ack(0 downto 0),
      free_queue_request_pipe_write_data => free_queue_request_pipe_write_data(7 downto 0),
      free_queue_put_pipe_write_req => free_queue_put_pipe_write_req(0 downto 0),
      free_queue_put_pipe_write_ack => free_queue_put_pipe_write_ack(0 downto 0),
      free_queue_put_pipe_write_data => free_queue_put_pipe_write_data(31 downto 0),
      op_lut_ctrl_pipe_write_req => op_lut_ctrl_pipe_write_req(0 downto 0),
      op_lut_ctrl_pipe_write_ack => op_lut_ctrl_pipe_write_ack(0 downto 0),
      op_lut_ctrl_pipe_write_data => op_lut_ctrl_pipe_write_data(7 downto 0),
      op_lut_data_pipe_write_req => op_lut_data_pipe_write_req(0 downto 0),
      op_lut_data_pipe_write_ack => op_lut_data_pipe_write_ack(0 downto 0),
      op_lut_data_pipe_write_data => op_lut_data_pipe_write_data(63 downto 0),
      tag_in => wrapper_output_tag_in,
      tag_out => wrapper_output_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_output_tag_in <= (others => '0');
  wrapper_output_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_output_start_req, start_ack => wrapper_output_start_ack,  fin_req => wrapper_output_fin_req,  fin_ack => wrapper_output_fin_ack);
  free_queue_ack_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_ack_pipe_read_req,
      read_ack => free_queue_ack_pipe_read_ack,
      read_data => free_queue_ack_pipe_read_data,
      write_req => free_queue_ack_pipe_write_req,
      write_ack => free_queue_ack_pipe_write_ack,
      write_data => free_queue_ack_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_get_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_get_pipe_read_req,
      read_ack => free_queue_get_pipe_read_ack,
      read_data => free_queue_get_pipe_read_data,
      write_req => free_queue_get_pipe_write_req,
      write_ack => free_queue_get_pipe_write_ack,
      write_data => free_queue_get_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_put_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_put_pipe_read_req,
      read_ack => free_queue_put_pipe_read_ack,
      read_data => free_queue_put_pipe_read_data,
      write_req => free_queue_put_pipe_write_req,
      write_ack => free_queue_put_pipe_write_ack,
      write_data => free_queue_put_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_request_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => free_queue_request_pipe_read_req,
      read_ack => free_queue_request_pipe_read_ack,
      read_data => free_queue_request_pipe_read_data,
      write_req => free_queue_request_pipe_write_req,
      write_ack => free_queue_request_pipe_write_ack,
      write_data => free_queue_request_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => in_ctrl_pipe_read_req,
      read_ack => in_ctrl_pipe_read_ack,
      read_data => in_ctrl_pipe_read_data,
      write_req => in_ctrl_pipe_write_req,
      write_ack => in_ctrl_pipe_write_ack,
      write_data => in_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  last_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => last_ctrl_pipe_read_req,
      read_ack => last_ctrl_pipe_read_ack,
      read_data => last_ctrl_pipe_read_data,
      write_req => last_ctrl_pipe_write_req,
      write_ack => last_ctrl_pipe_write_ack,
      write_data => last_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  midpipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => midpipe_pipe_read_req,
      read_ack => midpipe_pipe_read_ack,
      read_data => midpipe_pipe_read_data,
      write_req => midpipe_pipe_write_req,
      write_ack => midpipe_pipe_write_ack,
      write_data => midpipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  op_lut_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => op_lut_ctrl_pipe_read_req,
      read_ack => op_lut_ctrl_pipe_read_ack,
      read_data => op_lut_ctrl_pipe_read_data,
      write_req => op_lut_ctrl_pipe_write_req,
      write_ack => op_lut_ctrl_pipe_write_ack,
      write_data => op_lut_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  op_lut_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => op_lut_data_pipe_read_req,
      read_ack => op_lut_data_pipe_read_ack,
      read_data => op_lut_data_pipe_read_data,
      write_req => op_lut_data_pipe_write_req,
      write_ack => op_lut_data_pipe_write_ack,
      write_data => op_lut_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => out_ctrl_pipe_read_req,
      read_ack => out_ctrl_pipe_read_ack,
      read_data => out_ctrl_pipe_read_data,
      write_req => out_ctrl_pipe_write_req,
      write_ack => out_ctrl_pipe_write_ack,
      write_data => out_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  pkt_length_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => pkt_length_pipe_read_req,
      read_ack => pkt_length_pipe_read_ack,
      read_data => pkt_length_pipe_read_data,
      write_req => pkt_length_pipe_write_req,
      write_ack => pkt_length_pipe_write_ack,
      write_data => pkt_length_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  dummyWOM_memory_space_1: dummy_write_only_memory_subsystem -- 
    generic map(-- 
      num_stores => 1,
      addr_width => 4,
      data_width => 8,
      tag_width => 1
      ) -- 
    port map(-- 
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  RegisterBank_memory_space_2: register_bank -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 4,
      addr_width => 3,
      data_width => 8,
      tag_width => 2,
      num_registers => 4) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: memory_subsystem -- 
    generic map(-- 
      num_loads => 8,
      num_stores => 8,
      addr_width => 11,
      data_width => 8,
      tag_width => 2,
      number_of_banks => 4,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
