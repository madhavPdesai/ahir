library work;
use work.cpath_components.all;

entity start_cp is
  port (

    ip    : in bit_vector(275 downto 1);
    op    : out bit_vector(278 downto 1) := (others => '0');
    reset : in bit;
    clk   : in bit);
end start_cp;

architecture behavioral of start_cp is

  signal place_1_tip : bit_vector(0 downto 0);
  signal place_1_rst : bit_vector(0 downto 0);
  signal place_1_top : bit;
  signal place_100_tip : bit_vector(1 downto 0);
  signal place_100_rst : bit_vector(0 downto 0);
  signal place_100_top : bit;
  signal place_101_tip : bit_vector(0 downto 0);
  signal place_101_rst : bit_vector(0 downto 0);
  signal place_101_top : bit;
  signal place_105_tip : bit_vector(1 downto 0);
  signal place_105_rst : bit_vector(0 downto 0);
  signal place_105_top : bit;
  signal place_106_tip : bit_vector(0 downto 0);
  signal place_106_rst : bit_vector(0 downto 0);
  signal place_106_top : bit;
  signal place_107_tip : bit_vector(0 downto 0);
  signal place_107_rst : bit_vector(0 downto 0);
  signal place_107_top : bit;
  signal place_108_tip : bit_vector(0 downto 0);
  signal place_108_rst : bit_vector(0 downto 0);
  signal place_108_top : bit;
  signal place_109_tip : bit_vector(0 downto 0);
  signal place_109_rst : bit_vector(0 downto 0);
  signal place_109_top : bit;
  signal place_110_tip : bit_vector(0 downto 0);
  signal place_110_rst : bit_vector(0 downto 0);
  signal place_110_top : bit;
  signal place_111_tip : bit_vector(0 downto 0);
  signal place_111_rst : bit_vector(0 downto 0);
  signal place_111_top : bit;
  signal place_112_tip : bit_vector(0 downto 0);
  signal place_112_rst : bit_vector(0 downto 0);
  signal place_112_top : bit;
  signal place_113_tip : bit_vector(0 downto 0);
  signal place_113_rst : bit_vector(0 downto 0);
  signal place_113_top : bit;
  signal place_114_tip : bit_vector(0 downto 0);
  signal place_114_rst : bit_vector(0 downto 0);
  signal place_114_top : bit;
  signal place_115_tip : bit_vector(0 downto 0);
  signal place_115_rst : bit_vector(0 downto 0);
  signal place_115_top : bit;
  signal place_116_tip : bit_vector(0 downto 0);
  signal place_116_rst : bit_vector(0 downto 0);
  signal place_116_top : bit;
  signal place_117_tip : bit_vector(0 downto 0);
  signal place_117_rst : bit_vector(0 downto 0);
  signal place_117_top : bit;
  signal place_118_tip : bit_vector(0 downto 0);
  signal place_118_rst : bit_vector(0 downto 0);
  signal place_118_top : bit;
  signal place_119_tip : bit_vector(0 downto 0);
  signal place_119_rst : bit_vector(0 downto 0);
  signal place_119_top : bit;
  signal place_120_tip : bit_vector(0 downto 0);
  signal place_120_rst : bit_vector(0 downto 0);
  signal place_120_top : bit;
  signal place_121_tip : bit_vector(0 downto 0);
  signal place_121_rst : bit_vector(0 downto 0);
  signal place_121_top : bit;
  signal place_122_tip : bit_vector(0 downto 0);
  signal place_122_rst : bit_vector(1 downto 0);
  signal place_122_top : bit;
  signal place_123_tip : bit_vector(0 downto 0);
  signal place_123_rst : bit_vector(0 downto 0);
  signal place_123_top : bit;
  signal place_124_tip : bit_vector(0 downto 0);
  signal place_124_rst : bit_vector(0 downto 0);
  signal place_124_top : bit;
  signal place_126_tip : bit_vector(0 downto 0);
  signal place_126_rst : bit_vector(0 downto 0);
  signal place_126_top : bit;
  signal place_127_tip : bit_vector(0 downto 0);
  signal place_127_rst : bit_vector(0 downto 0);
  signal place_127_top : bit;
  signal place_128_tip : bit_vector(0 downto 0);
  signal place_128_rst : bit_vector(0 downto 0);
  signal place_128_top : bit;
  signal place_129_tip : bit_vector(0 downto 0);
  signal place_129_rst : bit_vector(1 downto 0);
  signal place_129_top : bit;
  signal place_130_tip : bit_vector(0 downto 0);
  signal place_130_rst : bit_vector(0 downto 0);
  signal place_130_top : bit;
  signal place_132_tip : bit_vector(0 downto 0);
  signal place_132_rst : bit_vector(0 downto 0);
  signal place_132_top : bit;
  signal place_133_tip : bit_vector(0 downto 0);
  signal place_133_rst : bit_vector(1 downto 0);
  signal place_133_top : bit;
  signal place_136_tip : bit_vector(1 downto 0);
  signal place_136_rst : bit_vector(0 downto 0);
  signal place_136_top : bit;
  signal place_137_tip : bit_vector(0 downto 0);
  signal place_137_rst : bit_vector(0 downto 0);
  signal place_137_top : bit;
  signal place_138_tip : bit_vector(0 downto 0);
  signal place_138_rst : bit_vector(0 downto 0);
  signal place_138_top : bit;
  signal place_139_tip : bit_vector(0 downto 0);
  signal place_139_rst : bit_vector(0 downto 0);
  signal place_139_top : bit;
  signal place_14_tip : bit_vector(1 downto 0);
  signal place_14_rst : bit_vector(0 downto 0);
  signal place_14_top : bit;
  signal place_140_tip : bit_vector(0 downto 0);
  signal place_140_rst : bit_vector(0 downto 0);
  signal place_140_top : bit;
  signal place_141_tip : bit_vector(0 downto 0);
  signal place_141_rst : bit_vector(0 downto 0);
  signal place_141_top : bit;
  signal place_142_tip : bit_vector(0 downto 0);
  signal place_142_rst : bit_vector(0 downto 0);
  signal place_142_top : bit;
  signal place_143_tip : bit_vector(0 downto 0);
  signal place_143_rst : bit_vector(0 downto 0);
  signal place_143_top : bit;
  signal place_144_tip : bit_vector(0 downto 0);
  signal place_144_rst : bit_vector(0 downto 0);
  signal place_144_top : bit;
  signal place_145_tip : bit_vector(0 downto 0);
  signal place_145_rst : bit_vector(0 downto 0);
  signal place_145_top : bit;
  signal place_146_tip : bit_vector(0 downto 0);
  signal place_146_rst : bit_vector(0 downto 0);
  signal place_146_top : bit;
  signal place_147_tip : bit_vector(0 downto 0);
  signal place_147_rst : bit_vector(0 downto 0);
  signal place_147_top : bit;
  signal place_148_tip : bit_vector(0 downto 0);
  signal place_148_rst : bit_vector(0 downto 0);
  signal place_148_top : bit;
  signal place_149_tip : bit_vector(0 downto 0);
  signal place_149_rst : bit_vector(0 downto 0);
  signal place_149_top : bit;
  signal place_150_tip : bit_vector(0 downto 0);
  signal place_150_rst : bit_vector(0 downto 0);
  signal place_150_top : bit;
  signal place_151_tip : bit_vector(0 downto 0);
  signal place_151_rst : bit_vector(0 downto 0);
  signal place_151_top : bit;
  signal place_152_tip : bit_vector(0 downto 0);
  signal place_152_rst : bit_vector(0 downto 0);
  signal place_152_top : bit;
  signal place_153_tip : bit_vector(0 downto 0);
  signal place_153_rst : bit_vector(0 downto 0);
  signal place_153_top : bit;
  signal place_154_tip : bit_vector(0 downto 0);
  signal place_154_rst : bit_vector(0 downto 0);
  signal place_154_top : bit;
  signal place_155_tip : bit_vector(0 downto 0);
  signal place_155_rst : bit_vector(0 downto 0);
  signal place_155_top : bit;
  signal place_156_tip : bit_vector(0 downto 0);
  signal place_156_rst : bit_vector(0 downto 0);
  signal place_156_top : bit;
  signal place_157_tip : bit_vector(0 downto 0);
  signal place_157_rst : bit_vector(0 downto 0);
  signal place_157_top : bit;
  signal place_158_tip : bit_vector(0 downto 0);
  signal place_158_rst : bit_vector(0 downto 0);
  signal place_158_top : bit;
  signal place_159_tip : bit_vector(0 downto 0);
  signal place_159_rst : bit_vector(0 downto 0);
  signal place_159_top : bit;
  signal place_16_tip : bit_vector(0 downto 0);
  signal place_16_rst : bit_vector(0 downto 0);
  signal place_16_top : bit;
  signal place_160_tip : bit_vector(0 downto 0);
  signal place_160_rst : bit_vector(0 downto 0);
  signal place_160_top : bit;
  signal place_161_tip : bit_vector(0 downto 0);
  signal place_161_rst : bit_vector(0 downto 0);
  signal place_161_top : bit;
  signal place_162_tip : bit_vector(0 downto 0);
  signal place_162_rst : bit_vector(0 downto 0);
  signal place_162_top : bit;
  signal place_163_tip : bit_vector(0 downto 0);
  signal place_163_rst : bit_vector(0 downto 0);
  signal place_163_top : bit;
  signal place_164_tip : bit_vector(0 downto 0);
  signal place_164_rst : bit_vector(0 downto 0);
  signal place_164_top : bit;
  signal place_165_tip : bit_vector(0 downto 0);
  signal place_165_rst : bit_vector(0 downto 0);
  signal place_165_top : bit;
  signal place_166_tip : bit_vector(0 downto 0);
  signal place_166_rst : bit_vector(0 downto 0);
  signal place_166_top : bit;
  signal place_167_tip : bit_vector(0 downto 0);
  signal place_167_rst : bit_vector(0 downto 0);
  signal place_167_top : bit;
  signal place_168_tip : bit_vector(0 downto 0);
  signal place_168_rst : bit_vector(0 downto 0);
  signal place_168_top : bit;
  signal place_169_tip : bit_vector(0 downto 0);
  signal place_169_rst : bit_vector(0 downto 0);
  signal place_169_top : bit;
  signal place_17_tip : bit_vector(0 downto 0);
  signal place_17_rst : bit_vector(0 downto 0);
  signal place_17_top : bit;
  signal place_170_tip : bit_vector(0 downto 0);
  signal place_170_rst : bit_vector(0 downto 0);
  signal place_170_top : bit;
  signal place_171_tip : bit_vector(0 downto 0);
  signal place_171_rst : bit_vector(0 downto 0);
  signal place_171_top : bit;
  signal place_172_tip : bit_vector(0 downto 0);
  signal place_172_rst : bit_vector(0 downto 0);
  signal place_172_top : bit;
  signal place_173_tip : bit_vector(0 downto 0);
  signal place_173_rst : bit_vector(0 downto 0);
  signal place_173_top : bit;
  signal place_174_tip : bit_vector(0 downto 0);
  signal place_174_rst : bit_vector(0 downto 0);
  signal place_174_top : bit;
  signal place_175_tip : bit_vector(0 downto 0);
  signal place_175_rst : bit_vector(0 downto 0);
  signal place_175_top : bit;
  signal place_176_tip : bit_vector(0 downto 0);
  signal place_176_rst : bit_vector(0 downto 0);
  signal place_176_top : bit;
  signal place_177_tip : bit_vector(0 downto 0);
  signal place_177_rst : bit_vector(0 downto 0);
  signal place_177_top : bit;
  signal place_178_tip : bit_vector(0 downto 0);
  signal place_178_rst : bit_vector(0 downto 0);
  signal place_178_top : bit;
  signal place_179_tip : bit_vector(0 downto 0);
  signal place_179_rst : bit_vector(1 downto 0);
  signal place_179_top : bit;
  signal place_180_tip : bit_vector(0 downto 0);
  signal place_180_rst : bit_vector(0 downto 0);
  signal place_180_top : bit;
  signal place_183_tip : bit_vector(0 downto 0);
  signal place_183_rst : bit_vector(0 downto 0);
  signal place_183_top : bit;
  signal place_184_tip : bit_vector(1 downto 0);
  signal place_184_rst : bit_vector(0 downto 0);
  signal place_184_top : bit;
  signal place_185_tip : bit_vector(0 downto 0);
  signal place_185_rst : bit_vector(0 downto 0);
  signal place_185_top : bit;
  signal place_186_tip : bit_vector(0 downto 0);
  signal place_186_rst : bit_vector(0 downto 0);
  signal place_186_top : bit;
  signal place_187_tip : bit_vector(0 downto 0);
  signal place_187_rst : bit_vector(0 downto 0);
  signal place_187_top : bit;
  signal place_188_tip : bit_vector(1 downto 0);
  signal place_188_rst : bit_vector(0 downto 0);
  signal place_188_top : bit;
  signal place_189_tip : bit_vector(0 downto 0);
  signal place_189_rst : bit_vector(0 downto 0);
  signal place_189_top : bit;
  signal place_190_tip : bit_vector(0 downto 0);
  signal place_190_rst : bit_vector(0 downto 0);
  signal place_190_top : bit;
  signal place_191_tip : bit_vector(0 downto 0);
  signal place_191_rst : bit_vector(0 downto 0);
  signal place_191_top : bit;
  signal place_192_tip : bit_vector(0 downto 0);
  signal place_192_rst : bit_vector(0 downto 0);
  signal place_192_top : bit;
  signal place_193_tip : bit_vector(1 downto 0);
  signal place_193_rst : bit_vector(0 downto 0);
  signal place_193_top : bit;
  signal place_194_tip : bit_vector(0 downto 0);
  signal place_194_rst : bit_vector(0 downto 0);
  signal place_194_top : bit;
  signal place_195_tip : bit_vector(0 downto 0);
  signal place_195_rst : bit_vector(0 downto 0);
  signal place_195_top : bit;
  signal place_196_tip : bit_vector(0 downto 0);
  signal place_196_rst : bit_vector(0 downto 0);
  signal place_196_top : bit;
  signal place_197_tip : bit_vector(0 downto 0);
  signal place_197_rst : bit_vector(0 downto 0);
  signal place_197_top : bit;
  signal place_198_tip : bit_vector(0 downto 0);
  signal place_198_rst : bit_vector(0 downto 0);
  signal place_198_top : bit;
  signal place_199_tip : bit_vector(0 downto 0);
  signal place_199_rst : bit_vector(0 downto 0);
  signal place_199_top : bit;
  signal place_20_tip : bit_vector(0 downto 0);
  signal place_20_rst : bit_vector(0 downto 0);
  signal place_20_top : bit;
  signal place_200_tip : bit_vector(0 downto 0);
  signal place_200_rst : bit_vector(0 downto 0);
  signal place_200_top : bit;
  signal place_201_tip : bit_vector(0 downto 0);
  signal place_201_rst : bit_vector(0 downto 0);
  signal place_201_top : bit;
  signal place_202_tip : bit_vector(0 downto 0);
  signal place_202_rst : bit_vector(0 downto 0);
  signal place_202_top : bit;
  signal place_203_tip : bit_vector(0 downto 0);
  signal place_203_rst : bit_vector(0 downto 0);
  signal place_203_top : bit;
  signal place_204_tip : bit_vector(0 downto 0);
  signal place_204_rst : bit_vector(0 downto 0);
  signal place_204_top : bit;
  signal place_205_tip : bit_vector(0 downto 0);
  signal place_205_rst : bit_vector(0 downto 0);
  signal place_205_top : bit;
  signal place_206_tip : bit_vector(0 downto 0);
  signal place_206_rst : bit_vector(0 downto 0);
  signal place_206_top : bit;
  signal place_208_tip : bit_vector(0 downto 0);
  signal place_208_rst : bit_vector(0 downto 0);
  signal place_208_top : bit;
  signal place_209_tip : bit_vector(1 downto 0);
  signal place_209_rst : bit_vector(0 downto 0);
  signal place_209_top : bit;
  signal place_210_tip : bit_vector(0 downto 0);
  signal place_210_rst : bit_vector(0 downto 0);
  signal place_210_top : bit;
  signal place_211_tip : bit_vector(0 downto 0);
  signal place_211_rst : bit_vector(0 downto 0);
  signal place_211_top : bit;
  signal place_212_tip : bit_vector(0 downto 0);
  signal place_212_rst : bit_vector(0 downto 0);
  signal place_212_top : bit;
  signal place_213_tip : bit_vector(1 downto 0);
  signal place_213_rst : bit_vector(0 downto 0);
  signal place_213_top : bit;
  signal place_214_tip : bit_vector(0 downto 0);
  signal place_214_rst : bit_vector(0 downto 0);
  signal place_214_top : bit;
  signal place_215_tip : bit_vector(0 downto 0);
  signal place_215_rst : bit_vector(0 downto 0);
  signal place_215_top : bit;
  signal place_216_tip : bit_vector(0 downto 0);
  signal place_216_rst : bit_vector(0 downto 0);
  signal place_216_top : bit;
  signal place_217_tip : bit_vector(0 downto 0);
  signal place_217_rst : bit_vector(0 downto 0);
  signal place_217_top : bit;
  signal place_218_tip : bit_vector(0 downto 0);
  signal place_218_rst : bit_vector(0 downto 0);
  signal place_218_top : bit;
  signal place_219_tip : bit_vector(0 downto 0);
  signal place_219_rst : bit_vector(0 downto 0);
  signal place_219_top : bit;
  signal place_22_tip : bit_vector(0 downto 0);
  signal place_22_rst : bit_vector(0 downto 0);
  signal place_22_top : bit;
  signal place_220_tip : bit_vector(0 downto 0);
  signal place_220_rst : bit_vector(0 downto 0);
  signal place_220_top : bit;
  signal place_221_tip : bit_vector(0 downto 0);
  signal place_221_rst : bit_vector(0 downto 0);
  signal place_221_top : bit;
  signal place_222_tip : bit_vector(0 downto 0);
  signal place_222_rst : bit_vector(1 downto 0);
  signal place_222_top : bit;
  signal place_223_tip : bit_vector(0 downto 0);
  signal place_223_rst : bit_vector(0 downto 0);
  signal place_223_top : bit;
  signal place_224_tip : bit_vector(0 downto 0);
  signal place_224_rst : bit_vector(0 downto 0);
  signal place_224_top : bit;
  signal place_225_tip : bit_vector(0 downto 0);
  signal place_225_rst : bit_vector(0 downto 0);
  signal place_225_top : bit;
  signal place_226_tip : bit_vector(0 downto 0);
  signal place_226_rst : bit_vector(0 downto 0);
  signal place_226_top : bit;
  signal place_227_tip : bit_vector(0 downto 0);
  signal place_227_rst : bit_vector(0 downto 0);
  signal place_227_top : bit;
  signal place_228_tip : bit_vector(0 downto 0);
  signal place_228_rst : bit_vector(0 downto 0);
  signal place_228_top : bit;
  signal place_229_tip : bit_vector(0 downto 0);
  signal place_229_rst : bit_vector(0 downto 0);
  signal place_229_top : bit;
  signal place_230_tip : bit_vector(0 downto 0);
  signal place_230_rst : bit_vector(0 downto 0);
  signal place_230_top : bit;
  signal place_231_tip : bit_vector(0 downto 0);
  signal place_231_rst : bit_vector(0 downto 0);
  signal place_231_top : bit;
  signal place_232_tip : bit_vector(1 downto 0);
  signal place_232_rst : bit_vector(0 downto 0);
  signal place_232_top : bit;
  signal place_233_tip : bit_vector(0 downto 0);
  signal place_233_rst : bit_vector(0 downto 0);
  signal place_233_top : bit;
  signal place_234_tip : bit_vector(0 downto 0);
  signal place_234_rst : bit_vector(0 downto 0);
  signal place_234_top : bit;
  signal place_235_tip : bit_vector(0 downto 0);
  signal place_235_rst : bit_vector(0 downto 0);
  signal place_235_top : bit;
  signal place_236_tip : bit_vector(1 downto 0);
  signal place_236_rst : bit_vector(0 downto 0);
  signal place_236_top : bit;
  signal place_237_tip : bit_vector(0 downto 0);
  signal place_237_rst : bit_vector(0 downto 0);
  signal place_237_top : bit;
  signal place_238_tip : bit_vector(0 downto 0);
  signal place_238_rst : bit_vector(0 downto 0);
  signal place_238_top : bit;
  signal place_239_tip : bit_vector(0 downto 0);
  signal place_239_rst : bit_vector(0 downto 0);
  signal place_239_top : bit;
  signal place_24_tip : bit_vector(0 downto 0);
  signal place_24_rst : bit_vector(0 downto 0);
  signal place_24_top : bit;
  signal place_240_tip : bit_vector(0 downto 0);
  signal place_240_rst : bit_vector(0 downto 0);
  signal place_240_top : bit;
  signal place_241_tip : bit_vector(0 downto 0);
  signal place_241_rst : bit_vector(0 downto 0);
  signal place_241_top : bit;
  signal place_242_tip : bit_vector(0 downto 0);
  signal place_242_rst : bit_vector(0 downto 0);
  signal place_242_top : bit;
  signal place_243_tip : bit_vector(0 downto 0);
  signal place_243_rst : bit_vector(0 downto 0);
  signal place_243_top : bit;
  signal place_244_tip : bit_vector(0 downto 0);
  signal place_244_rst : bit_vector(0 downto 0);
  signal place_244_top : bit;
  signal place_245_tip : bit_vector(0 downto 0);
  signal place_245_rst : bit_vector(0 downto 0);
  signal place_245_top : bit;
  signal place_246_tip : bit_vector(0 downto 0);
  signal place_246_rst : bit_vector(0 downto 0);
  signal place_246_top : bit;
  signal place_247_tip : bit_vector(0 downto 0);
  signal place_247_rst : bit_vector(0 downto 0);
  signal place_247_top : bit;
  signal place_248_tip : bit_vector(0 downto 0);
  signal place_248_rst : bit_vector(0 downto 0);
  signal place_248_top : bit;
  signal place_249_tip : bit_vector(0 downto 0);
  signal place_249_rst : bit_vector(0 downto 0);
  signal place_249_top : bit;
  signal place_25_tip : bit_vector(0 downto 0);
  signal place_25_rst : bit_vector(0 downto 0);
  signal place_25_top : bit;
  signal place_250_tip : bit_vector(0 downto 0);
  signal place_250_rst : bit_vector(0 downto 0);
  signal place_250_top : bit;
  signal place_251_tip : bit_vector(0 downto 0);
  signal place_251_rst : bit_vector(0 downto 0);
  signal place_251_top : bit;
  signal place_252_tip : bit_vector(0 downto 0);
  signal place_252_rst : bit_vector(0 downto 0);
  signal place_252_top : bit;
  signal place_253_tip : bit_vector(0 downto 0);
  signal place_253_rst : bit_vector(0 downto 0);
  signal place_253_top : bit;
  signal place_254_tip : bit_vector(0 downto 0);
  signal place_254_rst : bit_vector(0 downto 0);
  signal place_254_top : bit;
  signal place_255_tip : bit_vector(0 downto 0);
  signal place_255_rst : bit_vector(0 downto 0);
  signal place_255_top : bit;
  signal place_256_tip : bit_vector(0 downto 0);
  signal place_256_rst : bit_vector(1 downto 0);
  signal place_256_top : bit;
  signal place_257_tip : bit_vector(0 downto 0);
  signal place_257_rst : bit_vector(0 downto 0);
  signal place_257_top : bit;
  signal place_258_tip : bit_vector(0 downto 0);
  signal place_258_rst : bit_vector(0 downto 0);
  signal place_258_top : bit;
  signal place_259_tip : bit_vector(0 downto 0);
  signal place_259_rst : bit_vector(0 downto 0);
  signal place_259_top : bit;
  signal place_260_tip : bit_vector(0 downto 0);
  signal place_260_rst : bit_vector(0 downto 0);
  signal place_260_top : bit;
  signal place_261_tip : bit_vector(0 downto 0);
  signal place_261_rst : bit_vector(0 downto 0);
  signal place_261_top : bit;
  signal place_262_tip : bit_vector(0 downto 0);
  signal place_262_rst : bit_vector(0 downto 0);
  signal place_262_top : bit;
  signal place_263_tip : bit_vector(0 downto 0);
  signal place_263_rst : bit_vector(0 downto 0);
  signal place_263_top : bit;
  signal place_264_tip : bit_vector(0 downto 0);
  signal place_264_rst : bit_vector(0 downto 0);
  signal place_264_top : bit;
  signal place_265_tip : bit_vector(0 downto 0);
  signal place_265_rst : bit_vector(1 downto 0);
  signal place_265_top : bit;
  signal place_268_tip : bit_vector(1 downto 0);
  signal place_268_rst : bit_vector(0 downto 0);
  signal place_268_top : bit;
  signal place_269_tip : bit_vector(0 downto 0);
  signal place_269_rst : bit_vector(0 downto 0);
  signal place_269_top : bit;
  signal place_27_tip : bit_vector(0 downto 0);
  signal place_27_rst : bit_vector(0 downto 0);
  signal place_27_top : bit;
  signal place_270_tip : bit_vector(0 downto 0);
  signal place_270_rst : bit_vector(0 downto 0);
  signal place_270_top : bit;
  signal place_273_tip : bit_vector(1 downto 0);
  signal place_273_rst : bit_vector(0 downto 0);
  signal place_273_top : bit;
  signal place_274_tip : bit_vector(0 downto 0);
  signal place_274_rst : bit_vector(0 downto 0);
  signal place_274_top : bit;
  signal place_275_tip : bit_vector(0 downto 0);
  signal place_275_rst : bit_vector(0 downto 0);
  signal place_275_top : bit;
  signal place_276_tip : bit_vector(0 downto 0);
  signal place_276_rst : bit_vector(0 downto 0);
  signal place_276_top : bit;
  signal place_277_tip : bit_vector(0 downto 0);
  signal place_277_rst : bit_vector(0 downto 0);
  signal place_277_top : bit;
  signal place_278_tip : bit_vector(0 downto 0);
  signal place_278_rst : bit_vector(0 downto 0);
  signal place_278_top : bit;
  signal place_279_tip : bit_vector(0 downto 0);
  signal place_279_rst : bit_vector(0 downto 0);
  signal place_279_top : bit;
  signal place_280_tip : bit_vector(0 downto 0);
  signal place_280_rst : bit_vector(0 downto 0);
  signal place_280_top : bit;
  signal place_281_tip : bit_vector(0 downto 0);
  signal place_281_rst : bit_vector(0 downto 0);
  signal place_281_top : bit;
  signal place_282_tip : bit_vector(0 downto 0);
  signal place_282_rst : bit_vector(0 downto 0);
  signal place_282_top : bit;
  signal place_283_tip : bit_vector(0 downto 0);
  signal place_283_rst : bit_vector(0 downto 0);
  signal place_283_top : bit;
  signal place_284_tip : bit_vector(0 downto 0);
  signal place_284_rst : bit_vector(0 downto 0);
  signal place_284_top : bit;
  signal place_285_tip : bit_vector(0 downto 0);
  signal place_285_rst : bit_vector(0 downto 0);
  signal place_285_top : bit;
  signal place_286_tip : bit_vector(0 downto 0);
  signal place_286_rst : bit_vector(0 downto 0);
  signal place_286_top : bit;
  signal place_287_tip : bit_vector(0 downto 0);
  signal place_287_rst : bit_vector(0 downto 0);
  signal place_287_top : bit;
  signal place_288_tip : bit_vector(0 downto 0);
  signal place_288_rst : bit_vector(0 downto 0);
  signal place_288_top : bit;
  signal place_289_tip : bit_vector(0 downto 0);
  signal place_289_rst : bit_vector(0 downto 0);
  signal place_289_top : bit;
  signal place_290_tip : bit_vector(0 downto 0);
  signal place_290_rst : bit_vector(0 downto 0);
  signal place_290_top : bit;
  signal place_291_tip : bit_vector(0 downto 0);
  signal place_291_rst : bit_vector(0 downto 0);
  signal place_291_top : bit;
  signal place_292_tip : bit_vector(0 downto 0);
  signal place_292_rst : bit_vector(0 downto 0);
  signal place_292_top : bit;
  signal place_293_tip : bit_vector(0 downto 0);
  signal place_293_rst : bit_vector(0 downto 0);
  signal place_293_top : bit;
  signal place_294_tip : bit_vector(0 downto 0);
  signal place_294_rst : bit_vector(0 downto 0);
  signal place_294_top : bit;
  signal place_295_tip : bit_vector(0 downto 0);
  signal place_295_rst : bit_vector(0 downto 0);
  signal place_295_top : bit;
  signal place_296_tip : bit_vector(0 downto 0);
  signal place_296_rst : bit_vector(0 downto 0);
  signal place_296_top : bit;
  signal place_297_tip : bit_vector(0 downto 0);
  signal place_297_rst : bit_vector(0 downto 0);
  signal place_297_top : bit;
  signal place_298_tip : bit_vector(0 downto 0);
  signal place_298_rst : bit_vector(0 downto 0);
  signal place_298_top : bit;
  signal place_299_tip : bit_vector(0 downto 0);
  signal place_299_rst : bit_vector(0 downto 0);
  signal place_299_top : bit;
  signal place_30_tip : bit_vector(0 downto 0);
  signal place_30_rst : bit_vector(0 downto 0);
  signal place_30_top : bit;
  signal place_300_tip : bit_vector(0 downto 0);
  signal place_300_rst : bit_vector(0 downto 0);
  signal place_300_top : bit;
  signal place_301_tip : bit_vector(0 downto 0);
  signal place_301_rst : bit_vector(0 downto 0);
  signal place_301_top : bit;
  signal place_302_tip : bit_vector(0 downto 0);
  signal place_302_rst : bit_vector(0 downto 0);
  signal place_302_top : bit;
  signal place_303_tip : bit_vector(0 downto 0);
  signal place_303_rst : bit_vector(0 downto 0);
  signal place_303_top : bit;
  signal place_304_tip : bit_vector(0 downto 0);
  signal place_304_rst : bit_vector(0 downto 0);
  signal place_304_top : bit;
  signal place_305_tip : bit_vector(0 downto 0);
  signal place_305_rst : bit_vector(0 downto 0);
  signal place_305_top : bit;
  signal place_306_tip : bit_vector(0 downto 0);
  signal place_306_rst : bit_vector(0 downto 0);
  signal place_306_top : bit;
  signal place_307_tip : bit_vector(0 downto 0);
  signal place_307_rst : bit_vector(0 downto 0);
  signal place_307_top : bit;
  signal place_308_tip : bit_vector(0 downto 0);
  signal place_308_rst : bit_vector(0 downto 0);
  signal place_308_top : bit;
  signal place_309_tip : bit_vector(0 downto 0);
  signal place_309_rst : bit_vector(0 downto 0);
  signal place_309_top : bit;
  signal place_310_tip : bit_vector(0 downto 0);
  signal place_310_rst : bit_vector(1 downto 0);
  signal place_310_top : bit;
  signal place_311_tip : bit_vector(0 downto 0);
  signal place_311_rst : bit_vector(0 downto 0);
  signal place_311_top : bit;
  signal place_312_tip : bit_vector(0 downto 0);
  signal place_312_rst : bit_vector(0 downto 0);
  signal place_312_top : bit;
  signal place_313_tip : bit_vector(0 downto 0);
  signal place_313_rst : bit_vector(0 downto 0);
  signal place_313_top : bit;
  signal place_314_tip : bit_vector(0 downto 0);
  signal place_314_rst : bit_vector(0 downto 0);
  signal place_314_top : bit;
  signal place_315_tip : bit_vector(0 downto 0);
  signal place_315_rst : bit_vector(0 downto 0);
  signal place_315_top : bit;
  signal place_316_tip : bit_vector(0 downto 0);
  signal place_316_rst : bit_vector(0 downto 0);
  signal place_316_top : bit;
  signal place_317_tip : bit_vector(0 downto 0);
  signal place_317_rst : bit_vector(0 downto 0);
  signal place_317_top : bit;
  signal place_318_tip : bit_vector(0 downto 0);
  signal place_318_rst : bit_vector(0 downto 0);
  signal place_318_top : bit;
  signal place_319_tip : bit_vector(0 downto 0);
  signal place_319_rst : bit_vector(0 downto 0);
  signal place_319_top : bit;
  signal place_32_tip : bit_vector(0 downto 0);
  signal place_32_rst : bit_vector(0 downto 0);
  signal place_32_top : bit;
  signal place_320_tip : bit_vector(0 downto 0);
  signal place_320_rst : bit_vector(1 downto 0);
  signal place_320_top : bit;
  signal place_322_tip : bit_vector(0 downto 0);
  signal place_322_rst : bit_vector(0 downto 0);
  signal place_322_top : bit;
  signal place_323_tip : bit_vector(1 downto 0);
  signal place_323_rst : bit_vector(0 downto 0);
  signal place_323_top : bit;
  signal place_324_tip : bit_vector(0 downto 0);
  signal place_324_rst : bit_vector(0 downto 0);
  signal place_324_top : bit;
  signal place_325_tip : bit_vector(0 downto 0);
  signal place_325_rst : bit_vector(0 downto 0);
  signal place_325_top : bit;
  signal place_326_tip : bit_vector(0 downto 0);
  signal place_326_rst : bit_vector(0 downto 0);
  signal place_326_top : bit;
  signal place_327_tip : bit_vector(1 downto 0);
  signal place_327_rst : bit_vector(0 downto 0);
  signal place_327_top : bit;
  signal place_328_tip : bit_vector(0 downto 0);
  signal place_328_rst : bit_vector(0 downto 0);
  signal place_328_top : bit;
  signal place_329_tip : bit_vector(0 downto 0);
  signal place_329_rst : bit_vector(0 downto 0);
  signal place_329_top : bit;
  signal place_33_tip : bit_vector(0 downto 0);
  signal place_33_rst : bit_vector(0 downto 0);
  signal place_33_top : bit;
  signal place_330_tip : bit_vector(0 downto 0);
  signal place_330_rst : bit_vector(0 downto 0);
  signal place_330_top : bit;
  signal place_331_tip : bit_vector(0 downto 0);
  signal place_331_rst : bit_vector(0 downto 0);
  signal place_331_top : bit;
  signal place_332_tip : bit_vector(0 downto 0);
  signal place_332_rst : bit_vector(0 downto 0);
  signal place_332_top : bit;
  signal place_333_tip : bit_vector(0 downto 0);
  signal place_333_rst : bit_vector(0 downto 0);
  signal place_333_top : bit;
  signal place_334_tip : bit_vector(0 downto 0);
  signal place_334_rst : bit_vector(0 downto 0);
  signal place_334_top : bit;
  signal place_335_tip : bit_vector(0 downto 0);
  signal place_335_rst : bit_vector(0 downto 0);
  signal place_335_top : bit;
  signal place_336_tip : bit_vector(0 downto 0);
  signal place_336_rst : bit_vector(0 downto 0);
  signal place_336_top : bit;
  signal place_337_tip : bit_vector(0 downto 0);
  signal place_337_rst : bit_vector(0 downto 0);
  signal place_337_top : bit;
  signal place_338_tip : bit_vector(0 downto 0);
  signal place_338_rst : bit_vector(0 downto 0);
  signal place_338_top : bit;
  signal place_339_tip : bit_vector(0 downto 0);
  signal place_339_rst : bit_vector(0 downto 0);
  signal place_339_top : bit;
  signal place_340_tip : bit_vector(0 downto 0);
  signal place_340_rst : bit_vector(0 downto 0);
  signal place_340_top : bit;
  signal place_341_tip : bit_vector(0 downto 0);
  signal place_341_rst : bit_vector(0 downto 0);
  signal place_341_top : bit;
  signal place_342_tip : bit_vector(0 downto 0);
  signal place_342_rst : bit_vector(0 downto 0);
  signal place_342_top : bit;
  signal place_343_tip : bit_vector(0 downto 0);
  signal place_343_rst : bit_vector(0 downto 0);
  signal place_343_top : bit;
  signal place_344_tip : bit_vector(0 downto 0);
  signal place_344_rst : bit_vector(0 downto 0);
  signal place_344_top : bit;
  signal place_345_tip : bit_vector(0 downto 0);
  signal place_345_rst : bit_vector(0 downto 0);
  signal place_345_top : bit;
  signal place_346_tip : bit_vector(0 downto 0);
  signal place_346_rst : bit_vector(0 downto 0);
  signal place_346_top : bit;
  signal place_347_tip : bit_vector(0 downto 0);
  signal place_347_rst : bit_vector(0 downto 0);
  signal place_347_top : bit;
  signal place_349_tip : bit_vector(1 downto 0);
  signal place_349_rst : bit_vector(0 downto 0);
  signal place_349_top : bit;
  signal place_350_tip : bit_vector(0 downto 0);
  signal place_350_rst : bit_vector(0 downto 0);
  signal place_350_top : bit;
  signal place_351_tip : bit_vector(0 downto 0);
  signal place_351_rst : bit_vector(0 downto 0);
  signal place_351_top : bit;
  signal place_352_tip : bit_vector(0 downto 0);
  signal place_352_rst : bit_vector(0 downto 0);
  signal place_352_top : bit;
  signal place_354_tip : bit_vector(0 downto 0);
  signal place_354_rst : bit_vector(0 downto 0);
  signal place_354_top : bit;
  signal place_355_tip : bit_vector(0 downto 0);
  signal place_355_rst : bit_vector(0 downto 0);
  signal place_355_top : bit;
  signal place_356_tip : bit_vector(0 downto 0);
  signal place_356_rst : bit_vector(0 downto 0);
  signal place_356_top : bit;
  signal place_357_tip : bit_vector(0 downto 0);
  signal place_357_rst : bit_vector(0 downto 0);
  signal place_357_top : bit;
  signal place_358_tip : bit_vector(0 downto 0);
  signal place_358_rst : bit_vector(0 downto 0);
  signal place_358_top : bit;
  signal place_359_tip : bit_vector(0 downto 0);
  signal place_359_rst : bit_vector(0 downto 0);
  signal place_359_top : bit;
  signal place_36_tip : bit_vector(0 downto 0);
  signal place_36_rst : bit_vector(0 downto 0);
  signal place_36_top : bit;
  signal place_360_tip : bit_vector(0 downto 0);
  signal place_360_rst : bit_vector(0 downto 0);
  signal place_360_top : bit;
  signal place_361_tip : bit_vector(0 downto 0);
  signal place_361_rst : bit_vector(1 downto 0);
  signal place_361_top : bit;
  signal place_362_tip : bit_vector(0 downto 0);
  signal place_362_rst : bit_vector(0 downto 0);
  signal place_362_top : bit;
  signal place_363_tip : bit_vector(0 downto 0);
  signal place_363_rst : bit_vector(0 downto 0);
  signal place_363_top : bit;
  signal place_364_tip : bit_vector(0 downto 0);
  signal place_364_rst : bit_vector(0 downto 0);
  signal place_364_top : bit;
  signal place_365_tip : bit_vector(0 downto 0);
  signal place_365_rst : bit_vector(0 downto 0);
  signal place_365_top : bit;
  signal place_366_tip : bit_vector(0 downto 0);
  signal place_366_rst : bit_vector(0 downto 0);
  signal place_366_top : bit;
  signal place_367_tip : bit_vector(0 downto 0);
  signal place_367_rst : bit_vector(0 downto 0);
  signal place_367_top : bit;
  signal place_368_tip : bit_vector(0 downto 0);
  signal place_368_rst : bit_vector(0 downto 0);
  signal place_368_top : bit;
  signal place_369_tip : bit_vector(0 downto 0);
  signal place_369_rst : bit_vector(0 downto 0);
  signal place_369_top : bit;
  signal place_370_tip : bit_vector(0 downto 0);
  signal place_370_rst : bit_vector(0 downto 0);
  signal place_370_top : bit;
  signal place_371_tip : bit_vector(0 downto 0);
  signal place_371_rst : bit_vector(0 downto 0);
  signal place_371_top : bit;
  signal place_372_tip : bit_vector(0 downto 0);
  signal place_372_rst : bit_vector(0 downto 0);
  signal place_372_top : bit;
  signal place_373_tip : bit_vector(0 downto 0);
  signal place_373_rst : bit_vector(0 downto 0);
  signal place_373_top : bit;
  signal place_374_tip : bit_vector(0 downto 0);
  signal place_374_rst : bit_vector(0 downto 0);
  signal place_374_top : bit;
  signal place_375_tip : bit_vector(0 downto 0);
  signal place_375_rst : bit_vector(0 downto 0);
  signal place_375_top : bit;
  signal place_376_tip : bit_vector(0 downto 0);
  signal place_376_rst : bit_vector(0 downto 0);
  signal place_376_top : bit;
  signal place_377_tip : bit_vector(0 downto 0);
  signal place_377_rst : bit_vector(0 downto 0);
  signal place_377_top : bit;
  signal place_378_tip : bit_vector(0 downto 0);
  signal place_378_rst : bit_vector(0 downto 0);
  signal place_378_top : bit;
  signal place_379_tip : bit_vector(0 downto 0);
  signal place_379_rst : bit_vector(0 downto 0);
  signal place_379_top : bit;
  signal place_38_tip : bit_vector(0 downto 0);
  signal place_38_rst : bit_vector(0 downto 0);
  signal place_38_top : bit;
  signal place_380_tip : bit_vector(0 downto 0);
  signal place_380_rst : bit_vector(0 downto 0);
  signal place_380_top : bit;
  signal place_381_tip : bit_vector(0 downto 0);
  signal place_381_rst : bit_vector(0 downto 0);
  signal place_381_top : bit;
  signal place_382_tip : bit_vector(0 downto 0);
  signal place_382_rst : bit_vector(0 downto 0);
  signal place_382_top : bit;
  signal place_383_tip : bit_vector(0 downto 0);
  signal place_383_rst : bit_vector(0 downto 0);
  signal place_383_top : bit;
  signal place_384_tip : bit_vector(0 downto 0);
  signal place_384_rst : bit_vector(0 downto 0);
  signal place_384_top : bit;
  signal place_385_tip : bit_vector(0 downto 0);
  signal place_385_rst : bit_vector(0 downto 0);
  signal place_385_top : bit;
  signal place_386_tip : bit_vector(0 downto 0);
  signal place_386_rst : bit_vector(0 downto 0);
  signal place_386_top : bit;
  signal place_387_tip : bit_vector(0 downto 0);
  signal place_387_rst : bit_vector(0 downto 0);
  signal place_387_top : bit;
  signal place_388_tip : bit_vector(0 downto 0);
  signal place_388_rst : bit_vector(0 downto 0);
  signal place_388_top : bit;
  signal place_389_tip : bit_vector(0 downto 0);
  signal place_389_rst : bit_vector(0 downto 0);
  signal place_389_top : bit;
  signal place_390_tip : bit_vector(0 downto 0);
  signal place_390_rst : bit_vector(0 downto 0);
  signal place_390_top : bit;
  signal place_391_tip : bit_vector(0 downto 0);
  signal place_391_rst : bit_vector(1 downto 0);
  signal place_391_top : bit;
  signal place_392_tip : bit_vector(0 downto 0);
  signal place_392_rst : bit_vector(0 downto 0);
  signal place_392_top : bit;
  signal place_394_tip : bit_vector(0 downto 0);
  signal place_394_rst : bit_vector(0 downto 0);
  signal place_394_top : bit;
  signal place_396_tip : bit_vector(0 downto 0);
  signal place_396_rst : bit_vector(0 downto 0);
  signal place_396_top : bit;
  signal place_399_tip : bit_vector(1 downto 0);
  signal place_399_rst : bit_vector(0 downto 0);
  signal place_399_top : bit;
  signal place_40_tip : bit_vector(0 downto 0);
  signal place_40_rst : bit_vector(0 downto 0);
  signal place_40_top : bit;
  signal place_400_tip : bit_vector(0 downto 0);
  signal place_400_rst : bit_vector(0 downto 0);
  signal place_400_top : bit;
  signal place_401_tip : bit_vector(0 downto 0);
  signal place_401_rst : bit_vector(0 downto 0);
  signal place_401_top : bit;
  signal place_402_tip : bit_vector(0 downto 0);
  signal place_402_rst : bit_vector(0 downto 0);
  signal place_402_top : bit;
  signal place_403_tip : bit_vector(0 downto 0);
  signal place_403_rst : bit_vector(0 downto 0);
  signal place_403_top : bit;
  signal place_404_tip : bit_vector(0 downto 0);
  signal place_404_rst : bit_vector(0 downto 0);
  signal place_404_top : bit;
  signal place_405_tip : bit_vector(0 downto 0);
  signal place_405_rst : bit_vector(0 downto 0);
  signal place_405_top : bit;
  signal place_406_tip : bit_vector(0 downto 0);
  signal place_406_rst : bit_vector(0 downto 0);
  signal place_406_top : bit;
  signal place_407_tip : bit_vector(0 downto 0);
  signal place_407_rst : bit_vector(0 downto 0);
  signal place_407_top : bit;
  signal place_408_tip : bit_vector(0 downto 0);
  signal place_408_rst : bit_vector(0 downto 0);
  signal place_408_top : bit;
  signal place_409_tip : bit_vector(0 downto 0);
  signal place_409_rst : bit_vector(0 downto 0);
  signal place_409_top : bit;
  signal place_410_tip : bit_vector(0 downto 0);
  signal place_410_rst : bit_vector(0 downto 0);
  signal place_410_top : bit;
  signal place_411_tip : bit_vector(0 downto 0);
  signal place_411_rst : bit_vector(0 downto 0);
  signal place_411_top : bit;
  signal place_412_tip : bit_vector(0 downto 0);
  signal place_412_rst : bit_vector(0 downto 0);
  signal place_412_top : bit;
  signal place_413_tip : bit_vector(0 downto 0);
  signal place_413_rst : bit_vector(0 downto 0);
  signal place_413_top : bit;
  signal place_414_tip : bit_vector(0 downto 0);
  signal place_414_rst : bit_vector(0 downto 0);
  signal place_414_top : bit;
  signal place_415_tip : bit_vector(0 downto 0);
  signal place_415_rst : bit_vector(0 downto 0);
  signal place_415_top : bit;
  signal place_416_tip : bit_vector(0 downto 0);
  signal place_416_rst : bit_vector(0 downto 0);
  signal place_416_top : bit;
  signal place_417_tip : bit_vector(0 downto 0);
  signal place_417_rst : bit_vector(0 downto 0);
  signal place_417_top : bit;
  signal place_418_tip : bit_vector(0 downto 0);
  signal place_418_rst : bit_vector(0 downto 0);
  signal place_418_top : bit;
  signal place_419_tip : bit_vector(0 downto 0);
  signal place_419_rst : bit_vector(0 downto 0);
  signal place_419_top : bit;
  signal place_420_tip : bit_vector(0 downto 0);
  signal place_420_rst : bit_vector(0 downto 0);
  signal place_420_top : bit;
  signal place_421_tip : bit_vector(0 downto 0);
  signal place_421_rst : bit_vector(0 downto 0);
  signal place_421_top : bit;
  signal place_422_tip : bit_vector(0 downto 0);
  signal place_422_rst : bit_vector(0 downto 0);
  signal place_422_top : bit;
  signal place_423_tip : bit_vector(0 downto 0);
  signal place_423_rst : bit_vector(0 downto 0);
  signal place_423_top : bit;
  signal place_424_tip : bit_vector(0 downto 0);
  signal place_424_rst : bit_vector(0 downto 0);
  signal place_424_top : bit;
  signal place_425_tip : bit_vector(0 downto 0);
  signal place_425_rst : bit_vector(0 downto 0);
  signal place_425_top : bit;
  signal place_426_tip : bit_vector(0 downto 0);
  signal place_426_rst : bit_vector(0 downto 0);
  signal place_426_top : bit;
  signal place_427_tip : bit_vector(0 downto 0);
  signal place_427_rst : bit_vector(0 downto 0);
  signal place_427_top : bit;
  signal place_428_tip : bit_vector(0 downto 0);
  signal place_428_rst : bit_vector(0 downto 0);
  signal place_428_top : bit;
  signal place_429_tip : bit_vector(0 downto 0);
  signal place_429_rst : bit_vector(0 downto 0);
  signal place_429_top : bit;
  signal place_430_tip : bit_vector(0 downto 0);
  signal place_430_rst : bit_vector(0 downto 0);
  signal place_430_top : bit;
  signal place_431_tip : bit_vector(0 downto 0);
  signal place_431_rst : bit_vector(0 downto 0);
  signal place_431_top : bit;
  signal place_432_tip : bit_vector(0 downto 0);
  signal place_432_rst : bit_vector(0 downto 0);
  signal place_432_top : bit;
  signal place_433_tip : bit_vector(0 downto 0);
  signal place_433_rst : bit_vector(0 downto 0);
  signal place_433_top : bit;
  signal place_434_tip : bit_vector(0 downto 0);
  signal place_434_rst : bit_vector(0 downto 0);
  signal place_434_top : bit;
  signal place_435_tip : bit_vector(0 downto 0);
  signal place_435_rst : bit_vector(0 downto 0);
  signal place_435_top : bit;
  signal place_436_tip : bit_vector(0 downto 0);
  signal place_436_rst : bit_vector(0 downto 0);
  signal place_436_top : bit;
  signal place_437_tip : bit_vector(0 downto 0);
  signal place_437_rst : bit_vector(0 downto 0);
  signal place_437_top : bit;
  signal place_438_tip : bit_vector(0 downto 0);
  signal place_438_rst : bit_vector(0 downto 0);
  signal place_438_top : bit;
  signal place_439_tip : bit_vector(0 downto 0);
  signal place_439_rst : bit_vector(0 downto 0);
  signal place_439_top : bit;
  signal place_440_tip : bit_vector(0 downto 0);
  signal place_440_rst : bit_vector(0 downto 0);
  signal place_440_top : bit;
  signal place_441_tip : bit_vector(0 downto 0);
  signal place_441_rst : bit_vector(0 downto 0);
  signal place_441_top : bit;
  signal place_442_tip : bit_vector(0 downto 0);
  signal place_442_rst : bit_vector(0 downto 0);
  signal place_442_top : bit;
  signal place_443_tip : bit_vector(0 downto 0);
  signal place_443_rst : bit_vector(0 downto 0);
  signal place_443_top : bit;
  signal place_444_tip : bit_vector(0 downto 0);
  signal place_444_rst : bit_vector(0 downto 0);
  signal place_444_top : bit;
  signal place_445_tip : bit_vector(0 downto 0);
  signal place_445_rst : bit_vector(0 downto 0);
  signal place_445_top : bit;
  signal place_446_tip : bit_vector(0 downto 0);
  signal place_446_rst : bit_vector(0 downto 0);
  signal place_446_top : bit;
  signal place_447_tip : bit_vector(0 downto 0);
  signal place_447_rst : bit_vector(0 downto 0);
  signal place_447_top : bit;
  signal place_448_tip : bit_vector(0 downto 0);
  signal place_448_rst : bit_vector(0 downto 0);
  signal place_448_top : bit;
  signal place_449_tip : bit_vector(0 downto 0);
  signal place_449_rst : bit_vector(1 downto 0);
  signal place_449_top : bit;
  signal place_450_tip : bit_vector(0 downto 0);
  signal place_450_rst : bit_vector(0 downto 0);
  signal place_450_top : bit;
  signal place_451_tip : bit_vector(0 downto 0);
  signal place_451_rst : bit_vector(0 downto 0);
  signal place_451_top : bit;
  signal place_453_tip : bit_vector(0 downto 0);
  signal place_453_rst : bit_vector(0 downto 0);
  signal place_453_top : bit;
  signal place_454_tip : bit_vector(0 downto 0);
  signal place_454_rst : bit_vector(1 downto 0);
  signal place_454_top : bit;
  signal place_457_tip : bit_vector(1 downto 0);
  signal place_457_rst : bit_vector(0 downto 0);
  signal place_457_top : bit;
  signal place_458_tip : bit_vector(0 downto 0);
  signal place_458_rst : bit_vector(0 downto 0);
  signal place_458_top : bit;
  signal place_459_tip : bit_vector(0 downto 0);
  signal place_459_rst : bit_vector(0 downto 0);
  signal place_459_top : bit;
  signal place_46_tip : bit_vector(1 downto 0);
  signal place_46_rst : bit_vector(0 downto 0);
  signal place_46_top : bit;
  signal place_460_tip : bit_vector(0 downto 0);
  signal place_460_rst : bit_vector(0 downto 0);
  signal place_460_top : bit;
  signal place_462_tip : bit_vector(0 downto 0);
  signal place_462_rst : bit_vector(0 downto 0);
  signal place_462_top : bit;
  signal place_464_tip : bit_vector(1 downto 0);
  signal place_464_rst : bit_vector(0 downto 0);
  signal place_464_top : bit;
  signal place_465_tip : bit_vector(0 downto 0);
  signal place_465_rst : bit_vector(0 downto 0);
  signal place_465_top : bit;
  signal place_467_tip : bit_vector(0 downto 0);
  signal place_467_rst : bit_vector(0 downto 0);
  signal place_467_top : bit;
  signal place_469_tip : bit_vector(0 downto 0);
  signal place_469_rst : bit_vector(0 downto 0);
  signal place_469_top : bit;
  signal place_470_tip : bit_vector(0 downto 0);
  signal place_470_rst : bit_vector(1 downto 0);
  signal place_470_top : bit;
  signal place_471_tip : bit_vector(0 downto 0);
  signal place_471_rst : bit_vector(0 downto 0);
  signal place_471_top : bit;
  signal place_472_tip : bit_vector(0 downto 0);
  signal place_472_rst : bit_vector(0 downto 0);
  signal place_472_top : bit;
  signal place_473_tip : bit_vector(0 downto 0);
  signal place_473_rst : bit_vector(0 downto 0);
  signal place_473_top : bit;
  signal place_474_tip : bit_vector(0 downto 0);
  signal place_474_rst : bit_vector(0 downto 0);
  signal place_474_top : bit;
  signal place_475_tip : bit_vector(0 downto 0);
  signal place_475_rst : bit_vector(0 downto 0);
  signal place_475_top : bit;
  signal place_476_tip : bit_vector(0 downto 0);
  signal place_476_rst : bit_vector(0 downto 0);
  signal place_476_top : bit;
  signal place_477_tip : bit_vector(0 downto 0);
  signal place_477_rst : bit_vector(0 downto 0);
  signal place_477_top : bit;
  signal place_478_tip : bit_vector(0 downto 0);
  signal place_478_rst : bit_vector(0 downto 0);
  signal place_478_top : bit;
  signal place_479_tip : bit_vector(0 downto 0);
  signal place_479_rst : bit_vector(0 downto 0);
  signal place_479_top : bit;
  signal place_48_tip : bit_vector(0 downto 0);
  signal place_48_rst : bit_vector(0 downto 0);
  signal place_48_top : bit;
  signal place_480_tip : bit_vector(0 downto 0);
  signal place_480_rst : bit_vector(0 downto 0);
  signal place_480_top : bit;
  signal place_481_tip : bit_vector(0 downto 0);
  signal place_481_rst : bit_vector(0 downto 0);
  signal place_481_top : bit;
  signal place_482_tip : bit_vector(0 downto 0);
  signal place_482_rst : bit_vector(0 downto 0);
  signal place_482_top : bit;
  signal place_483_tip : bit_vector(0 downto 0);
  signal place_483_rst : bit_vector(0 downto 0);
  signal place_483_top : bit;
  signal place_484_tip : bit_vector(0 downto 0);
  signal place_484_rst : bit_vector(0 downto 0);
  signal place_484_top : bit;
  signal place_485_tip : bit_vector(0 downto 0);
  signal place_485_rst : bit_vector(0 downto 0);
  signal place_485_top : bit;
  signal place_486_tip : bit_vector(0 downto 0);
  signal place_486_rst : bit_vector(0 downto 0);
  signal place_486_top : bit;
  signal place_487_tip : bit_vector(0 downto 0);
  signal place_487_rst : bit_vector(0 downto 0);
  signal place_487_top : bit;
  signal place_488_tip : bit_vector(0 downto 0);
  signal place_488_rst : bit_vector(0 downto 0);
  signal place_488_top : bit;
  signal place_489_tip : bit_vector(0 downto 0);
  signal place_489_rst : bit_vector(0 downto 0);
  signal place_489_top : bit;
  signal place_490_tip : bit_vector(0 downto 0);
  signal place_490_rst : bit_vector(0 downto 0);
  signal place_490_top : bit;
  signal place_491_tip : bit_vector(0 downto 0);
  signal place_491_rst : bit_vector(0 downto 0);
  signal place_491_top : bit;
  signal place_492_tip : bit_vector(0 downto 0);
  signal place_492_rst : bit_vector(0 downto 0);
  signal place_492_top : bit;
  signal place_493_tip : bit_vector(0 downto 0);
  signal place_493_rst : bit_vector(0 downto 0);
  signal place_493_top : bit;
  signal place_494_tip : bit_vector(0 downto 0);
  signal place_494_rst : bit_vector(0 downto 0);
  signal place_494_top : bit;
  signal place_495_tip : bit_vector(0 downto 0);
  signal place_495_rst : bit_vector(0 downto 0);
  signal place_495_top : bit;
  signal place_496_tip : bit_vector(0 downto 0);
  signal place_496_rst : bit_vector(0 downto 0);
  signal place_496_top : bit;
  signal place_497_tip : bit_vector(0 downto 0);
  signal place_497_rst : bit_vector(0 downto 0);
  signal place_497_top : bit;
  signal place_498_tip : bit_vector(0 downto 0);
  signal place_498_rst : bit_vector(0 downto 0);
  signal place_498_top : bit;
  signal place_499_tip : bit_vector(0 downto 0);
  signal place_499_rst : bit_vector(0 downto 0);
  signal place_499_top : bit;
  signal place_5_tip : bit_vector(0 downto 0);
  signal place_5_rst : bit_vector(0 downto 0);
  signal place_5_top : bit;
  signal place_500_tip : bit_vector(0 downto 0);
  signal place_500_rst : bit_vector(0 downto 0);
  signal place_500_top : bit;
  signal place_501_tip : bit_vector(0 downto 0);
  signal place_501_rst : bit_vector(0 downto 0);
  signal place_501_top : bit;
  signal place_502_tip : bit_vector(0 downto 0);
  signal place_502_rst : bit_vector(0 downto 0);
  signal place_502_top : bit;
  signal place_503_tip : bit_vector(0 downto 0);
  signal place_503_rst : bit_vector(0 downto 0);
  signal place_503_top : bit;
  signal place_504_tip : bit_vector(0 downto 0);
  signal place_504_rst : bit_vector(0 downto 0);
  signal place_504_top : bit;
  signal place_505_tip : bit_vector(0 downto 0);
  signal place_505_rst : bit_vector(0 downto 0);
  signal place_505_top : bit;
  signal place_506_tip : bit_vector(0 downto 0);
  signal place_506_rst : bit_vector(0 downto 0);
  signal place_506_top : bit;
  signal place_507_tip : bit_vector(0 downto 0);
  signal place_507_rst : bit_vector(0 downto 0);
  signal place_507_top : bit;
  signal place_508_tip : bit_vector(0 downto 0);
  signal place_508_rst : bit_vector(0 downto 0);
  signal place_508_top : bit;
  signal place_509_tip : bit_vector(0 downto 0);
  signal place_509_rst : bit_vector(0 downto 0);
  signal place_509_top : bit;
  signal place_510_tip : bit_vector(0 downto 0);
  signal place_510_rst : bit_vector(0 downto 0);
  signal place_510_top : bit;
  signal place_511_tip : bit_vector(0 downto 0);
  signal place_511_rst : bit_vector(0 downto 0);
  signal place_511_top : bit;
  signal place_512_tip : bit_vector(0 downto 0);
  signal place_512_rst : bit_vector(0 downto 0);
  signal place_512_top : bit;
  signal place_513_tip : bit_vector(0 downto 0);
  signal place_513_rst : bit_vector(0 downto 0);
  signal place_513_top : bit;
  signal place_514_tip : bit_vector(0 downto 0);
  signal place_514_rst : bit_vector(1 downto 0);
  signal place_514_top : bit;
  signal place_515_tip : bit_vector(0 downto 0);
  signal place_515_rst : bit_vector(0 downto 0);
  signal place_515_top : bit;
  signal place_516_tip : bit_vector(0 downto 0);
  signal place_516_rst : bit_vector(0 downto 0);
  signal place_516_top : bit;
  signal place_517_tip : bit_vector(1 downto 0);
  signal place_517_rst : bit_vector(0 downto 0);
  signal place_517_top : bit;
  signal place_518_tip : bit_vector(0 downto 0);
  signal place_518_rst : bit_vector(0 downto 0);
  signal place_518_top : bit;
  signal place_519_tip : bit_vector(0 downto 0);
  signal place_519_rst : bit_vector(0 downto 0);
  signal place_519_top : bit;
  signal place_52_tip : bit_vector(0 downto 0);
  signal place_52_rst : bit_vector(0 downto 0);
  signal place_52_top : bit;
  signal place_520_tip : bit_vector(1 downto 0);
  signal place_520_rst : bit_vector(0 downto 0);
  signal place_520_top : bit;
  signal place_521_tip : bit_vector(0 downto 0);
  signal place_521_rst : bit_vector(0 downto 0);
  signal place_521_top : bit;
  signal place_522_tip : bit_vector(0 downto 0);
  signal place_522_rst : bit_vector(0 downto 0);
  signal place_522_top : bit;
  signal place_524_tip : bit_vector(0 downto 0);
  signal place_524_rst : bit_vector(0 downto 0);
  signal place_524_top : bit;
  signal place_525_tip : bit_vector(0 downto 0);
  signal place_525_rst : bit_vector(0 downto 0);
  signal place_525_top : bit;
  signal place_526_tip : bit_vector(0 downto 0);
  signal place_526_rst : bit_vector(0 downto 0);
  signal place_526_top : bit;
  signal place_527_tip : bit_vector(0 downto 0);
  signal place_527_rst : bit_vector(0 downto 0);
  signal place_527_top : bit;
  signal place_528_tip : bit_vector(0 downto 0);
  signal place_528_rst : bit_vector(0 downto 0);
  signal place_528_top : bit;
  signal place_529_tip : bit_vector(0 downto 0);
  signal place_529_rst : bit_vector(0 downto 0);
  signal place_529_top : bit;
  signal place_530_tip : bit_vector(0 downto 0);
  signal place_530_rst : bit_vector(0 downto 0);
  signal place_530_top : bit;
  signal place_531_tip : bit_vector(0 downto 0);
  signal place_531_rst : bit_vector(0 downto 0);
  signal place_531_top : bit;
  signal place_532_tip : bit_vector(0 downto 0);
  signal place_532_rst : bit_vector(0 downto 0);
  signal place_532_top : bit;
  signal place_533_tip : bit_vector(0 downto 0);
  signal place_533_rst : bit_vector(0 downto 0);
  signal place_533_top : bit;
  signal place_534_tip : bit_vector(0 downto 0);
  signal place_534_rst : bit_vector(0 downto 0);
  signal place_534_top : bit;
  signal place_535_tip : bit_vector(0 downto 0);
  signal place_535_rst : bit_vector(0 downto 0);
  signal place_535_top : bit;
  signal place_536_tip : bit_vector(0 downto 0);
  signal place_536_rst : bit_vector(0 downto 0);
  signal place_536_top : bit;
  signal place_537_tip : bit_vector(0 downto 0);
  signal place_537_rst : bit_vector(1 downto 0);
  signal place_537_top : bit;
  signal place_538_tip : bit_vector(0 downto 0);
  signal place_538_rst : bit_vector(0 downto 0);
  signal place_538_top : bit;
  signal place_539_tip : bit_vector(0 downto 0);
  signal place_539_rst : bit_vector(0 downto 0);
  signal place_539_top : bit;
  signal place_54_tip : bit_vector(0 downto 0);
  signal place_54_rst : bit_vector(0 downto 0);
  signal place_54_top : bit;
  signal place_540_tip : bit_vector(0 downto 0);
  signal place_540_rst : bit_vector(0 downto 0);
  signal place_540_top : bit;
  signal place_541_tip : bit_vector(0 downto 0);
  signal place_541_rst : bit_vector(0 downto 0);
  signal place_541_top : bit;
  signal place_542_tip : bit_vector(0 downto 0);
  signal place_542_rst : bit_vector(0 downto 0);
  signal place_542_top : bit;
  signal place_543_tip : bit_vector(0 downto 0);
  signal place_543_rst : bit_vector(0 downto 0);
  signal place_543_top : bit;
  signal place_544_tip : bit_vector(0 downto 0);
  signal place_544_rst : bit_vector(0 downto 0);
  signal place_544_top : bit;
  signal place_545_tip : bit_vector(0 downto 0);
  signal place_545_rst : bit_vector(0 downto 0);
  signal place_545_top : bit;
  signal place_546_tip : bit_vector(0 downto 0);
  signal place_546_rst : bit_vector(0 downto 0);
  signal place_546_top : bit;
  signal place_547_tip : bit_vector(0 downto 0);
  signal place_547_rst : bit_vector(0 downto 0);
  signal place_547_top : bit;
  signal place_548_tip : bit_vector(0 downto 0);
  signal place_548_rst : bit_vector(0 downto 0);
  signal place_548_top : bit;
  signal place_549_tip : bit_vector(0 downto 0);
  signal place_549_rst : bit_vector(0 downto 0);
  signal place_549_top : bit;
  signal place_550_tip : bit_vector(0 downto 0);
  signal place_550_rst : bit_vector(0 downto 0);
  signal place_550_top : bit;
  signal place_551_tip : bit_vector(0 downto 0);
  signal place_551_rst : bit_vector(0 downto 0);
  signal place_551_top : bit;
  signal place_552_tip : bit_vector(0 downto 0);
  signal place_552_rst : bit_vector(0 downto 0);
  signal place_552_top : bit;
  signal place_553_tip : bit_vector(0 downto 0);
  signal place_553_rst : bit_vector(0 downto 0);
  signal place_553_top : bit;
  signal place_554_tip : bit_vector(0 downto 0);
  signal place_554_rst : bit_vector(0 downto 0);
  signal place_554_top : bit;
  signal place_555_tip : bit_vector(0 downto 0);
  signal place_555_rst : bit_vector(0 downto 0);
  signal place_555_top : bit;
  signal place_556_tip : bit_vector(0 downto 0);
  signal place_556_rst : bit_vector(0 downto 0);
  signal place_556_top : bit;
  signal place_557_tip : bit_vector(0 downto 0);
  signal place_557_rst : bit_vector(0 downto 0);
  signal place_557_top : bit;
  signal place_558_tip : bit_vector(0 downto 0);
  signal place_558_rst : bit_vector(0 downto 0);
  signal place_558_top : bit;
  signal place_559_tip : bit_vector(0 downto 0);
  signal place_559_rst : bit_vector(0 downto 0);
  signal place_559_top : bit;
  signal place_560_tip : bit_vector(0 downto 0);
  signal place_560_rst : bit_vector(0 downto 0);
  signal place_560_top : bit;
  signal place_561_tip : bit_vector(0 downto 0);
  signal place_561_rst : bit_vector(0 downto 0);
  signal place_561_top : bit;
  signal place_562_tip : bit_vector(0 downto 0);
  signal place_562_rst : bit_vector(0 downto 0);
  signal place_562_top : bit;
  signal place_563_tip : bit_vector(0 downto 0);
  signal place_563_rst : bit_vector(0 downto 0);
  signal place_563_top : bit;
  signal place_564_tip : bit_vector(0 downto 0);
  signal place_564_rst : bit_vector(0 downto 0);
  signal place_564_top : bit;
  signal place_565_tip : bit_vector(0 downto 0);
  signal place_565_rst : bit_vector(0 downto 0);
  signal place_565_top : bit;
  signal place_566_tip : bit_vector(0 downto 0);
  signal place_566_rst : bit_vector(0 downto 0);
  signal place_566_top : bit;
  signal place_567_tip : bit_vector(0 downto 0);
  signal place_567_rst : bit_vector(0 downto 0);
  signal place_567_top : bit;
  signal place_568_tip : bit_vector(0 downto 0);
  signal place_568_rst : bit_vector(0 downto 0);
  signal place_568_top : bit;
  signal place_569_tip : bit_vector(0 downto 0);
  signal place_569_rst : bit_vector(0 downto 0);
  signal place_569_top : bit;
  signal place_570_tip : bit_vector(0 downto 0);
  signal place_570_rst : bit_vector(0 downto 0);
  signal place_570_top : bit;
  signal place_571_tip : bit_vector(0 downto 0);
  signal place_571_rst : bit_vector(0 downto 0);
  signal place_571_top : bit;
  signal place_572_tip : bit_vector(0 downto 0);
  signal place_572_rst : bit_vector(1 downto 0);
  signal place_572_top : bit;
  signal place_573_tip : bit_vector(0 downto 0);
  signal place_573_rst : bit_vector(0 downto 0);
  signal place_573_top : bit;
  signal place_574_tip : bit_vector(0 downto 0);
  signal place_574_rst : bit_vector(0 downto 0);
  signal place_574_top : bit;
  signal place_575_tip : bit_vector(0 downto 0);
  signal place_575_rst : bit_vector(0 downto 0);
  signal place_575_top : bit;
  signal place_576_tip : bit_vector(0 downto 0);
  signal place_576_rst : bit_vector(0 downto 0);
  signal place_576_top : bit;
  signal place_577_tip : bit_vector(0 downto 0);
  signal place_577_rst : bit_vector(0 downto 0);
  signal place_577_top : bit;
  signal place_578_tip : bit_vector(0 downto 0);
  signal place_578_rst : bit_vector(0 downto 0);
  signal place_578_top : bit;
  signal place_579_tip : bit_vector(0 downto 0);
  signal place_579_rst : bit_vector(0 downto 0);
  signal place_579_top : bit;
  signal place_580_tip : bit_vector(0 downto 0);
  signal place_580_rst : bit_vector(0 downto 0);
  signal place_580_top : bit;
  signal place_581_tip : bit_vector(0 downto 0);
  signal place_581_rst : bit_vector(0 downto 0);
  signal place_581_top : bit;
  signal place_582_tip : bit_vector(0 downto 0);
  signal place_582_rst : bit_vector(0 downto 0);
  signal place_582_top : bit;
  signal place_583_tip : bit_vector(0 downto 0);
  signal place_583_rst : bit_vector(0 downto 0);
  signal place_583_top : bit;
  signal place_584_tip : bit_vector(0 downto 0);
  signal place_584_rst : bit_vector(0 downto 0);
  signal place_584_top : bit;
  signal place_585_tip : bit_vector(0 downto 0);
  signal place_585_rst : bit_vector(0 downto 0);
  signal place_585_top : bit;
  signal place_586_tip : bit_vector(0 downto 0);
  signal place_586_rst : bit_vector(0 downto 0);
  signal place_586_top : bit;
  signal place_587_tip : bit_vector(0 downto 0);
  signal place_587_rst : bit_vector(0 downto 0);
  signal place_587_top : bit;
  signal place_588_tip : bit_vector(0 downto 0);
  signal place_588_rst : bit_vector(0 downto 0);
  signal place_588_top : bit;
  signal place_589_tip : bit_vector(0 downto 0);
  signal place_589_rst : bit_vector(0 downto 0);
  signal place_589_top : bit;
  signal place_59_tip : bit_vector(0 downto 0);
  signal place_59_rst : bit_vector(0 downto 0);
  signal place_59_top : bit;
  signal place_590_tip : bit_vector(0 downto 0);
  signal place_590_rst : bit_vector(0 downto 0);
  signal place_590_top : bit;
  signal place_591_tip : bit_vector(0 downto 0);
  signal place_591_rst : bit_vector(0 downto 0);
  signal place_591_top : bit;
  signal place_592_tip : bit_vector(0 downto 0);
  signal place_592_rst : bit_vector(0 downto 0);
  signal place_592_top : bit;
  signal place_593_tip : bit_vector(0 downto 0);
  signal place_593_rst : bit_vector(0 downto 0);
  signal place_593_top : bit;
  signal place_594_tip : bit_vector(0 downto 0);
  signal place_594_rst : bit_vector(0 downto 0);
  signal place_594_top : bit;
  signal place_595_tip : bit_vector(0 downto 0);
  signal place_595_rst : bit_vector(0 downto 0);
  signal place_595_top : bit;
  signal place_596_tip : bit_vector(0 downto 0);
  signal place_596_rst : bit_vector(0 downto 0);
  signal place_596_top : bit;
  signal place_597_tip : bit_vector(0 downto 0);
  signal place_597_rst : bit_vector(0 downto 0);
  signal place_597_top : bit;
  signal place_598_tip : bit_vector(0 downto 0);
  signal place_598_rst : bit_vector(0 downto 0);
  signal place_598_top : bit;
  signal place_599_tip : bit_vector(0 downto 0);
  signal place_599_rst : bit_vector(0 downto 0);
  signal place_599_top : bit;
  signal place_600_tip : bit_vector(0 downto 0);
  signal place_600_rst : bit_vector(0 downto 0);
  signal place_600_top : bit;
  signal place_601_tip : bit_vector(0 downto 0);
  signal place_601_rst : bit_vector(0 downto 0);
  signal place_601_top : bit;
  signal place_602_tip : bit_vector(0 downto 0);
  signal place_602_rst : bit_vector(0 downto 0);
  signal place_602_top : bit;
  signal place_603_tip : bit_vector(0 downto 0);
  signal place_603_rst : bit_vector(0 downto 0);
  signal place_603_top : bit;
  signal place_604_tip : bit_vector(0 downto 0);
  signal place_604_rst : bit_vector(0 downto 0);
  signal place_604_top : bit;
  signal place_605_tip : bit_vector(0 downto 0);
  signal place_605_rst : bit_vector(0 downto 0);
  signal place_605_top : bit;
  signal place_606_tip : bit_vector(0 downto 0);
  signal place_606_rst : bit_vector(0 downto 0);
  signal place_606_top : bit;
  signal place_607_tip : bit_vector(0 downto 0);
  signal place_607_rst : bit_vector(0 downto 0);
  signal place_607_top : bit;
  signal place_608_tip : bit_vector(0 downto 0);
  signal place_608_rst : bit_vector(1 downto 0);
  signal place_608_top : bit;
  signal place_609_tip : bit_vector(0 downto 0);
  signal place_609_rst : bit_vector(0 downto 0);
  signal place_609_top : bit;
  signal place_61_tip : bit_vector(0 downto 0);
  signal place_61_rst : bit_vector(0 downto 0);
  signal place_61_top : bit;
  signal place_610_tip : bit_vector(0 downto 0);
  signal place_610_rst : bit_vector(0 downto 0);
  signal place_610_top : bit;
  signal place_612_tip : bit_vector(0 downto 0);
  signal place_612_rst : bit_vector(0 downto 0);
  signal place_612_top : bit;
  signal place_613_tip : bit_vector(0 downto 0);
  signal place_613_rst : bit_vector(0 downto 0);
  signal place_613_top : bit;
  signal place_614_tip : bit_vector(0 downto 0);
  signal place_614_rst : bit_vector(0 downto 0);
  signal place_614_top : bit;
  signal place_615_tip : bit_vector(0 downto 0);
  signal place_615_rst : bit_vector(1 downto 0);
  signal place_615_top : bit;
  signal place_617_tip : bit_vector(0 downto 0);
  signal place_617_rst : bit_vector(0 downto 0);
  signal place_617_top : bit;
  signal place_618_tip : bit_vector(1 downto 0);
  signal place_618_rst : bit_vector(0 downto 0);
  signal place_618_top : bit;
  signal place_619_tip : bit_vector(0 downto 0);
  signal place_619_rst : bit_vector(0 downto 0);
  signal place_619_top : bit;
  signal place_620_tip : bit_vector(0 downto 0);
  signal place_620_rst : bit_vector(0 downto 0);
  signal place_620_top : bit;
  signal place_621_tip : bit_vector(0 downto 0);
  signal place_621_rst : bit_vector(0 downto 0);
  signal place_621_top : bit;
  signal place_622_tip : bit_vector(1 downto 0);
  signal place_622_rst : bit_vector(0 downto 0);
  signal place_622_top : bit;
  signal place_623_tip : bit_vector(0 downto 0);
  signal place_623_rst : bit_vector(0 downto 0);
  signal place_623_top : bit;
  signal place_624_tip : bit_vector(0 downto 0);
  signal place_624_rst : bit_vector(0 downto 0);
  signal place_624_top : bit;
  signal place_625_tip : bit_vector(0 downto 0);
  signal place_625_rst : bit_vector(0 downto 0);
  signal place_625_top : bit;
  signal place_626_tip : bit_vector(0 downto 0);
  signal place_626_rst : bit_vector(0 downto 0);
  signal place_626_top : bit;
  signal place_627_tip : bit_vector(0 downto 0);
  signal place_627_rst : bit_vector(0 downto 0);
  signal place_627_top : bit;
  signal place_628_tip : bit_vector(0 downto 0);
  signal place_628_rst : bit_vector(0 downto 0);
  signal place_628_top : bit;
  signal place_629_tip : bit_vector(0 downto 0);
  signal place_629_rst : bit_vector(0 downto 0);
  signal place_629_top : bit;
  signal place_63_tip : bit_vector(2 downto 0);
  signal place_63_rst : bit_vector(0 downto 0);
  signal place_63_top : bit;
  signal place_630_tip : bit_vector(0 downto 0);
  signal place_630_rst : bit_vector(0 downto 0);
  signal place_630_top : bit;
  signal place_631_tip : bit_vector(0 downto 0);
  signal place_631_rst : bit_vector(0 downto 0);
  signal place_631_top : bit;
  signal place_632_tip : bit_vector(0 downto 0);
  signal place_632_rst : bit_vector(1 downto 0);
  signal place_632_top : bit;
  signal place_635_tip : bit_vector(1 downto 0);
  signal place_635_rst : bit_vector(0 downto 0);
  signal place_635_top : bit;
  signal place_636_tip : bit_vector(0 downto 0);
  signal place_636_rst : bit_vector(0 downto 0);
  signal place_636_top : bit;
  signal place_637_tip : bit_vector(0 downto 0);
  signal place_637_rst : bit_vector(0 downto 0);
  signal place_637_top : bit;
  signal place_638_tip : bit_vector(0 downto 0);
  signal place_638_rst : bit_vector(0 downto 0);
  signal place_638_top : bit;
  signal place_639_tip : bit_vector(0 downto 0);
  signal place_639_rst : bit_vector(0 downto 0);
  signal place_639_top : bit;
  signal place_640_tip : bit_vector(0 downto 0);
  signal place_640_rst : bit_vector(0 downto 0);
  signal place_640_top : bit;
  signal place_641_tip : bit_vector(0 downto 0);
  signal place_641_rst : bit_vector(0 downto 0);
  signal place_641_top : bit;
  signal place_642_tip : bit_vector(0 downto 0);
  signal place_642_rst : bit_vector(0 downto 0);
  signal place_642_top : bit;
  signal place_643_tip : bit_vector(0 downto 0);
  signal place_643_rst : bit_vector(0 downto 0);
  signal place_643_top : bit;
  signal place_644_tip : bit_vector(0 downto 0);
  signal place_644_rst : bit_vector(0 downto 0);
  signal place_644_top : bit;
  signal place_645_tip : bit_vector(0 downto 0);
  signal place_645_rst : bit_vector(0 downto 0);
  signal place_645_top : bit;
  signal place_646_tip : bit_vector(0 downto 0);
  signal place_646_rst : bit_vector(0 downto 0);
  signal place_646_top : bit;
  signal place_647_tip : bit_vector(0 downto 0);
  signal place_647_rst : bit_vector(0 downto 0);
  signal place_647_top : bit;
  signal place_648_tip : bit_vector(0 downto 0);
  signal place_648_rst : bit_vector(0 downto 0);
  signal place_648_top : bit;
  signal place_649_tip : bit_vector(0 downto 0);
  signal place_649_rst : bit_vector(0 downto 0);
  signal place_649_top : bit;
  signal place_65_tip : bit_vector(0 downto 0);
  signal place_65_rst : bit_vector(0 downto 0);
  signal place_65_top : bit;
  signal place_650_tip : bit_vector(0 downto 0);
  signal place_650_rst : bit_vector(0 downto 0);
  signal place_650_top : bit;
  signal place_651_tip : bit_vector(0 downto 0);
  signal place_651_rst : bit_vector(0 downto 0);
  signal place_651_top : bit;
  signal place_652_tip : bit_vector(0 downto 0);
  signal place_652_rst : bit_vector(0 downto 0);
  signal place_652_top : bit;
  signal place_653_tip : bit_vector(0 downto 0);
  signal place_653_rst : bit_vector(0 downto 0);
  signal place_653_top : bit;
  signal place_654_tip : bit_vector(0 downto 0);
  signal place_654_rst : bit_vector(0 downto 0);
  signal place_654_top : bit;
  signal place_655_tip : bit_vector(0 downto 0);
  signal place_655_rst : bit_vector(0 downto 0);
  signal place_655_top : bit;
  signal place_656_tip : bit_vector(0 downto 0);
  signal place_656_rst : bit_vector(0 downto 0);
  signal place_656_top : bit;
  signal place_657_tip : bit_vector(0 downto 0);
  signal place_657_rst : bit_vector(0 downto 0);
  signal place_657_top : bit;
  signal place_658_tip : bit_vector(0 downto 0);
  signal place_658_rst : bit_vector(0 downto 0);
  signal place_658_top : bit;
  signal place_659_tip : bit_vector(0 downto 0);
  signal place_659_rst : bit_vector(0 downto 0);
  signal place_659_top : bit;
  signal place_66_tip : bit_vector(0 downto 0);
  signal place_66_rst : bit_vector(0 downto 0);
  signal place_66_top : bit;
  signal place_660_tip : bit_vector(0 downto 0);
  signal place_660_rst : bit_vector(0 downto 0);
  signal place_660_top : bit;
  signal place_661_tip : bit_vector(0 downto 0);
  signal place_661_rst : bit_vector(0 downto 0);
  signal place_661_top : bit;
  signal place_662_tip : bit_vector(0 downto 0);
  signal place_662_rst : bit_vector(0 downto 0);
  signal place_662_top : bit;
  signal place_663_tip : bit_vector(0 downto 0);
  signal place_663_rst : bit_vector(0 downto 0);
  signal place_663_top : bit;
  signal place_664_tip : bit_vector(0 downto 0);
  signal place_664_rst : bit_vector(0 downto 0);
  signal place_664_top : bit;
  signal place_665_tip : bit_vector(0 downto 0);
  signal place_665_rst : bit_vector(0 downto 0);
  signal place_665_top : bit;
  signal place_666_tip : bit_vector(0 downto 0);
  signal place_666_rst : bit_vector(0 downto 0);
  signal place_666_top : bit;
  signal place_667_tip : bit_vector(0 downto 0);
  signal place_667_rst : bit_vector(1 downto 0);
  signal place_667_top : bit;
  signal place_668_tip : bit_vector(0 downto 0);
  signal place_668_rst : bit_vector(0 downto 0);
  signal place_668_top : bit;
  signal place_669_tip : bit_vector(0 downto 0);
  signal place_669_rst : bit_vector(0 downto 0);
  signal place_669_top : bit;
  signal place_671_tip : bit_vector(0 downto 0);
  signal place_671_rst : bit_vector(0 downto 0);
  signal place_671_top : bit;
  signal place_673_tip : bit_vector(1 downto 0);
  signal place_673_rst : bit_vector(0 downto 0);
  signal place_673_top : bit;
  signal place_674_tip : bit_vector(0 downto 0);
  signal place_674_rst : bit_vector(0 downto 0);
  signal place_674_top : bit;
  signal place_675_tip : bit_vector(0 downto 0);
  signal place_675_rst : bit_vector(0 downto 0);
  signal place_675_top : bit;
  signal place_676_tip : bit_vector(0 downto 0);
  signal place_676_rst : bit_vector(0 downto 0);
  signal place_676_top : bit;
  signal place_677_tip : bit_vector(0 downto 0);
  signal place_677_rst : bit_vector(0 downto 0);
  signal place_677_top : bit;
  signal place_678_tip : bit_vector(0 downto 0);
  signal place_678_rst : bit_vector(0 downto 0);
  signal place_678_top : bit;
  signal place_679_tip : bit_vector(0 downto 0);
  signal place_679_rst : bit_vector(0 downto 0);
  signal place_679_top : bit;
  signal place_680_tip : bit_vector(0 downto 0);
  signal place_680_rst : bit_vector(0 downto 0);
  signal place_680_top : bit;
  signal place_681_tip : bit_vector(0 downto 0);
  signal place_681_rst : bit_vector(0 downto 0);
  signal place_681_top : bit;
  signal place_682_tip : bit_vector(0 downto 0);
  signal place_682_rst : bit_vector(1 downto 0);
  signal place_682_top : bit;
  signal place_684_tip : bit_vector(0 downto 0);
  signal place_684_rst : bit_vector(0 downto 0);
  signal place_684_top : bit;
  signal place_685_tip : bit_vector(1 downto 0);
  signal place_685_rst : bit_vector(0 downto 0);
  signal place_685_top : bit;
  signal place_686_tip : bit_vector(0 downto 0);
  signal place_686_rst : bit_vector(0 downto 0);
  signal place_686_top : bit;
  signal place_687_tip : bit_vector(0 downto 0);
  signal place_687_rst : bit_vector(0 downto 0);
  signal place_687_top : bit;
  signal place_688_tip : bit_vector(0 downto 0);
  signal place_688_rst : bit_vector(0 downto 0);
  signal place_688_top : bit;
  signal place_689_tip : bit_vector(1 downto 0);
  signal place_689_rst : bit_vector(0 downto 0);
  signal place_689_top : bit;
  signal place_69_tip : bit_vector(0 downto 0);
  signal place_69_rst : bit_vector(0 downto 0);
  signal place_69_top : bit;
  signal place_690_tip : bit_vector(0 downto 0);
  signal place_690_rst : bit_vector(0 downto 0);
  signal place_690_top : bit;
  signal place_691_tip : bit_vector(0 downto 0);
  signal place_691_rst : bit_vector(0 downto 0);
  signal place_691_top : bit;
  signal place_692_tip : bit_vector(0 downto 0);
  signal place_692_rst : bit_vector(0 downto 0);
  signal place_692_top : bit;
  signal place_693_tip : bit_vector(0 downto 0);
  signal place_693_rst : bit_vector(0 downto 0);
  signal place_693_top : bit;
  signal place_694_tip : bit_vector(0 downto 0);
  signal place_694_rst : bit_vector(0 downto 0);
  signal place_694_top : bit;
  signal place_695_tip : bit_vector(0 downto 0);
  signal place_695_rst : bit_vector(0 downto 0);
  signal place_695_top : bit;
  signal place_696_tip : bit_vector(0 downto 0);
  signal place_696_rst : bit_vector(0 downto 0);
  signal place_696_top : bit;
  signal place_697_tip : bit_vector(0 downto 0);
  signal place_697_rst : bit_vector(0 downto 0);
  signal place_697_top : bit;
  signal place_698_tip : bit_vector(0 downto 0);
  signal place_698_rst : bit_vector(1 downto 0);
  signal place_698_top : bit;
  signal place_7_tip : bit_vector(0 downto 0);
  signal place_7_rst : bit_vector(0 downto 0);
  signal place_7_top : bit;
  signal place_701_tip : bit_vector(1 downto 0);
  signal place_701_rst : bit_vector(0 downto 0);
  signal place_701_top : bit;
  signal place_702_tip : bit_vector(0 downto 0);
  signal place_702_rst : bit_vector(0 downto 0);
  signal place_702_top : bit;
  signal place_703_tip : bit_vector(0 downto 0);
  signal place_703_rst : bit_vector(0 downto 0);
  signal place_703_top : bit;
  signal place_704_tip : bit_vector(0 downto 0);
  signal place_704_rst : bit_vector(0 downto 0);
  signal place_704_top : bit;
  signal place_705_tip : bit_vector(0 downto 0);
  signal place_705_rst : bit_vector(0 downto 0);
  signal place_705_top : bit;
  signal place_706_tip : bit_vector(0 downto 0);
  signal place_706_rst : bit_vector(0 downto 0);
  signal place_706_top : bit;
  signal place_707_tip : bit_vector(0 downto 0);
  signal place_707_rst : bit_vector(0 downto 0);
  signal place_707_top : bit;
  signal place_708_tip : bit_vector(0 downto 0);
  signal place_708_rst : bit_vector(0 downto 0);
  signal place_708_top : bit;
  signal place_709_tip : bit_vector(0 downto 0);
  signal place_709_rst : bit_vector(0 downto 0);
  signal place_709_top : bit;
  signal place_710_tip : bit_vector(0 downto 0);
  signal place_710_rst : bit_vector(0 downto 0);
  signal place_710_top : bit;
  signal place_711_tip : bit_vector(0 downto 0);
  signal place_711_rst : bit_vector(0 downto 0);
  signal place_711_top : bit;
  signal place_712_tip : bit_vector(0 downto 0);
  signal place_712_rst : bit_vector(0 downto 0);
  signal place_712_top : bit;
  signal place_713_tip : bit_vector(0 downto 0);
  signal place_713_rst : bit_vector(0 downto 0);
  signal place_713_top : bit;
  signal place_714_tip : bit_vector(0 downto 0);
  signal place_714_rst : bit_vector(0 downto 0);
  signal place_714_top : bit;
  signal place_715_tip : bit_vector(0 downto 0);
  signal place_715_rst : bit_vector(0 downto 0);
  signal place_715_top : bit;
  signal place_716_tip : bit_vector(0 downto 0);
  signal place_716_rst : bit_vector(0 downto 0);
  signal place_716_top : bit;
  signal place_717_tip : bit_vector(0 downto 0);
  signal place_717_rst : bit_vector(0 downto 0);
  signal place_717_top : bit;
  signal place_718_tip : bit_vector(0 downto 0);
  signal place_718_rst : bit_vector(0 downto 0);
  signal place_718_top : bit;
  signal place_719_tip : bit_vector(0 downto 0);
  signal place_719_rst : bit_vector(0 downto 0);
  signal place_719_top : bit;
  signal place_72_tip : bit_vector(0 downto 0);
  signal place_72_rst : bit_vector(0 downto 0);
  signal place_72_top : bit;
  signal place_720_tip : bit_vector(0 downto 0);
  signal place_720_rst : bit_vector(0 downto 0);
  signal place_720_top : bit;
  signal place_721_tip : bit_vector(0 downto 0);
  signal place_721_rst : bit_vector(0 downto 0);
  signal place_721_top : bit;
  signal place_722_tip : bit_vector(0 downto 0);
  signal place_722_rst : bit_vector(0 downto 0);
  signal place_722_top : bit;
  signal place_723_tip : bit_vector(0 downto 0);
  signal place_723_rst : bit_vector(0 downto 0);
  signal place_723_top : bit;
  signal place_724_tip : bit_vector(0 downto 0);
  signal place_724_rst : bit_vector(0 downto 0);
  signal place_724_top : bit;
  signal place_725_tip : bit_vector(0 downto 0);
  signal place_725_rst : bit_vector(0 downto 0);
  signal place_725_top : bit;
  signal place_726_tip : bit_vector(0 downto 0);
  signal place_726_rst : bit_vector(0 downto 0);
  signal place_726_top : bit;
  signal place_727_tip : bit_vector(0 downto 0);
  signal place_727_rst : bit_vector(0 downto 0);
  signal place_727_top : bit;
  signal place_728_tip : bit_vector(0 downto 0);
  signal place_728_rst : bit_vector(0 downto 0);
  signal place_728_top : bit;
  signal place_729_tip : bit_vector(0 downto 0);
  signal place_729_rst : bit_vector(0 downto 0);
  signal place_729_top : bit;
  signal place_730_tip : bit_vector(0 downto 0);
  signal place_730_rst : bit_vector(0 downto 0);
  signal place_730_top : bit;
  signal place_731_tip : bit_vector(0 downto 0);
  signal place_731_rst : bit_vector(0 downto 0);
  signal place_731_top : bit;
  signal place_732_tip : bit_vector(0 downto 0);
  signal place_732_rst : bit_vector(0 downto 0);
  signal place_732_top : bit;
  signal place_733_tip : bit_vector(0 downto 0);
  signal place_733_rst : bit_vector(0 downto 0);
  signal place_733_top : bit;
  signal place_734_tip : bit_vector(0 downto 0);
  signal place_734_rst : bit_vector(0 downto 0);
  signal place_734_top : bit;
  signal place_735_tip : bit_vector(0 downto 0);
  signal place_735_rst : bit_vector(0 downto 0);
  signal place_735_top : bit;
  signal place_736_tip : bit_vector(0 downto 0);
  signal place_736_rst : bit_vector(0 downto 0);
  signal place_736_top : bit;
  signal place_737_tip : bit_vector(0 downto 0);
  signal place_737_rst : bit_vector(0 downto 0);
  signal place_737_top : bit;
  signal place_738_tip : bit_vector(0 downto 0);
  signal place_738_rst : bit_vector(1 downto 0);
  signal place_738_top : bit;
  signal place_739_tip : bit_vector(0 downto 0);
  signal place_739_rst : bit_vector(0 downto 0);
  signal place_739_top : bit;
  signal place_74_tip : bit_vector(0 downto 0);
  signal place_74_rst : bit_vector(0 downto 0);
  signal place_74_top : bit;
  signal place_740_tip : bit_vector(0 downto 0);
  signal place_740_rst : bit_vector(0 downto 0);
  signal place_740_top : bit;
  signal place_742_tip : bit_vector(0 downto 0);
  signal place_742_rst : bit_vector(0 downto 0);
  signal place_742_top : bit;
  signal place_744_tip : bit_vector(1 downto 0);
  signal place_744_rst : bit_vector(0 downto 0);
  signal place_744_top : bit;
  signal place_745_tip : bit_vector(0 downto 0);
  signal place_745_rst : bit_vector(0 downto 0);
  signal place_745_top : bit;
  signal place_746_tip : bit_vector(0 downto 0);
  signal place_746_rst : bit_vector(0 downto 0);
  signal place_746_top : bit;
  signal place_747_tip : bit_vector(0 downto 0);
  signal place_747_rst : bit_vector(0 downto 0);
  signal place_747_top : bit;
  signal place_748_tip : bit_vector(0 downto 0);
  signal place_748_rst : bit_vector(0 downto 0);
  signal place_748_top : bit;
  signal place_749_tip : bit_vector(0 downto 0);
  signal place_749_rst : bit_vector(0 downto 0);
  signal place_749_top : bit;
  signal place_75_tip : bit_vector(0 downto 0);
  signal place_75_rst : bit_vector(0 downto 0);
  signal place_75_top : bit;
  signal place_750_tip : bit_vector(0 downto 0);
  signal place_750_rst : bit_vector(0 downto 0);
  signal place_750_top : bit;
  signal place_751_tip : bit_vector(0 downto 0);
  signal place_751_rst : bit_vector(0 downto 0);
  signal place_751_top : bit;
  signal place_752_tip : bit_vector(0 downto 0);
  signal place_752_rst : bit_vector(0 downto 0);
  signal place_752_top : bit;
  signal place_753_tip : bit_vector(0 downto 0);
  signal place_753_rst : bit_vector(1 downto 0);
  signal place_753_top : bit;
  signal place_77_tip : bit_vector(0 downto 0);
  signal place_77_rst : bit_vector(0 downto 0);
  signal place_77_top : bit;
  signal place_81_tip : bit_vector(0 downto 0);
  signal place_81_rst : bit_vector(0 downto 0);
  signal place_81_top : bit;
  signal place_83_tip : bit_vector(0 downto 0);
  signal place_83_rst : bit_vector(0 downto 0);
  signal place_83_top : bit;
  signal place_84_tip : bit_vector(0 downto 0);
  signal place_84_rst : bit_vector(0 downto 0);
  signal place_84_top : bit;
  signal place_86_tip : bit_vector(0 downto 0);
  signal place_86_rst : bit_vector(0 downto 0);
  signal place_86_top : bit;
  signal place_87_tip : bit_vector(0 downto 0);
  signal place_87_rst : bit_vector(0 downto 0);
  signal place_87_top : bit;
  signal place_88_tip : bit_vector(0 downto 0);
  signal place_88_rst : bit_vector(0 downto 0);
  signal place_88_top : bit;
  signal place_89_tip : bit_vector(0 downto 0);
  signal place_89_rst : bit_vector(0 downto 0);
  signal place_89_top : bit;
  signal place_9_tip : bit_vector(0 downto 0);
  signal place_9_rst : bit_vector(0 downto 0);
  signal place_9_top : bit;
  signal place_90_tip : bit_vector(0 downto 0);
  signal place_90_rst : bit_vector(0 downto 0);
  signal place_90_top : bit;
  signal place_91_tip : bit_vector(0 downto 0);
  signal place_91_rst : bit_vector(0 downto 0);
  signal place_91_top : bit;
  signal place_92_tip : bit_vector(0 downto 0);
  signal place_92_rst : bit_vector(0 downto 0);
  signal place_92_top : bit;
  signal place_93_tip : bit_vector(0 downto 0);
  signal place_93_rst : bit_vector(0 downto 0);
  signal place_93_top : bit;
  signal place_94_tip : bit_vector(0 downto 0);
  signal place_94_rst : bit_vector(0 downto 0);
  signal place_94_top : bit;
  signal place_95_tip : bit_vector(0 downto 0);
  signal place_95_rst : bit_vector(0 downto 0);
  signal place_95_top : bit;
  signal place_96_tip : bit_vector(0 downto 0);
  signal place_96_rst : bit_vector(0 downto 0);
  signal place_96_top : bit;
  signal place_97_tip : bit_vector(0 downto 0);
  signal place_97_rst : bit_vector(0 downto 0);
  signal place_97_top : bit;
  signal place_99_tip : bit_vector(0 downto 0);
  signal place_99_rst : bit_vector(0 downto 0);
  signal place_99_top : bit;

  signal cbr_10_oper_tmp_d_42_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_10_oper_tmp_d_42_bool_d_req_ge : bit;
  signal cbr_10_oper_tmp_d_42_bool_d_req_top : bit;
  signal cbr_11_oper_tmp_d_54_bool_d_req_tip : bit_vector(2 downto 0);
  signal cbr_11_oper_tmp_d_54_bool_d_req_ge : bit;
  signal cbr_11_oper_tmp_d_54_bool_d_req_top : bit;
  signal cbr_12_oper_tmp_d_4223_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_12_oper_tmp_d_4223_bool_d_req_ge : bit;
  signal cbr_12_oper_tmp_d_4223_bool_d_req_top : bit;
  signal cbr_13_oper_exitcond128_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_13_oper_exitcond128_bool_d_req_ge : bit;
  signal cbr_13_oper_exitcond128_bool_d_req_top : bit;
  signal cbr_14_oper_exitcond131_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_14_oper_exitcond131_bool_d_req_ge : bit;
  signal cbr_14_oper_exitcond131_bool_d_req_top : bit;
  signal cbr_15_oper_tmp_d_92_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_15_oper_tmp_d_92_bool_d_req_ge : bit;
  signal cbr_15_oper_tmp_d_92_bool_d_req_top : bit;
  signal cbr_16_oper_tmp_d_11348_bool_d_req_tip : bit_vector(2 downto 0);
  signal cbr_16_oper_tmp_d_11348_bool_d_req_ge : bit;
  signal cbr_16_oper_tmp_d_11348_bool_d_req_top : bit;
  signal cbr_17_oper_tmp_d_113_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_17_oper_tmp_d_113_bool_d_req_ge : bit;
  signal cbr_17_oper_tmp_d_113_bool_d_req_top : bit;
  signal cbr_18_oper_exitcond142_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_18_oper_exitcond142_bool_d_req_ge : bit;
  signal cbr_18_oper_exitcond142_bool_d_req_top : bit;
  signal cbr_19_oper_tmp_d_149_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_19_oper_tmp_d_149_bool_d_req_ge : bit;
  signal cbr_19_oper_tmp_d_149_bool_d_req_top : bit;
  signal cbr_20_oper_tmp_d_14574_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_20_oper_tmp_d_14574_bool_d_req_ge : bit;
  signal cbr_20_oper_tmp_d_14574_bool_d_req_top : bit;
  signal cbr_21_oper_tmp_d_166_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_21_oper_tmp_d_166_bool_d_req_ge : bit;
  signal cbr_21_oper_tmp_d_166_bool_d_req_top : bit;
  signal cbr_22_oper_tmp_d_14578_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_22_oper_tmp_d_14578_bool_d_req_ge : bit;
  signal cbr_22_oper_tmp_d_14578_bool_d_req_top : bit;
  signal cbr_23_oper_tmp_d_14580_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_23_oper_tmp_d_14580_bool_d_req_ge : bit;
  signal cbr_23_oper_tmp_d_14580_bool_d_req_top : bit;
  signal cbr_24_oper_exitcond145_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_24_oper_exitcond145_bool_d_req_ge : bit;
  signal cbr_24_oper_exitcond145_bool_d_req_top : bit;
  signal cbr_25_oper_tmp_d_202_bool_d_req_tip : bit_vector(2 downto 0);
  signal cbr_25_oper_tmp_d_202_bool_d_req_ge : bit;
  signal cbr_25_oper_tmp_d_202_bool_d_req_top : bit;
  signal cbr_26_oper_tmp_d_20299_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_26_oper_tmp_d_20299_bool_d_req_ge : bit;
  signal cbr_26_oper_tmp_d_20299_bool_d_req_top : bit;
  signal cbr_27_oper_exitcond150_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_27_oper_exitcond150_bool_d_req_ge : bit;
  signal cbr_27_oper_exitcond150_bool_d_req_top : bit;
  signal cbr_28_oper_tmp_d_221_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_28_oper_tmp_d_221_bool_d_req_ge : bit;
  signal cbr_28_oper_tmp_d_221_bool_d_req_top : bit;
  signal cbr_29_oper_tmp_d_221111_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_29_oper_tmp_d_221111_bool_d_req_ge : bit;
  signal cbr_29_oper_tmp_d_221111_bool_d_req_top : bit;
  signal cbr_30_oper_exitcond158_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_30_oper_exitcond158_bool_d_req_ge : bit;
  signal cbr_30_oper_exitcond158_bool_d_req_top : bit;
  signal cbr_6_oper_exitcond_bool_d_req_tip : bit_vector(2 downto 0);
  signal cbr_6_oper_exitcond_bool_d_req_ge : bit;
  signal cbr_6_oper_exitcond_bool_d_req_top : bit;
  signal cbr_7_oper_exitcond120_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_7_oper_exitcond120_bool_d_req_ge : bit;
  signal cbr_7_oper_exitcond120_bool_d_req_top : bit;
  signal cbr_8_oper_tmp_d_16_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_8_oper_tmp_d_16_bool_d_req_ge : bit;
  signal cbr_8_oper_tmp_d_16_bool_d_req_top : bit;
  signal cbr_9_oper_tmp_d_1614_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_9_oper_tmp_d_1614_bool_d_req_ge : bit;
  signal cbr_9_oper_tmp_d_1614_bool_d_req_top : bit;
  signal else_d_0_d_entry_tip : bit_vector(0 downto 0);
  signal else_d_0_d_entry_ge : bit;
  signal else_d_0_d_entry_top : bit;
  signal else_d_0_to_else_d_1_src_tip : bit_vector(0 downto 0);
  signal else_d_0_to_else_d_1_src_ge : bit;
  signal else_d_0_to_else_d_1_src_top : bit;
  signal else_d_0_to_then_d_2_src_tip : bit_vector(0 downto 0);
  signal else_d_0_to_then_d_2_src_ge : bit;
  signal else_d_0_to_then_d_2_src_top : bit;
  signal else_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal else_d_1_d_entry_ge : bit;
  signal else_d_1_d_entry_top : bit;
  signal else_d_1_to_loopexit_d_10_src_tip : bit_vector(0 downto 0);
  signal else_d_1_to_loopexit_d_10_src_ge : bit;
  signal else_d_1_to_loopexit_d_10_src_top : bit;
  signal else_d_1_to_no_exit_d_10_d_backedge_src_tip : bit_vector(0 downto 0);
  signal else_d_1_to_no_exit_d_10_d_backedge_src_ge : bit;
  signal else_d_1_to_no_exit_d_10_d_backedge_src_top : bit;
  signal fin_tip : bit_vector(0 downto 0);
  signal fin_ge : bit;
  signal fin_top : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar118_d_ph_d_ph_mux_1_d_ack_ge : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_ack_top : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar118_d_ph_d_ph_mux_1_d_req0_ge : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_req0_top : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar118_d_ph_d_ph_mux_1_d_req1_ge : bit;
  signal indvar118_d_ph_d_ph_mux_1_d_req1_top : bit;
  signal indvar121_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar121_mux_1_d_ack_ge : bit;
  signal indvar121_mux_1_d_ack_top : bit;
  signal indvar121_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar121_mux_1_d_req0_ge : bit;
  signal indvar121_mux_1_d_req0_top : bit;
  signal indvar121_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar121_mux_1_d_req1_ge : bit;
  signal indvar121_mux_1_d_req1_top : bit;
  signal indvar123_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar123_mux_1_d_ack_ge : bit;
  signal indvar123_mux_1_d_ack_top : bit;
  signal indvar123_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar123_mux_1_d_req0_ge : bit;
  signal indvar123_mux_1_d_req0_top : bit;
  signal indvar123_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar123_mux_1_d_req1_ge : bit;
  signal indvar123_mux_1_d_req1_top : bit;
  signal indvar126_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar126_mux_1_d_ack_ge : bit;
  signal indvar126_mux_1_d_ack_top : bit;
  signal indvar126_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar126_mux_1_d_req0_ge : bit;
  signal indvar126_mux_1_d_req0_top : bit;
  signal indvar126_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar126_mux_1_d_req1_ge : bit;
  signal indvar126_mux_1_d_req1_top : bit;
  signal indvar129_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar129_mux_1_d_ack_ge : bit;
  signal indvar129_mux_1_d_ack_top : bit;
  signal indvar129_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar129_mux_1_d_req0_ge : bit;
  signal indvar129_mux_1_d_req0_top : bit;
  signal indvar129_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar129_mux_1_d_req1_ge : bit;
  signal indvar129_mux_1_d_req1_top : bit;
  signal indvar132_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar132_mux_1_d_ack_ge : bit;
  signal indvar132_mux_1_d_ack_top : bit;
  signal indvar132_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar132_mux_1_d_req0_ge : bit;
  signal indvar132_mux_1_d_req0_top : bit;
  signal indvar132_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar132_mux_1_d_req1_ge : bit;
  signal indvar132_mux_1_d_req1_top : bit;
  signal indvar134_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar134_mux_1_d_ack_ge : bit;
  signal indvar134_mux_1_d_ack_top : bit;
  signal indvar134_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar134_mux_1_d_req0_ge : bit;
  signal indvar134_mux_1_d_req0_top : bit;
  signal indvar134_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar134_mux_1_d_req1_ge : bit;
  signal indvar134_mux_1_d_req1_top : bit;
  signal indvar138_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar138_mux_1_d_ack_ge : bit;
  signal indvar138_mux_1_d_ack_top : bit;
  signal indvar138_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar138_mux_1_d_req0_ge : bit;
  signal indvar138_mux_1_d_req0_top : bit;
  signal indvar138_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar138_mux_1_d_req1_ge : bit;
  signal indvar138_mux_1_d_req1_top : bit;
  signal indvar143_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar143_mux_1_d_ack_ge : bit;
  signal indvar143_mux_1_d_ack_top : bit;
  signal indvar143_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar143_mux_1_d_req0_ge : bit;
  signal indvar143_mux_1_d_req0_top : bit;
  signal indvar143_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar143_mux_1_d_req1_ge : bit;
  signal indvar143_mux_1_d_req1_top : bit;
  signal indvar146_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar146_mux_1_d_ack_ge : bit;
  signal indvar146_mux_1_d_ack_top : bit;
  signal indvar146_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar146_mux_1_d_req0_ge : bit;
  signal indvar146_mux_1_d_req0_top : bit;
  signal indvar146_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar146_mux_1_d_req1_ge : bit;
  signal indvar146_mux_1_d_req1_top : bit;
  signal indvar148_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar148_mux_1_d_ack_ge : bit;
  signal indvar148_mux_1_d_ack_top : bit;
  signal indvar148_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar148_mux_1_d_req0_ge : bit;
  signal indvar148_mux_1_d_req0_top : bit;
  signal indvar148_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar148_mux_1_d_req1_ge : bit;
  signal indvar148_mux_1_d_req1_top : bit;
  signal indvar151_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar151_mux_1_d_ack_ge : bit;
  signal indvar151_mux_1_d_ack_top : bit;
  signal indvar151_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar151_mux_1_d_req0_ge : bit;
  signal indvar151_mux_1_d_req0_top : bit;
  signal indvar151_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar151_mux_1_d_req1_ge : bit;
  signal indvar151_mux_1_d_req1_top : bit;
  signal indvar153_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar153_mux_1_d_ack_ge : bit;
  signal indvar153_mux_1_d_ack_top : bit;
  signal indvar153_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar153_mux_1_d_req0_ge : bit;
  signal indvar153_mux_1_d_req0_top : bit;
  signal indvar153_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar153_mux_1_d_req1_ge : bit;
  signal indvar153_mux_1_d_req1_top : bit;
  signal indvar_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal indvar_mux_1_d_ack_ge : bit;
  signal indvar_mux_1_d_ack_top : bit;
  signal indvar_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal indvar_mux_1_d_req0_ge : bit;
  signal indvar_mux_1_d_req0_top : bit;
  signal indvar_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal indvar_mux_1_d_req1_ge : bit;
  signal indvar_mux_1_d_req1_top : bit;
  signal init_tip : bit_vector(0 downto 0);
  signal init_ge : bit;
  signal init_top : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_d_ph_mux_1_d_ack_ge : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_ack_top : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_d_ph_mux_1_d_req0_ge : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_req0_top : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_d_ph_mux_1_d_req1_ge : bit;
  signal j_d_3_d_in_d_ph_mux_1_d_req1_top : bit;
  signal j_d_3_d_in_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_mux_1_d_ack_ge : bit;
  signal j_d_3_d_in_mux_1_d_ack_top : bit;
  signal j_d_3_d_in_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_mux_1_d_req0_ge : bit;
  signal j_d_3_d_in_mux_1_d_req0_top : bit;
  signal j_d_3_d_in_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal j_d_3_d_in_mux_1_d_req1_ge : bit;
  signal j_d_3_d_in_mux_1_d_req1_top : bit;
  signal j_d_9_d_2_d_be_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_1_d_ack_ge : bit;
  signal j_d_9_d_2_d_be_mux_1_d_ack_top : bit;
  signal j_d_9_d_2_d_be_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_1_d_req0_ge : bit;
  signal j_d_9_d_2_d_be_mux_1_d_req0_top : bit;
  signal j_d_9_d_2_d_be_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_1_d_req1_ge : bit;
  signal j_d_9_d_2_d_be_mux_1_d_req1_top : bit;
  signal j_d_9_d_2_d_be_mux_2_d_ack_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_2_d_ack_ge : bit;
  signal j_d_9_d_2_d_be_mux_2_d_ack_top : bit;
  signal j_d_9_d_2_d_be_mux_2_d_req0_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_2_d_req0_ge : bit;
  signal j_d_9_d_2_d_be_mux_2_d_req0_top : bit;
  signal j_d_9_d_2_d_be_mux_2_d_req1_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_d_be_mux_2_d_req1_ge : bit;
  signal j_d_9_d_2_d_be_mux_2_d_req1_top : bit;
  signal j_d_9_d_2_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_mux_1_d_ack_ge : bit;
  signal j_d_9_d_2_mux_1_d_ack_top : bit;
  signal j_d_9_d_2_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_mux_1_d_req0_ge : bit;
  signal j_d_9_d_2_mux_1_d_req0_top : bit;
  signal j_d_9_d_2_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal j_d_9_d_2_mux_1_d_req1_ge : bit;
  signal j_d_9_d_2_mux_1_d_req1_top : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal k_d_1_d_in_d_ph_mux_1_d_ack_ge : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_ack_top : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal k_d_1_d_in_d_ph_mux_1_d_req0_ge : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_req0_top : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal k_d_1_d_in_d_ph_mux_1_d_req1_ge : bit;
  signal k_d_1_d_in_d_ph_mux_1_d_req1_top : bit;
  signal k_d_2_d_3_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal k_d_2_d_3_mux_1_d_ack_ge : bit;
  signal k_d_2_d_3_mux_1_d_ack_top : bit;
  signal k_d_2_d_3_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal k_d_2_d_3_mux_1_d_req0_ge : bit;
  signal k_d_2_d_3_mux_1_d_req0_top : bit;
  signal k_d_2_d_3_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal k_d_2_d_3_mux_1_d_req1_ge : bit;
  signal k_d_2_d_3_mux_1_d_req1_top : bit;
  signal k_d_3_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal k_d_3_d_0_mux_1_d_ack_ge : bit;
  signal k_d_3_d_0_mux_1_d_ack_top : bit;
  signal k_d_3_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal k_d_3_d_0_mux_1_d_req0_ge : bit;
  signal k_d_3_d_0_mux_1_d_req0_top : bit;
  signal k_d_3_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal k_d_3_d_0_mux_1_d_req1_ge : bit;
  signal k_d_3_d_0_mux_1_d_req1_top : bit;
  signal k_d_4_d_3_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal k_d_4_d_3_mux_1_d_ack_ge : bit;
  signal k_d_4_d_3_mux_1_d_ack_top : bit;
  signal k_d_4_d_3_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal k_d_4_d_3_mux_1_d_req0_ge : bit;
  signal k_d_4_d_3_mux_1_d_req0_top : bit;
  signal k_d_4_d_3_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal k_d_4_d_3_mux_1_d_req1_ge : bit;
  signal k_d_4_d_3_mux_1_d_req1_top : bit;
  signal k_d_5_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal k_d_5_d_0_mux_1_d_ack_ge : bit;
  signal k_d_5_d_0_mux_1_d_ack_top : bit;
  signal k_d_5_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal k_d_5_d_0_mux_1_d_req0_ge : bit;
  signal k_d_5_d_0_mux_1_d_req0_top : bit;
  signal k_d_5_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal k_d_5_d_0_mux_1_d_req1_ge : bit;
  signal k_d_5_d_0_mux_1_d_req1_top : bit;
  signal load_A_d_ack_tip : bit_vector(0 downto 0);
  signal load_A_d_ack_ge : bit;
  signal load_A_d_ack_top : bit;
  signal load_A_d_req_tip : bit_vector(0 downto 0);
  signal load_A_d_req_ge : bit;
  signal load_A_d_req_top : bit;
  signal load_ccoeff_d_ack_tip : bit_vector(0 downto 0);
  signal load_ccoeff_d_ack_ge : bit;
  signal load_ccoeff_d_ack_top : bit;
  signal load_ccoeff_d_req_tip : bit_vector(0 downto 0);
  signal load_ccoeff_d_req_ge : bit;
  signal load_ccoeff_d_req_top : bit;
  signal load_l_array_d_ack_tip : bit_vector(0 downto 0);
  signal load_l_array_d_ack_ge : bit;
  signal load_l_array_d_ack_top : bit;
  signal load_l_array_d_req_tip : bit_vector(0 downto 0);
  signal load_l_array_d_req_ge : bit;
  signal load_l_array_d_req_top : bit;
  signal load_noofelem_d_ack_tip : bit_vector(0 downto 0);
  signal load_noofelem_d_ack_ge : bit;
  signal load_noofelem_d_ack_top : bit;
  signal load_noofelem_d_req_tip : bit_vector(0 downto 0);
  signal load_noofelem_d_req_ge : bit;
  signal load_noofelem_d_req_top : bit;
  signal load_rcoeff_d_ack_tip : bit_vector(0 downto 0);
  signal load_rcoeff_d_ack_ge : bit;
  signal load_rcoeff_d_ack_top : bit;
  signal load_rcoeff_d_req_tip : bit_vector(0 downto 0);
  signal load_rcoeff_d_req_ge : bit;
  signal load_rcoeff_d_req_top : bit;
  signal load_start_call_divide_0_return_d_ack_tip : bit_vector(0 downto 0);
  signal load_start_call_divide_0_return_d_ack_ge : bit;
  signal load_start_call_divide_0_return_d_ack_top : bit;
  signal load_start_call_divide_0_return_d_req_tip : bit_vector(0 downto 0);
  signal load_start_call_divide_0_return_d_req_ge : bit;
  signal load_start_call_divide_0_return_d_req_top : bit;
  signal load_tmp_d_103_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_103_d_ack_ge : bit;
  signal load_tmp_d_103_d_ack_top : bit;
  signal load_tmp_d_103_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_103_d_req_ge : bit;
  signal load_tmp_d_103_d_req_top : bit;
  signal load_tmp_d_108_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_108_d_ack_ge : bit;
  signal load_tmp_d_108_d_ack_top : bit;
  signal load_tmp_d_108_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_108_d_req_ge : bit;
  signal load_tmp_d_108_d_req_top : bit;
  signal load_tmp_d_123_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_123_d_ack_ge : bit;
  signal load_tmp_d_123_d_ack_top : bit;
  signal load_tmp_d_123_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_123_d_req_ge : bit;
  signal load_tmp_d_123_d_req_top : bit;
  signal load_tmp_d_128_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_128_d_ack_ge : bit;
  signal load_tmp_d_128_d_ack_top : bit;
  signal load_tmp_d_128_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_128_d_req_ge : bit;
  signal load_tmp_d_128_d_req_top : bit;
  signal load_tmp_d_133_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_133_d_ack_ge : bit;
  signal load_tmp_d_133_d_ack_top : bit;
  signal load_tmp_d_133_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_133_d_req_ge : bit;
  signal load_tmp_d_133_d_req_top : bit;
  signal load_tmp_d_159_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_159_d_ack_ge : bit;
  signal load_tmp_d_159_d_ack_top : bit;
  signal load_tmp_d_159_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_159_d_req_ge : bit;
  signal load_tmp_d_159_d_req_top : bit;
  signal load_tmp_d_180_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_180_d_ack_ge : bit;
  signal load_tmp_d_180_d_ack_top : bit;
  signal load_tmp_d_180_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_180_d_req_ge : bit;
  signal load_tmp_d_180_d_req_top : bit;
  signal load_tmp_d_193_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_193_d_ack_ge : bit;
  signal load_tmp_d_193_d_ack_top : bit;
  signal load_tmp_d_193_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_193_d_req_ge : bit;
  signal load_tmp_d_193_d_req_top : bit;
  signal load_tmp_d_211_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_211_d_ack_ge : bit;
  signal load_tmp_d_211_d_ack_top : bit;
  signal load_tmp_d_211_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_211_d_req_ge : bit;
  signal load_tmp_d_211_d_req_top : bit;
  signal load_tmp_d_21_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_21_d_ack_ge : bit;
  signal load_tmp_d_21_d_ack_top : bit;
  signal load_tmp_d_21_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_21_d_req_ge : bit;
  signal load_tmp_d_21_d_req_top : bit;
  signal load_tmp_d_230_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_230_d_ack_ge : bit;
  signal load_tmp_d_230_d_ack_top : bit;
  signal load_tmp_d_230_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_230_d_req_ge : bit;
  signal load_tmp_d_230_d_req_top : bit;
  signal load_tmp_d_26_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_26_d_ack_ge : bit;
  signal load_tmp_d_26_d_ack_top : bit;
  signal load_tmp_d_26_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_26_d_req_ge : bit;
  signal load_tmp_d_26_d_req_top : bit;
  signal load_tmp_d_31_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_31_d_ack_ge : bit;
  signal load_tmp_d_31_d_ack_top : bit;
  signal load_tmp_d_31_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_31_d_req_ge : bit;
  signal load_tmp_d_31_d_req_top : bit;
  signal load_tmp_d_48_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_48_d_ack_ge : bit;
  signal load_tmp_d_48_d_ack_top : bit;
  signal load_tmp_d_48_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_48_d_req_ge : bit;
  signal load_tmp_d_48_d_req_top : bit;
  signal load_tmp_d_53_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_53_d_ack_ge : bit;
  signal load_tmp_d_53_d_ack_top : bit;
  signal load_tmp_d_53_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_53_d_req_ge : bit;
  signal load_tmp_d_53_d_req_top : bit;
  signal load_tmp_d_66_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_66_d_ack_ge : bit;
  signal load_tmp_d_66_d_ack_top : bit;
  signal load_tmp_d_66_d_req_tip : bit_vector(0 downto 0);
  signal load_tmp_d_66_d_req_ge : bit;
  signal load_tmp_d_66_d_req_top : bit;
  signal load_tmp_d_75_d_ack_tip : bit_vector(0 downto 0);
  signal load_tmp_d_75_d_ack_ge : bit;
  signal load_tmp_d_75_d_ack_top : bit;
  signal load_tmp_d_75_d_req_tip : bit_vector(1 downto 0);
  signal load_tmp_d_75_d_req_ge : bit;
  signal load_tmp_d_75_d_req_top : bit;
  signal load_u_array_d_ack_tip : bit_vector(0 downto 0);
  signal load_u_array_d_ack_ge : bit;
  signal load_u_array_d_ack_top : bit;
  signal load_u_array_d_req_tip : bit_vector(0 downto 0);
  signal load_u_array_d_req_ge : bit;
  signal load_u_array_d_req_top : bit;
  signal loopentry_d_12_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_12_d_entry_ge : bit;
  signal loopentry_d_12_d_entry_top : bit;
  signal loopentry_d_12_d_loopexit_to_loopentry_d_12_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_12_d_loopexit_to_loopentry_d_12_src_ge : bit;
  signal loopentry_d_12_d_loopexit_to_loopentry_d_12_src_top : bit;
  signal loopentry_d_12_d_pre_tip : bit_vector(1 downto 0);
  signal loopentry_d_12_d_pre_ge : bit;
  signal loopentry_d_12_d_pre_top : bit;
  signal loopentry_d_12_to_loopexit_d_12_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_12_to_loopexit_d_12_src_ge : bit;
  signal loopentry_d_12_to_loopexit_d_12_src_top : bit;
  signal loopentry_d_12_to_no_exit_d_12_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_12_to_no_exit_d_12_d_preheader_src_ge : bit;
  signal loopentry_d_12_to_no_exit_d_12_d_preheader_src_top : bit;
  signal loopentry_d_14_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_14_d_entry_ge : bit;
  signal loopentry_d_14_d_entry_top : bit;
  signal loopentry_d_14_d_loopexit_to_loopentry_d_14_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_14_d_loopexit_to_loopentry_d_14_src_ge : bit;
  signal loopentry_d_14_d_loopexit_to_loopentry_d_14_src_top : bit;
  signal loopentry_d_14_d_pre_tip : bit_vector(1 downto 0);
  signal loopentry_d_14_d_pre_ge : bit;
  signal loopentry_d_14_d_pre_top : bit;
  signal loopentry_d_14_to_loopexit_d_14_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_14_to_loopexit_d_14_src_ge : bit;
  signal loopentry_d_14_to_loopexit_d_14_src_top : bit;
  signal loopentry_d_14_to_no_exit_d_14_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_14_to_no_exit_d_14_d_preheader_src_ge : bit;
  signal loopentry_d_14_to_no_exit_d_14_d_preheader_src_top : bit;
  signal loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_ge : bit;
  signal loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_top : bit;
  signal loopentry_d_2_to_no_exit_d_2_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_2_to_no_exit_d_2_d_preheader_src_ge : bit;
  signal loopentry_d_2_to_no_exit_d_2_d_preheader_src_top : bit;
  signal loopentry_d_4_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_d_entry_ge : bit;
  signal loopentry_d_4_d_entry_top : bit;
  signal loopentry_d_4_d_loopexit_to_loopentry_d_4_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_d_loopexit_to_loopentry_d_4_src_ge : bit;
  signal loopentry_d_4_d_loopexit_to_loopentry_d_4_src_top : bit;
  signal loopentry_d_4_d_outer_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_d_outer_d_entry_ge : bit;
  signal loopentry_d_4_d_outer_d_entry_top : bit;
  signal loopentry_d_4_d_outer_d_pre_tip : bit_vector(2 downto 0);
  signal loopentry_d_4_d_outer_d_pre_ge : bit;
  signal loopentry_d_4_d_outer_d_pre_top : bit;
  signal loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_ge : bit;
  signal loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top : bit;
  signal loopentry_d_4_d_outer_to_loopentry_d_4_src_tip : bit_vector(3 downto 0);
  signal loopentry_d_4_d_outer_to_loopentry_d_4_src_ge : bit;
  signal loopentry_d_4_d_outer_to_loopentry_d_4_src_top : bit;
  signal loopentry_d_4_d_pre_tip : bit_vector(1 downto 0);
  signal loopentry_d_4_d_pre_ge : bit;
  signal loopentry_d_4_d_pre_top : bit;
  signal loopentry_d_4_to_no_exit_d_4_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_to_no_exit_d_4_d_preheader_src_ge : bit;
  signal loopentry_d_4_to_no_exit_d_4_d_preheader_src_top : bit;
  signal loopentry_d_4_to_no_exit_d_5_d_preheader_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_4_to_no_exit_d_5_d_preheader_src_ge : bit;
  signal loopentry_d_4_to_no_exit_d_5_d_preheader_src_top : bit;
  signal loopentry_d_7_d_outer_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_7_d_outer_d_entry_ge : bit;
  signal loopentry_d_7_d_outer_d_entry_top : bit;
  signal loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_ge : bit;
  signal loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_top : bit;
  signal loopentry_d_7_d_outer_d_pre_tip : bit_vector(1 downto 0);
  signal loopentry_d_7_d_outer_d_pre_ge : bit;
  signal loopentry_d_7_d_outer_d_pre_top : bit;
  signal loopentry_d_7_d_outer_to_loopentry_d_7_src_tip : bit_vector(3 downto 0);
  signal loopentry_d_7_d_outer_to_loopentry_d_7_src_ge : bit;
  signal loopentry_d_7_d_outer_to_loopentry_d_7_src_top : bit;
  signal loopentry_d_7_to_loopexit_d_7_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_7_to_loopexit_d_7_src_ge : bit;
  signal loopentry_d_7_to_loopexit_d_7_src_top : bit;
  signal loopentry_d_7_to_no_exit_d_7_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_7_to_no_exit_d_7_src_ge : bit;
  signal loopentry_d_7_to_no_exit_d_7_src_top : bit;
  signal loopexit_d_10_to_loopentry_d_12_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_10_to_loopentry_d_12_d_loopexit_src_ge : bit;
  signal loopexit_d_10_to_loopentry_d_12_d_loopexit_src_top : bit;
  signal loopexit_d_10_to_no_exit_d_10_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_10_to_no_exit_d_10_d_outer_src_ge : bit;
  signal loopexit_d_10_to_no_exit_d_10_d_outer_src_top : bit;
  signal loopexit_d_12_d_entry_tip : bit_vector(0 downto 0);
  signal loopexit_d_12_d_entry_ge : bit;
  signal loopexit_d_12_d_entry_top : bit;
  signal loopexit_d_12_to_loopentry_d_12_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_12_to_loopentry_d_12_src_ge : bit;
  signal loopexit_d_12_to_loopentry_d_12_src_top : bit;
  signal loopexit_d_12_to_loopentry_d_14_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_12_to_loopentry_d_14_d_loopexit_src_ge : bit;
  signal loopexit_d_12_to_loopentry_d_14_d_loopexit_src_top : bit;
  signal loopexit_d_14_d_entry_tip : bit_vector(0 downto 0);
  signal loopexit_d_14_d_entry_ge : bit;
  signal loopexit_d_14_d_entry_top : bit;
  signal loopexit_d_14_to_loopentry_d_14_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_14_to_loopentry_d_14_src_ge : bit;
  signal loopexit_d_14_to_loopentry_d_14_src_top : bit;
  signal loopexit_d_14_to_return_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_14_to_return_src_ge : bit;
  signal loopexit_d_14_to_return_src_top : bit;
  signal loopexit_d_1_to_loopentry_d_2_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_to_loopentry_d_2_src_ge : bit;
  signal loopexit_d_1_to_loopentry_d_2_src_top : bit;
  signal loopexit_d_1_to_no_exit_d_1_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_1_to_no_exit_d_1_d_outer_src_ge : bit;
  signal loopexit_d_1_to_no_exit_d_1_d_outer_src_top : bit;
  signal loopexit_d_5_d_entry_tip : bit_vector(0 downto 0);
  signal loopexit_d_5_d_entry_ge : bit;
  signal loopexit_d_5_d_entry_top : bit;
  signal loopexit_d_5_to_loopentry_d_4_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_5_to_loopentry_d_4_d_outer_src_ge : bit;
  signal loopexit_d_5_to_loopentry_d_4_d_outer_src_top : bit;
  signal loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_ge : bit;
  signal loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_top : bit;
  signal loopexit_d_7_to_loopentry_d_7_d_outer_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_7_to_loopentry_d_7_d_outer_src_ge : bit;
  signal loopexit_d_7_to_loopentry_d_7_d_outer_src_top : bit;
  signal loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_ge : bit;
  signal loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_top : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_2_mux_1_d_ack_ge : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_ack_top : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_2_mux_1_d_req0_ge : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_req0_top : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_2_mux_1_d_req1_ge : bit;
  signal maxcoeff_d_2_d_2_mux_1_d_req1_top : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_ge : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_top : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_ge : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_top : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_ge : bit;
  signal maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_top : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_ph_mux_1_d_ack_ge : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_ack_top : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_ph_mux_1_d_req0_ge : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_req0_top : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_d_ph_mux_1_d_req1_ge : bit;
  signal maxcoeff_d_2_d_ph_mux_1_d_req1_top : bit;
  signal maxcoeff_d_2_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_mux_1_d_ack_ge : bit;
  signal maxcoeff_d_2_mux_1_d_ack_top : bit;
  signal maxcoeff_d_2_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_mux_1_d_req0_ge : bit;
  signal maxcoeff_d_2_mux_1_d_req0_top : bit;
  signal maxcoeff_d_2_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal maxcoeff_d_2_mux_1_d_req1_ge : bit;
  signal maxcoeff_d_2_mux_1_d_req1_top : bit;
  signal no_exit_d_10_to_else_d_0_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_10_to_else_d_0_src_ge : bit;
  signal no_exit_d_10_to_else_d_0_src_top : bit;
  signal no_exit_d_10_to_then_d_1_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_10_to_then_d_1_src_ge : bit;
  signal no_exit_d_10_to_then_d_1_src_top : bit;
  signal no_exit_d_12_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_12_d_entry_ge : bit;
  signal no_exit_d_12_d_entry_top : bit;
  signal no_exit_d_12_to_loopexit_d_12_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_12_to_loopexit_d_12_d_loopexit_src_ge : bit;
  signal no_exit_d_12_to_loopexit_d_12_d_loopexit_src_top : bit;
  signal no_exit_d_12_to_no_exit_d_12_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_12_to_no_exit_d_12_src_ge : bit;
  signal no_exit_d_12_to_no_exit_d_12_src_top : bit;
  signal no_exit_d_14_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_14_d_entry_ge : bit;
  signal no_exit_d_14_d_entry_top : bit;
  signal no_exit_d_14_to_loopexit_d_14_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_14_to_loopexit_d_14_d_loopexit_src_ge : bit;
  signal no_exit_d_14_to_loopexit_d_14_d_loopexit_src_top : bit;
  signal no_exit_d_14_to_no_exit_d_14_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_14_to_no_exit_d_14_src_ge : bit;
  signal no_exit_d_14_to_no_exit_d_14_src_top : bit;
  signal no_exit_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_d_entry_ge : bit;
  signal no_exit_d_1_d_entry_top : bit;
  signal no_exit_d_1_to_loopexit_d_1_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_to_loopexit_d_1_src_ge : bit;
  signal no_exit_d_1_to_loopexit_d_1_src_top : bit;
  signal no_exit_d_1_to_no_exit_d_1_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_1_to_no_exit_d_1_src_ge : bit;
  signal no_exit_d_1_to_no_exit_d_1_src_top : bit;
  signal no_exit_d_2_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_d_entry_ge : bit;
  signal no_exit_d_2_d_entry_top : bit;
  signal no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_ge : bit;
  signal no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_top : bit;
  signal no_exit_d_2_to_no_exit_d_2_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_2_to_no_exit_d_2_src_ge : bit;
  signal no_exit_d_2_to_no_exit_d_2_src_top : bit;
  signal no_exit_d_4_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_4_d_entry_ge : bit;
  signal no_exit_d_4_d_entry_top : bit;
  signal no_exit_d_4_d_pre_tip : bit_vector(1 downto 0);
  signal no_exit_d_4_d_pre_ge : bit;
  signal no_exit_d_4_d_pre_top : bit;
  signal no_exit_d_4_d_preheader_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_4_d_preheader_d_entry_ge : bit;
  signal no_exit_d_4_d_preheader_d_entry_top : bit;
  signal no_exit_d_4_d_preheader_to_no_exit_d_4_src_tip : bit_vector(1 downto 0);
  signal no_exit_d_4_d_preheader_to_no_exit_d_4_src_ge : bit;
  signal no_exit_d_4_d_preheader_to_no_exit_d_4_src_top : bit;
  signal no_exit_d_4_to_loopentry_d_4_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_4_to_loopentry_d_4_d_loopexit_src_ge : bit;
  signal no_exit_d_4_to_loopentry_d_4_d_loopexit_src_top : bit;
  signal no_exit_d_4_to_then_d_0_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_4_to_then_d_0_src_ge : bit;
  signal no_exit_d_4_to_then_d_0_src_top : bit;
  signal no_exit_d_5_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_5_d_entry_ge : bit;
  signal no_exit_d_5_d_entry_top : bit;
  signal no_exit_d_5_to_loopexit_d_5_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_5_to_loopexit_d_5_src_ge : bit;
  signal no_exit_d_5_to_loopexit_d_5_src_top : bit;
  signal no_exit_d_5_to_no_exit_d_5_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_5_to_no_exit_d_5_src_ge : bit;
  signal no_exit_d_5_to_no_exit_d_5_src_top : bit;
  signal no_exit_d_7_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_7_d_entry_ge : bit;
  signal no_exit_d_7_d_entry_top : bit;
  signal no_exit_d_7_to_loopentry_d_7_d_backedge_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_7_to_loopentry_d_7_d_backedge_src_ge : bit;
  signal no_exit_d_7_to_loopentry_d_7_d_backedge_src_top : bit;
  signal no_exit_d_7_to_no_exit_d_8_d_preheader_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_7_to_no_exit_d_8_d_preheader_src_ge : bit;
  signal no_exit_d_7_to_no_exit_d_8_d_preheader_src_top : bit;
  signal no_exit_d_8_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_8_d_entry_ge : bit;
  signal no_exit_d_8_d_entry_top : bit;
  signal no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_ge : bit;
  signal no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_top : bit;
  signal no_exit_d_8_to_no_exit_d_8_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_8_to_no_exit_d_8_src_ge : bit;
  signal no_exit_d_8_to_no_exit_d_8_src_top : bit;
  signal oper_exitcond120_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond120_bool_d_ack_ge : bit;
  signal oper_exitcond120_bool_d_ack_top : bit;
  signal oper_exitcond120_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond120_bool_d_req_ge : bit;
  signal oper_exitcond120_bool_d_req_top : bit;
  signal oper_exitcond128_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond128_bool_d_ack_ge : bit;
  signal oper_exitcond128_bool_d_ack_top : bit;
  signal oper_exitcond128_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond128_bool_d_req_ge : bit;
  signal oper_exitcond128_bool_d_req_top : bit;
  signal oper_exitcond131_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond131_bool_d_ack_ge : bit;
  signal oper_exitcond131_bool_d_ack_top : bit;
  signal oper_exitcond131_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond131_bool_d_req_ge : bit;
  signal oper_exitcond131_bool_d_req_top : bit;
  signal oper_exitcond142_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond142_bool_d_ack_ge : bit;
  signal oper_exitcond142_bool_d_ack_top : bit;
  signal oper_exitcond142_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond142_bool_d_req_ge : bit;
  signal oper_exitcond142_bool_d_req_top : bit;
  signal oper_exitcond145_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond145_bool_d_ack_ge : bit;
  signal oper_exitcond145_bool_d_ack_top : bit;
  signal oper_exitcond145_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond145_bool_d_req_ge : bit;
  signal oper_exitcond145_bool_d_req_top : bit;
  signal oper_exitcond150_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond150_bool_d_ack_ge : bit;
  signal oper_exitcond150_bool_d_ack_top : bit;
  signal oper_exitcond150_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond150_bool_d_req_ge : bit;
  signal oper_exitcond150_bool_d_req_top : bit;
  signal oper_exitcond158_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond158_bool_d_ack_ge : bit;
  signal oper_exitcond158_bool_d_ack_top : bit;
  signal oper_exitcond158_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond158_bool_d_req_ge : bit;
  signal oper_exitcond158_bool_d_req_top : bit;
  signal oper_exitcond_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_exitcond_bool_d_ack_ge : bit;
  signal oper_exitcond_bool_d_ack_top : bit;
  signal oper_exitcond_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_exitcond_bool_d_req_ge : bit;
  signal oper_exitcond_bool_d_req_top : bit;
  signal oper_inc_d_11_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_11_int_d_ack_ge : bit;
  signal oper_inc_d_11_int_d_ack_top : bit;
  signal oper_inc_d_11_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_11_int_d_req_ge : bit;
  signal oper_inc_d_11_int_d_req_top : bit;
  signal oper_inc_d_12_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_12_int_d_ack_ge : bit;
  signal oper_inc_d_12_int_d_ack_top : bit;
  signal oper_inc_d_12_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_12_int_d_req_ge : bit;
  signal oper_inc_d_12_int_d_req_top : bit;
  signal oper_inc_d_14_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_14_int_d_ack_ge : bit;
  signal oper_inc_d_14_int_d_ack_top : bit;
  signal oper_inc_d_14_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_14_int_d_req_ge : bit;
  signal oper_inc_d_14_int_d_req_top : bit;
  signal oper_inc_d_15_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_15_int_d_ack_ge : bit;
  signal oper_inc_d_15_int_d_ack_top : bit;
  signal oper_inc_d_15_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_15_int_d_req_ge : bit;
  signal oper_inc_d_15_int_d_req_top : bit;
  signal oper_inc_d_2_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_2_int_d_ack_ge : bit;
  signal oper_inc_d_2_int_d_ack_top : bit;
  signal oper_inc_d_2_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_2_int_d_req_ge : bit;
  signal oper_inc_d_2_int_d_req_top : bit;
  signal oper_inc_d_5_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_5_int_d_ack_ge : bit;
  signal oper_inc_d_5_int_d_ack_top : bit;
  signal oper_inc_d_5_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_5_int_d_req_ge : bit;
  signal oper_inc_d_5_int_d_req_top : bit;
  signal oper_inc_d_960_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_960_int_d_ack_ge : bit;
  signal oper_inc_d_960_int_d_ack_top : bit;
  signal oper_inc_d_960_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_960_int_d_req_ge : bit;
  signal oper_inc_d_960_int_d_req_top : bit;
  signal oper_inc_d_976_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_976_int_d_ack_ge : bit;
  signal oper_inc_d_976_int_d_ack_top : bit;
  signal oper_inc_d_976_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_976_int_d_req_ge : bit;
  signal oper_inc_d_976_int_d_req_top : bit;
  signal oper_inc_d_9_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_9_int_d_ack_ge : bit;
  signal oper_inc_d_9_int_d_ack_top : bit;
  signal oper_inc_d_9_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_9_int_d_req_ge : bit;
  signal oper_inc_d_9_int_d_req_top : bit;
  signal oper_indvar_d_next119_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next119_uint_d_ack_ge : bit;
  signal oper_indvar_d_next119_uint_d_ack_top : bit;
  signal oper_indvar_d_next119_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next119_uint_d_req_ge : bit;
  signal oper_indvar_d_next119_uint_d_req_top : bit;
  signal oper_indvar_d_next122_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next122_uint_d_ack_ge : bit;
  signal oper_indvar_d_next122_uint_d_ack_top : bit;
  signal oper_indvar_d_next122_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next122_uint_d_req_ge : bit;
  signal oper_indvar_d_next122_uint_d_req_top : bit;
  signal oper_indvar_d_next124_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next124_uint_d_ack_ge : bit;
  signal oper_indvar_d_next124_uint_d_ack_top : bit;
  signal oper_indvar_d_next124_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next124_uint_d_req_ge : bit;
  signal oper_indvar_d_next124_uint_d_req_top : bit;
  signal oper_indvar_d_next127_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next127_uint_d_ack_ge : bit;
  signal oper_indvar_d_next127_uint_d_ack_top : bit;
  signal oper_indvar_d_next127_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next127_uint_d_req_ge : bit;
  signal oper_indvar_d_next127_uint_d_req_top : bit;
  signal oper_indvar_d_next130_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next130_uint_d_ack_ge : bit;
  signal oper_indvar_d_next130_uint_d_ack_top : bit;
  signal oper_indvar_d_next130_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next130_uint_d_req_ge : bit;
  signal oper_indvar_d_next130_uint_d_req_top : bit;
  signal oper_indvar_d_next133_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next133_uint_d_ack_ge : bit;
  signal oper_indvar_d_next133_uint_d_ack_top : bit;
  signal oper_indvar_d_next133_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next133_uint_d_req_ge : bit;
  signal oper_indvar_d_next133_uint_d_req_top : bit;
  signal oper_indvar_d_next139_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next139_uint_d_ack_ge : bit;
  signal oper_indvar_d_next139_uint_d_ack_top : bit;
  signal oper_indvar_d_next139_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next139_uint_d_req_ge : bit;
  signal oper_indvar_d_next139_uint_d_req_top : bit;
  signal oper_indvar_d_next144_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next144_uint_d_ack_ge : bit;
  signal oper_indvar_d_next144_uint_d_ack_top : bit;
  signal oper_indvar_d_next144_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next144_uint_d_req_ge : bit;
  signal oper_indvar_d_next144_uint_d_req_top : bit;
  signal oper_indvar_d_next147_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next147_uint_d_ack_ge : bit;
  signal oper_indvar_d_next147_uint_d_ack_top : bit;
  signal oper_indvar_d_next147_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next147_uint_d_req_ge : bit;
  signal oper_indvar_d_next147_uint_d_req_top : bit;
  signal oper_indvar_d_next149_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next149_uint_d_ack_ge : bit;
  signal oper_indvar_d_next149_uint_d_ack_top : bit;
  signal oper_indvar_d_next149_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next149_uint_d_req_ge : bit;
  signal oper_indvar_d_next149_uint_d_req_top : bit;
  signal oper_indvar_d_next152_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next152_uint_d_ack_ge : bit;
  signal oper_indvar_d_next152_uint_d_ack_top : bit;
  signal oper_indvar_d_next152_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next152_uint_d_req_ge : bit;
  signal oper_indvar_d_next152_uint_d_req_top : bit;
  signal oper_indvar_d_next157_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next157_uint_d_ack_ge : bit;
  signal oper_indvar_d_next157_uint_d_ack_top : bit;
  signal oper_indvar_d_next157_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next157_uint_d_req_ge : bit;
  signal oper_indvar_d_next157_uint_d_req_top : bit;
  signal oper_indvar_d_next_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next_uint_d_ack_ge : bit;
  signal oper_indvar_d_next_uint_d_ack_top : bit;
  signal oper_indvar_d_next_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_indvar_d_next_uint_d_req_ge : bit;
  signal oper_indvar_d_next_uint_d_req_top : bit;
  signal oper_j_d_321_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_j_d_321_int_d_ack_ge : bit;
  signal oper_j_d_321_int_d_ack_top : bit;
  signal oper_j_d_321_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_j_d_321_int_d_req_ge : bit;
  signal oper_j_d_321_int_d_req_top : bit;
  signal oper_j_d_3_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_j_d_3_int_d_ack_ge : bit;
  signal oper_j_d_3_int_d_ack_top : bit;
  signal oper_j_d_3_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_j_d_3_int_d_req_ge : bit;
  signal oper_j_d_3_int_d_req_top : bit;
  signal oper_j_d_746_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_j_d_746_int_d_ack_ge : bit;
  signal oper_j_d_746_int_d_ack_top : bit;
  signal oper_j_d_746_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_j_d_746_int_d_req_ge : bit;
  signal oper_j_d_746_int_d_req_top : bit;
  signal oper_j_d_7_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_j_d_7_int_d_ack_ge : bit;
  signal oper_j_d_7_int_d_ack_top : bit;
  signal oper_j_d_7_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_j_d_7_int_d_req_ge : bit;
  signal oper_j_d_7_int_d_req_top : bit;
  signal oper_k_d_1_d_in_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_k_d_1_d_in_int_d_ack_ge : bit;
  signal oper_k_d_1_d_in_int_d_ack_top : bit;
  signal oper_k_d_1_d_in_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_k_d_1_d_in_int_d_req_ge : bit;
  signal oper_k_d_1_d_in_int_d_req_top : bit;
  signal oper_k_d_1_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_k_d_1_int_d_ack_ge : bit;
  signal oper_k_d_1_int_d_ack_top : bit;
  signal oper_k_d_1_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_k_d_1_int_d_req_ge : bit;
  signal oper_k_d_1_int_d_req_top : bit;
  signal oper_k_d_2_d_2_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_k_d_2_d_2_int_d_ack_ge : bit;
  signal oper_k_d_2_d_2_int_d_ack_top : bit;
  signal oper_k_d_2_d_2_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_k_d_2_d_2_int_d_req_ge : bit;
  signal oper_k_d_2_d_2_int_d_req_top : bit;
  signal oper_k_d_4_d_2_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_k_d_4_d_2_int_d_ack_ge : bit;
  signal oper_k_d_4_d_2_int_d_ack_top : bit;
  signal oper_k_d_4_d_2_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_k_d_4_d_2_int_d_req_ge : bit;
  signal oper_k_d_4_d_2_int_d_req_top : bit;
  signal oper_tmp_d_107_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_107_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_107_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_107_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_107_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_107_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_11348_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11348_bool_d_ack_ge : bit;
  signal oper_tmp_d_11348_bool_d_ack_top : bit;
  signal oper_tmp_d_11348_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11348_bool_d_req_ge : bit;
  signal oper_tmp_d_11348_bool_d_req_top : bit;
  signal oper_tmp_d_113_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_113_bool_d_ack_ge : bit;
  signal oper_tmp_d_113_bool_d_ack_top : bit;
  signal oper_tmp_d_113_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_113_bool_d_req_ge : bit;
  signal oper_tmp_d_113_bool_d_req_top : bit;
  signal oper_tmp_d_118_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_118_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_118_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_118_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_118_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_118_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_11_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_11_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_11_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_11_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_11_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_11_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_125_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_125_uint_d_ack_ge : bit;
  signal oper_tmp_d_125_uint_d_ack_top : bit;
  signal oper_tmp_d_125_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_125_uint_d_req_ge : bit;
  signal oper_tmp_d_125_uint_d_req_top : bit;
  signal oper_tmp_d_132_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_132_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_132_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_132_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_132_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_132_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_132_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_132_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_134_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_134_float_d_ack_ge : bit;
  signal oper_tmp_d_134_float_d_ack_top : bit;
  signal oper_tmp_d_134_float_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_134_float_d_req_ge : bit;
  signal oper_tmp_d_134_float_d_req_top : bit;
  signal oper_tmp_d_135_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_135_float_d_ack_ge : bit;
  signal oper_tmp_d_135_float_d_ack_top : bit;
  signal oper_tmp_d_135_float_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_135_float_d_req_ge : bit;
  signal oper_tmp_d_135_float_d_req_top : bit;
  signal oper_tmp_d_136_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_136_uint_d_ack_ge : bit;
  signal oper_tmp_d_136_uint_d_ack_top : bit;
  signal oper_tmp_d_136_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_136_uint_d_req_ge : bit;
  signal oper_tmp_d_136_uint_d_req_top : bit;
  signal oper_tmp_d_137_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_137_uint_d_ack_ge : bit;
  signal oper_tmp_d_137_uint_d_ack_top : bit;
  signal oper_tmp_d_137_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_137_uint_d_req_ge : bit;
  signal oper_tmp_d_137_uint_d_req_top : bit;
  signal oper_tmp_d_14574_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14574_bool_d_ack_ge : bit;
  signal oper_tmp_d_14574_bool_d_ack_top : bit;
  signal oper_tmp_d_14574_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14574_bool_d_req_ge : bit;
  signal oper_tmp_d_14574_bool_d_req_top : bit;
  signal oper_tmp_d_14578_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14578_bool_d_ack_ge : bit;
  signal oper_tmp_d_14578_bool_d_ack_top : bit;
  signal oper_tmp_d_14578_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14578_bool_d_req_ge : bit;
  signal oper_tmp_d_14578_bool_d_req_top : bit;
  signal oper_tmp_d_14580_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14580_bool_d_ack_ge : bit;
  signal oper_tmp_d_14580_bool_d_ack_top : bit;
  signal oper_tmp_d_14580_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14580_bool_d_req_ge : bit;
  signal oper_tmp_d_14580_bool_d_req_top : bit;
  signal oper_tmp_d_149_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_149_bool_d_ack_ge : bit;
  signal oper_tmp_d_149_bool_d_ack_top : bit;
  signal oper_tmp_d_149_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_149_bool_d_req_ge : bit;
  signal oper_tmp_d_149_bool_d_req_top : bit;
  signal oper_tmp_d_154_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_154_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_154_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_154_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_154_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_154_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_155_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_155_uint_d_ack_ge : bit;
  signal oper_tmp_d_155_uint_d_ack_top : bit;
  signal oper_tmp_d_155_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_155_uint_d_req_ge : bit;
  signal oper_tmp_d_155_uint_d_req_top : bit;
  signal oper_tmp_d_158_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_158_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_158_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_158_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_158_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_158_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_158_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_158_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_1614_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1614_bool_d_ack_ge : bit;
  signal oper_tmp_d_1614_bool_d_ack_top : bit;
  signal oper_tmp_d_1614_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1614_bool_d_req_ge : bit;
  signal oper_tmp_d_1614_bool_d_req_top : bit;
  signal oper_tmp_d_163_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_163_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_163_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_163_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_163_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_163_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_166_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_166_bool_d_ack_ge : bit;
  signal oper_tmp_d_166_bool_d_ack_top : bit;
  signal oper_tmp_d_166_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_166_bool_d_req_ge : bit;
  signal oper_tmp_d_166_bool_d_req_top : bit;
  signal oper_tmp_d_16_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_16_bool_d_ack_ge : bit;
  signal oper_tmp_d_16_bool_d_ack_top : bit;
  signal oper_tmp_d_16_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_16_bool_d_req_ge : bit;
  signal oper_tmp_d_16_bool_d_req_top : bit;
  signal oper_tmp_d_171_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_171_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_171_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_171_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_171_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_171_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_175_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_175_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_175_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_175_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_175_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_175_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_175_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_175_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_179_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_179_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_179_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_179_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_179_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_179_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_179_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_179_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_188_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_188_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_188_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_188_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_188_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_188_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_188_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_188_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_192_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_192_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_192_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_192_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_192_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_192_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_192_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_192_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_20299_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_20299_bool_d_ack_ge : bit;
  signal oper_tmp_d_20299_bool_d_ack_top : bit;
  signal oper_tmp_d_20299_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_20299_bool_d_req_ge : bit;
  signal oper_tmp_d_20299_bool_d_req_top : bit;
  signal oper_tmp_d_202_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_202_bool_d_ack_ge : bit;
  signal oper_tmp_d_202_bool_d_ack_top : bit;
  signal oper_tmp_d_202_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_202_bool_d_req_ge : bit;
  signal oper_tmp_d_202_bool_d_req_top : bit;
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_ack_ge : bit;
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_ack_top : bit;
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_req_ge : bit;
  signal oper_tmp_d_206_d_lvl_d_0_uint_d_req_top : bit;
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_ack_ge : bit;
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_ack_top : bit;
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_req_ge : bit;
  signal oper_tmp_d_20_d_lvl_d_0_uint_d_req_top : bit;
  signal oper_tmp_d_210_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_210_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_210_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_210_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_210_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_210_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_221111_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_221111_bool_d_ack_ge : bit;
  signal oper_tmp_d_221111_bool_d_ack_top : bit;
  signal oper_tmp_d_221111_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_221111_bool_d_req_ge : bit;
  signal oper_tmp_d_221111_bool_d_req_top : bit;
  signal oper_tmp_d_221_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_221_bool_d_ack_ge : bit;
  signal oper_tmp_d_221_bool_d_ack_top : bit;
  signal oper_tmp_d_221_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_221_bool_d_req_ge : bit;
  signal oper_tmp_d_221_bool_d_req_top : bit;
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_ack_ge : bit;
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_ack_top : bit;
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_req_ge : bit;
  signal oper_tmp_d_225_d_lvl_d_0_uint_d_req_top : bit;
  signal oper_tmp_d_229_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_229_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_229_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_229_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_229_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_229_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_229_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_229_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_ack_ge : bit;
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_ack_top : bit;
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_req_ge : bit;
  signal oper_tmp_d_25_d_lvl_d_0_uint_d_req_top : bit;
  signal oper_tmp_d_27_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_27_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_27_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_27_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_27_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_27_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_27_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_27_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_ack_ge : bit;
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_ack_top : bit;
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_req_ge : bit;
  signal oper_tmp_d_30_d_lvl_d_0_uint_d_req_top : bit;
  signal oper_tmp_d_4223_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_4223_bool_d_ack_ge : bit;
  signal oper_tmp_d_4223_bool_d_ack_top : bit;
  signal oper_tmp_d_4223_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_4223_bool_d_req_ge : bit;
  signal oper_tmp_d_4223_bool_d_req_top : bit;
  signal oper_tmp_d_42_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_42_bool_d_ack_ge : bit;
  signal oper_tmp_d_42_bool_d_ack_top : bit;
  signal oper_tmp_d_42_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_42_bool_d_req_ge : bit;
  signal oper_tmp_d_42_bool_d_req_top : bit;
  signal oper_tmp_d_47_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_47_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_47_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_47_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_47_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_47_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_52_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_52_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_52_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_52_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_52_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_52_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_54_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_54_bool_d_ack_ge : bit;
  signal oper_tmp_d_54_bool_d_ack_top : bit;
  signal oper_tmp_d_54_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_54_bool_d_req_ge : bit;
  signal oper_tmp_d_54_bool_d_req_top : bit;
  signal oper_tmp_d_65_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_65_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_65_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_65_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_65_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_65_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_74_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_74_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_74_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_74_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_74_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_74_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_92_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_92_bool_d_ack_ge : bit;
  signal oper_tmp_d_92_bool_d_ack_top : bit;
  signal oper_tmp_d_92_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_92_bool_d_req_ge : bit;
  signal oper_tmp_d_92_bool_d_req_top : bit;
  signal oper_tmp_d_97_d_id_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_id_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_97_d_id_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_97_d_id_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_id_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_97_d_id_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_ack_ge : bit;
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_ack_top : bit;
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_req_ge : bit;
  signal oper_tmp_d_97_d_lvl_d_1_uint_d_req_top : bit;
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_ack_ge : bit;
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_ack_top : bit;
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_req_ge : bit;
  signal oper_tmp_d_97_d_lvl_d_2_uint_d_req_top : bit;
  signal oper_tmp_d_uint_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_uint_d_ack_ge : bit;
  signal oper_tmp_d_uint_d_ack_top : bit;
  signal oper_tmp_d_uint_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_uint_d_req_ge : bit;
  signal oper_tmp_d_uint_d_req_top : bit;
  signal start_call_divide_0_actual_0_wr_d_ack_tip : bit_vector(0 downto 0);
  signal start_call_divide_0_actual_0_wr_d_ack_ge : bit;
  signal start_call_divide_0_actual_0_wr_d_ack_top : bit;
  signal start_call_divide_0_actual_0_wr_d_req_tip : bit_vector(1 downto 0);
  signal start_call_divide_0_actual_0_wr_d_req_ge : bit;
  signal start_call_divide_0_actual_0_wr_d_req_top : bit;
  signal start_call_divide_0_actual_1_wr_d_ack_tip : bit_vector(0 downto 0);
  signal start_call_divide_0_actual_1_wr_d_ack_ge : bit;
  signal start_call_divide_0_actual_1_wr_d_ack_top : bit;
  signal start_call_divide_0_actual_1_wr_d_req_tip : bit_vector(1 downto 0);
  signal start_call_divide_0_actual_1_wr_d_req_ge : bit;
  signal start_call_divide_0_actual_1_wr_d_req_top : bit;
  signal start_call_divide_0_d_ack_tip : bit_vector(0 downto 0);
  signal start_call_divide_0_d_ack_ge : bit;
  signal start_call_divide_0_d_ack_top : bit;
  signal start_call_divide_0_d_req_tip : bit_vector(0 downto 0);
  signal start_call_divide_0_d_req_ge : bit;
  signal start_call_divide_0_d_req_top : bit;
  signal store_0_d_ack_tip : bit_vector(0 downto 0);
  signal store_0_d_ack_ge : bit;
  signal store_0_d_ack_top : bit;
  signal store_0_d_req_tip : bit_vector(0 downto 0);
  signal store_0_d_req_ge : bit;
  signal store_0_d_req_top : bit;
  signal store_10_d_ack_tip : bit_vector(0 downto 0);
  signal store_10_d_ack_ge : bit;
  signal store_10_d_ack_top : bit;
  signal store_10_d_req_tip : bit_vector(0 downto 0);
  signal store_10_d_req_ge : bit;
  signal store_10_d_req_top : bit;
  signal store_11_d_ack_tip : bit_vector(0 downto 0);
  signal store_11_d_ack_ge : bit;
  signal store_11_d_ack_top : bit;
  signal store_11_d_req_tip : bit_vector(2 downto 0);
  signal store_11_d_req_ge : bit;
  signal store_11_d_req_top : bit;
  signal store_12_d_ack_tip : bit_vector(0 downto 0);
  signal store_12_d_ack_ge : bit;
  signal store_12_d_ack_top : bit;
  signal store_12_d_req_tip : bit_vector(2 downto 0);
  signal store_12_d_req_ge : bit;
  signal store_12_d_req_top : bit;
  signal store_13_d_ack_tip : bit_vector(0 downto 0);
  signal store_13_d_ack_ge : bit;
  signal store_13_d_ack_top : bit;
  signal store_13_d_req_tip : bit_vector(2 downto 0);
  signal store_13_d_req_ge : bit;
  signal store_13_d_req_top : bit;
  signal store_1_d_ack_tip : bit_vector(0 downto 0);
  signal store_1_d_ack_ge : bit;
  signal store_1_d_ack_top : bit;
  signal store_1_d_req_tip : bit_vector(2 downto 0);
  signal store_1_d_req_ge : bit;
  signal store_1_d_req_top : bit;
  signal store_2_d_ack_tip : bit_vector(0 downto 0);
  signal store_2_d_ack_ge : bit;
  signal store_2_d_ack_top : bit;
  signal store_2_d_req_tip : bit_vector(2 downto 0);
  signal store_2_d_req_ge : bit;
  signal store_2_d_req_top : bit;
  signal store_3_d_ack_tip : bit_vector(0 downto 0);
  signal store_3_d_ack_ge : bit;
  signal store_3_d_ack_top : bit;
  signal store_3_d_req_tip : bit_vector(2 downto 0);
  signal store_3_d_req_ge : bit;
  signal store_3_d_req_top : bit;
  signal store_4_d_ack_tip : bit_vector(0 downto 0);
  signal store_4_d_ack_ge : bit;
  signal store_4_d_ack_top : bit;
  signal store_4_d_req_tip : bit_vector(2 downto 0);
  signal store_4_d_req_ge : bit;
  signal store_4_d_req_top : bit;
  signal store_5_d_ack_tip : bit_vector(0 downto 0);
  signal store_5_d_ack_ge : bit;
  signal store_5_d_ack_top : bit;
  signal store_5_d_req_tip : bit_vector(2 downto 0);
  signal store_5_d_req_ge : bit;
  signal store_5_d_req_top : bit;
  signal store_6_d_ack_tip : bit_vector(0 downto 0);
  signal store_6_d_ack_ge : bit;
  signal store_6_d_ack_top : bit;
  signal store_6_d_req_tip : bit_vector(2 downto 0);
  signal store_6_d_req_ge : bit;
  signal store_6_d_req_top : bit;
  signal store_7_d_ack_tip : bit_vector(0 downto 0);
  signal store_7_d_ack_ge : bit;
  signal store_7_d_ack_top : bit;
  signal store_7_d_req_tip : bit_vector(1 downto 0);
  signal store_7_d_req_ge : bit;
  signal store_7_d_req_top : bit;
  signal store_8_d_ack_tip : bit_vector(0 downto 0);
  signal store_8_d_ack_ge : bit;
  signal store_8_d_ack_top : bit;
  signal store_8_d_req_tip : bit_vector(0 downto 0);
  signal store_8_d_req_ge : bit;
  signal store_8_d_req_top : bit;
  signal store_9_d_ack_tip : bit_vector(0 downto 0);
  signal store_9_d_ack_ge : bit;
  signal store_9_d_ack_top : bit;
  signal store_9_d_req_tip : bit_vector(2 downto 0);
  signal store_9_d_req_ge : bit;
  signal store_9_d_req_top : bit;
  signal tc_i_d_1_d_0_d_ack_tip : bit_vector(0 downto 0);
  signal tc_i_d_1_d_0_d_ack_ge : bit;
  signal tc_i_d_1_d_0_d_ack_top : bit;
  signal tc_i_d_1_d_0_d_req_tip : bit_vector(0 downto 0);
  signal tc_i_d_1_d_0_d_req_ge : bit;
  signal tc_i_d_1_d_0_d_req_top : bit;
  signal tc_i_d_2_d_0_d_ph_d_ack_tip : bit_vector(0 downto 0);
  signal tc_i_d_2_d_0_d_ph_d_ack_ge : bit;
  signal tc_i_d_2_d_0_d_ph_d_ack_top : bit;
  signal tc_i_d_2_d_0_d_ph_d_req_tip : bit_vector(0 downto 0);
  signal tc_i_d_2_d_0_d_ph_d_req_ge : bit;
  signal tc_i_d_2_d_0_d_ph_d_req_top : bit;
  signal tc_i_d_3_d_0_d_ph_d_ack_tip : bit_vector(0 downto 0);
  signal tc_i_d_3_d_0_d_ph_d_ack_ge : bit;
  signal tc_i_d_3_d_0_d_ph_d_ack_top : bit;
  signal tc_i_d_3_d_0_d_ph_d_req_tip : bit_vector(0 downto 0);
  signal tc_i_d_3_d_0_d_ph_d_req_ge : bit;
  signal tc_i_d_3_d_0_d_ph_d_req_top : bit;
  signal tc_i_d_4_d_0_d_ack_tip : bit_vector(0 downto 0);
  signal tc_i_d_4_d_0_d_ack_ge : bit;
  signal tc_i_d_4_d_0_d_ack_top : bit;
  signal tc_i_d_4_d_0_d_req_tip : bit_vector(0 downto 0);
  signal tc_i_d_4_d_0_d_req_ge : bit;
  signal tc_i_d_4_d_0_d_req_top : bit;
  signal tc_i_d_5_d_0_d_ack_tip : bit_vector(0 downto 0);
  signal tc_i_d_5_d_0_d_ack_ge : bit;
  signal tc_i_d_5_d_0_d_ack_top : bit;
  signal tc_i_d_5_d_0_d_req_tip : bit_vector(0 downto 0);
  signal tc_i_d_5_d_0_d_req_ge : bit;
  signal tc_i_d_5_d_0_d_req_top : bit;
  signal tc_indvar138_d_ack_tip : bit_vector(0 downto 0);
  signal tc_indvar138_d_ack_ge : bit;
  signal tc_indvar138_d_ack_top : bit;
  signal tc_indvar138_d_req_tip : bit_vector(0 downto 0);
  signal tc_indvar138_d_req_ge : bit;
  signal tc_indvar138_d_req_top : bit;
  signal tc_indvar151_d_ack_tip : bit_vector(0 downto 0);
  signal tc_indvar151_d_ack_ge : bit;
  signal tc_indvar151_d_ack_top : bit;
  signal tc_indvar151_d_req_tip : bit_vector(0 downto 0);
  signal tc_indvar151_d_req_ge : bit;
  signal tc_indvar151_d_req_top : bit;
  signal tc_j_d_11_d_2_d_ack_tip : bit_vector(0 downto 0);
  signal tc_j_d_11_d_2_d_ack_ge : bit;
  signal tc_j_d_11_d_2_d_ack_top : bit;
  signal tc_j_d_11_d_2_d_req_tip : bit_vector(0 downto 0);
  signal tc_j_d_11_d_2_d_req_ge : bit;
  signal tc_j_d_11_d_2_d_req_top : bit;
  signal tc_j_d_13_d_2_d_ack_tip : bit_vector(0 downto 0);
  signal tc_j_d_13_d_2_d_ack_ge : bit;
  signal tc_j_d_13_d_2_d_ack_top : bit;
  signal tc_j_d_13_d_2_d_req_tip : bit_vector(0 downto 0);
  signal tc_j_d_13_d_2_d_req_ge : bit;
  signal tc_j_d_13_d_2_d_req_top : bit;
  signal tc_j_d_3_d_2_d_ack_tip : bit_vector(0 downto 0);
  signal tc_j_d_3_d_2_d_ack_ge : bit;
  signal tc_j_d_3_d_2_d_ack_top : bit;
  signal tc_j_d_3_d_2_d_req_tip : bit_vector(0 downto 0);
  signal tc_j_d_3_d_2_d_req_ge : bit;
  signal tc_j_d_3_d_2_d_req_top : bit;
  signal tc_j_d_3_d_in_d_ack_tip : bit_vector(0 downto 0);
  signal tc_j_d_3_d_in_d_ack_ge : bit;
  signal tc_j_d_3_d_in_d_ack_top : bit;
  signal tc_j_d_3_d_in_d_req_tip : bit_vector(0 downto 0);
  signal tc_j_d_3_d_in_d_req_ge : bit;
  signal tc_j_d_3_d_in_d_req_top : bit;
  signal tc_j_d_7_d_1_d_ack_tip : bit_vector(0 downto 0);
  signal tc_j_d_7_d_1_d_ack_ge : bit;
  signal tc_j_d_7_d_1_d_ack_top : bit;
  signal tc_j_d_7_d_1_d_req_tip : bit_vector(0 downto 0);
  signal tc_j_d_7_d_1_d_req_ge : bit;
  signal tc_j_d_7_d_1_d_req_top : bit;
  signal tc_p_d_0_d_0_d_ph_d_ack_tip : bit_vector(0 downto 0);
  signal tc_p_d_0_d_0_d_ph_d_ack_ge : bit;
  signal tc_p_d_0_d_0_d_ph_d_ack_top : bit;
  signal tc_p_d_0_d_0_d_ph_d_req_tip : bit_vector(0 downto 0);
  signal tc_p_d_0_d_0_d_ph_d_req_ge : bit;
  signal tc_p_d_0_d_0_d_ph_d_req_top : bit;
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_ack_top : bit;
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_req_ge : bit;
  signal tc_tmp_d_118_d_id_d_1_d_cast_d_req_top : bit;
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_154_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_158_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_163_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_171_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_175_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_179_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_188_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_192_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_ack_top : bit;
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_req_ge : bit;
  signal tc_tmp_d_206_d_id_d_0_d_cast_d_req_top : bit;
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_ack_top : bit;
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_req_ge : bit;
  signal tc_tmp_d_225_d_id_d_0_d_cast_d_req_top : bit;
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_ack_top : bit;
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_req_ge : bit;
  signal tc_tmp_d_27_d_id_d_1_d_cast_d_req_top : bit;
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_ack_top : bit;
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_req_ge : bit;
  signal tc_tmp_d_27_d_id_d_2_d_cast_d_req_top : bit;
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_ack_top : bit;
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_req_ge : bit;
  signal tc_tmp_d_74_d_id_d_1_d_cast_d_req_top : bit;
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_ack_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_ack_ge : bit;
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_ack_top : bit;
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_req_tip : bit_vector(0 downto 0);
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_req_ge : bit;
  signal tc_tmp_d_97_d_id_d_1_d_cast_d_req_top : bit;
  signal then_d_0_d_entry_tip : bit_vector(0 downto 0);
  signal then_d_0_d_entry_ge : bit;
  signal then_d_0_d_entry_top : bit;
  signal then_d_0_to_no_exit_d_4_src_tip : bit_vector(0 downto 0);
  signal then_d_0_to_no_exit_d_4_src_ge : bit;
  signal then_d_0_to_no_exit_d_4_src_top : bit;
  signal then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_tip : bit_vector(0 downto 0);
  signal then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_ge : bit;
  signal then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_top : bit;
  signal then_d_1_d_entry_tip : bit_vector(0 downto 0);
  signal then_d_1_d_entry_ge : bit;
  signal then_d_1_d_entry_top : bit;
  signal then_d_1_to_loopexit_d_10_src_tip : bit_vector(0 downto 0);
  signal then_d_1_to_loopexit_d_10_src_ge : bit;
  signal then_d_1_to_loopexit_d_10_src_top : bit;
  signal then_d_1_to_no_exit_d_10_d_backedge_src_tip : bit_vector(0 downto 0);
  signal then_d_1_to_no_exit_d_10_d_backedge_src_ge : bit;
  signal then_d_1_to_no_exit_d_10_d_backedge_src_top : bit;
  signal then_d_2_d_entry_tip : bit_vector(0 downto 0);
  signal then_d_2_d_entry_ge : bit;
  signal then_d_2_d_entry_top : bit;
  signal then_d_2_to_loopexit_d_10_src_tip : bit_vector(0 downto 0);
  signal then_d_2_to_loopexit_d_10_src_ge : bit;
  signal then_d_2_to_loopexit_d_10_src_top : bit;
  signal then_d_2_to_no_exit_d_10_d_backedge_src_tip : bit_vector(0 downto 0);
  signal then_d_2_to_no_exit_d_10_d_backedge_src_ge : bit;
  signal then_d_2_to_no_exit_d_10_d_backedge_src_top : bit;

begin


  place_1 : place
  generic map(1, 1, '0')
  port map(place_1_tip, place_1_rst, place_1_top, reset, clk);

  place_100 : place
  generic map(2, 1, '0')
  port map(place_100_tip, place_100_rst, place_100_top, reset, clk);

  place_101 : place
  generic map(1, 1, '0')
  port map(place_101_tip, place_101_rst, place_101_top, reset, clk);

  place_105 : place
  generic map(2, 1, '0')
  port map(place_105_tip, place_105_rst, place_105_top, reset, clk);

  place_106 : place
  generic map(1, 1, '0')
  port map(place_106_tip, place_106_rst, place_106_top, reset, clk);

  place_107 : place
  generic map(1, 1, '0')
  port map(place_107_tip, place_107_rst, place_107_top, reset, clk);

  place_108 : place
  generic map(1, 1, '0')
  port map(place_108_tip, place_108_rst, place_108_top, reset, clk);

  place_109 : place
  generic map(1, 1, '0')
  port map(place_109_tip, place_109_rst, place_109_top, reset, clk);

  place_110 : place
  generic map(1, 1, '0')
  port map(place_110_tip, place_110_rst, place_110_top, reset, clk);

  place_111 : place
  generic map(1, 1, '0')
  port map(place_111_tip, place_111_rst, place_111_top, reset, clk);

  place_112 : place
  generic map(1, 1, '0')
  port map(place_112_tip, place_112_rst, place_112_top, reset, clk);

  place_113 : place
  generic map(1, 1, '0')
  port map(place_113_tip, place_113_rst, place_113_top, reset, clk);

  place_114 : place
  generic map(1, 1, '0')
  port map(place_114_tip, place_114_rst, place_114_top, reset, clk);

  place_115 : place
  generic map(1, 1, '0')
  port map(place_115_tip, place_115_rst, place_115_top, reset, clk);

  place_116 : place
  generic map(1, 1, '0')
  port map(place_116_tip, place_116_rst, place_116_top, reset, clk);

  place_117 : place
  generic map(1, 1, '0')
  port map(place_117_tip, place_117_rst, place_117_top, reset, clk);

  place_118 : place
  generic map(1, 1, '0')
  port map(place_118_tip, place_118_rst, place_118_top, reset, clk);

  place_119 : place
  generic map(1, 1, '0')
  port map(place_119_tip, place_119_rst, place_119_top, reset, clk);

  place_120 : place
  generic map(1, 1, '0')
  port map(place_120_tip, place_120_rst, place_120_top, reset, clk);

  place_121 : place
  generic map(1, 1, '0')
  port map(place_121_tip, place_121_rst, place_121_top, reset, clk);

  place_122 : place
  generic map(1, 2, '0')
  port map(place_122_tip, place_122_rst, place_122_top, reset, clk);

  place_123 : place
  generic map(1, 1, '0')
  port map(place_123_tip, place_123_rst, place_123_top, reset, clk);

  place_124 : place
  generic map(1, 1, '0')
  port map(place_124_tip, place_124_rst, place_124_top, reset, clk);

  place_126 : place
  generic map(1, 1, '0')
  port map(place_126_tip, place_126_rst, place_126_top, reset, clk);

  place_127 : place
  generic map(1, 1, '0')
  port map(place_127_tip, place_127_rst, place_127_top, reset, clk);

  place_128 : place
  generic map(1, 1, '0')
  port map(place_128_tip, place_128_rst, place_128_top, reset, clk);

  place_129 : place
  generic map(1, 2, '0')
  port map(place_129_tip, place_129_rst, place_129_top, reset, clk);

  place_130 : place
  generic map(1, 1, '0')
  port map(place_130_tip, place_130_rst, place_130_top, reset, clk);

  place_132 : place
  generic map(1, 1, '0')
  port map(place_132_tip, place_132_rst, place_132_top, reset, clk);

  place_133 : place
  generic map(1, 2, '0')
  port map(place_133_tip, place_133_rst, place_133_top, reset, clk);

  place_136 : place
  generic map(2, 1, '0')
  port map(place_136_tip, place_136_rst, place_136_top, reset, clk);

  place_137 : place
  generic map(1, 1, '0')
  port map(place_137_tip, place_137_rst, place_137_top, reset, clk);

  place_138 : place
  generic map(1, 1, '0')
  port map(place_138_tip, place_138_rst, place_138_top, reset, clk);

  place_139 : place
  generic map(1, 1, '0')
  port map(place_139_tip, place_139_rst, place_139_top, reset, clk);

  place_14 : place
  generic map(2, 1, '0')
  port map(place_14_tip, place_14_rst, place_14_top, reset, clk);

  place_140 : place
  generic map(1, 1, '0')
  port map(place_140_tip, place_140_rst, place_140_top, reset, clk);

  place_141 : place
  generic map(1, 1, '0')
  port map(place_141_tip, place_141_rst, place_141_top, reset, clk);

  place_142 : place
  generic map(1, 1, '0')
  port map(place_142_tip, place_142_rst, place_142_top, reset, clk);

  place_143 : place
  generic map(1, 1, '0')
  port map(place_143_tip, place_143_rst, place_143_top, reset, clk);

  place_144 : place
  generic map(1, 1, '0')
  port map(place_144_tip, place_144_rst, place_144_top, reset, clk);

  place_145 : place
  generic map(1, 1, '0')
  port map(place_145_tip, place_145_rst, place_145_top, reset, clk);

  place_146 : place
  generic map(1, 1, '0')
  port map(place_146_tip, place_146_rst, place_146_top, reset, clk);

  place_147 : place
  generic map(1, 1, '0')
  port map(place_147_tip, place_147_rst, place_147_top, reset, clk);

  place_148 : place
  generic map(1, 1, '0')
  port map(place_148_tip, place_148_rst, place_148_top, reset, clk);

  place_149 : place
  generic map(1, 1, '0')
  port map(place_149_tip, place_149_rst, place_149_top, reset, clk);

  place_150 : place
  generic map(1, 1, '0')
  port map(place_150_tip, place_150_rst, place_150_top, reset, clk);

  place_151 : place
  generic map(1, 1, '0')
  port map(place_151_tip, place_151_rst, place_151_top, reset, clk);

  place_152 : place
  generic map(1, 1, '0')
  port map(place_152_tip, place_152_rst, place_152_top, reset, clk);

  place_153 : place
  generic map(1, 1, '0')
  port map(place_153_tip, place_153_rst, place_153_top, reset, clk);

  place_154 : place
  generic map(1, 1, '0')
  port map(place_154_tip, place_154_rst, place_154_top, reset, clk);

  place_155 : place
  generic map(1, 1, '0')
  port map(place_155_tip, place_155_rst, place_155_top, reset, clk);

  place_156 : place
  generic map(1, 1, '0')
  port map(place_156_tip, place_156_rst, place_156_top, reset, clk);

  place_157 : place
  generic map(1, 1, '0')
  port map(place_157_tip, place_157_rst, place_157_top, reset, clk);

  place_158 : place
  generic map(1, 1, '0')
  port map(place_158_tip, place_158_rst, place_158_top, reset, clk);

  place_159 : place
  generic map(1, 1, '0')
  port map(place_159_tip, place_159_rst, place_159_top, reset, clk);

  place_16 : place
  generic map(1, 1, '0')
  port map(place_16_tip, place_16_rst, place_16_top, reset, clk);

  place_160 : place
  generic map(1, 1, '0')
  port map(place_160_tip, place_160_rst, place_160_top, reset, clk);

  place_161 : place
  generic map(1, 1, '0')
  port map(place_161_tip, place_161_rst, place_161_top, reset, clk);

  place_162 : place
  generic map(1, 1, '0')
  port map(place_162_tip, place_162_rst, place_162_top, reset, clk);

  place_163 : place
  generic map(1, 1, '0')
  port map(place_163_tip, place_163_rst, place_163_top, reset, clk);

  place_164 : place
  generic map(1, 1, '0')
  port map(place_164_tip, place_164_rst, place_164_top, reset, clk);

  place_165 : place
  generic map(1, 1, '0')
  port map(place_165_tip, place_165_rst, place_165_top, reset, clk);

  place_166 : place
  generic map(1, 1, '0')
  port map(place_166_tip, place_166_rst, place_166_top, reset, clk);

  place_167 : place
  generic map(1, 1, '0')
  port map(place_167_tip, place_167_rst, place_167_top, reset, clk);

  place_168 : place
  generic map(1, 1, '0')
  port map(place_168_tip, place_168_rst, place_168_top, reset, clk);

  place_169 : place
  generic map(1, 1, '0')
  port map(place_169_tip, place_169_rst, place_169_top, reset, clk);

  place_17 : place
  generic map(1, 1, '0')
  port map(place_17_tip, place_17_rst, place_17_top, reset, clk);

  place_170 : place
  generic map(1, 1, '0')
  port map(place_170_tip, place_170_rst, place_170_top, reset, clk);

  place_171 : place
  generic map(1, 1, '0')
  port map(place_171_tip, place_171_rst, place_171_top, reset, clk);

  place_172 : place
  generic map(1, 1, '0')
  port map(place_172_tip, place_172_rst, place_172_top, reset, clk);

  place_173 : place
  generic map(1, 1, '0')
  port map(place_173_tip, place_173_rst, place_173_top, reset, clk);

  place_174 : place
  generic map(1, 1, '0')
  port map(place_174_tip, place_174_rst, place_174_top, reset, clk);

  place_175 : place
  generic map(1, 1, '0')
  port map(place_175_tip, place_175_rst, place_175_top, reset, clk);

  place_176 : place
  generic map(1, 1, '0')
  port map(place_176_tip, place_176_rst, place_176_top, reset, clk);

  place_177 : place
  generic map(1, 1, '0')
  port map(place_177_tip, place_177_rst, place_177_top, reset, clk);

  place_178 : place
  generic map(1, 1, '0')
  port map(place_178_tip, place_178_rst, place_178_top, reset, clk);

  place_179 : place
  generic map(1, 2, '0')
  port map(place_179_tip, place_179_rst, place_179_top, reset, clk);

  place_180 : place
  generic map(1, 1, '0')
  port map(place_180_tip, place_180_rst, place_180_top, reset, clk);

  place_183 : place
  generic map(1, 1, '0')
  port map(place_183_tip, place_183_rst, place_183_top, reset, clk);

  place_184 : place
  generic map(2, 1, '0')
  port map(place_184_tip, place_184_rst, place_184_top, reset, clk);

  place_185 : place
  generic map(1, 1, '0')
  port map(place_185_tip, place_185_rst, place_185_top, reset, clk);

  place_186 : place
  generic map(1, 1, '0')
  port map(place_186_tip, place_186_rst, place_186_top, reset, clk);

  place_187 : place
  generic map(1, 1, '0')
  port map(place_187_tip, place_187_rst, place_187_top, reset, clk);

  place_188 : place
  generic map(2, 1, '0')
  port map(place_188_tip, place_188_rst, place_188_top, reset, clk);

  place_189 : place
  generic map(1, 1, '0')
  port map(place_189_tip, place_189_rst, place_189_top, reset, clk);

  place_190 : place
  generic map(1, 1, '0')
  port map(place_190_tip, place_190_rst, place_190_top, reset, clk);

  place_191 : place
  generic map(1, 1, '0')
  port map(place_191_tip, place_191_rst, place_191_top, reset, clk);

  place_192 : place
  generic map(1, 1, '0')
  port map(place_192_tip, place_192_rst, place_192_top, reset, clk);

  place_193 : place
  generic map(2, 1, '0')
  port map(place_193_tip, place_193_rst, place_193_top, reset, clk);

  place_194 : place
  generic map(1, 1, '0')
  port map(place_194_tip, place_194_rst, place_194_top, reset, clk);

  place_195 : place
  generic map(1, 1, '0')
  port map(place_195_tip, place_195_rst, place_195_top, reset, clk);

  place_196 : place
  generic map(1, 1, '0')
  port map(place_196_tip, place_196_rst, place_196_top, reset, clk);

  place_197 : place
  generic map(1, 1, '0')
  port map(place_197_tip, place_197_rst, place_197_top, reset, clk);

  place_198 : place
  generic map(1, 1, '0')
  port map(place_198_tip, place_198_rst, place_198_top, reset, clk);

  place_199 : place
  generic map(1, 1, '0')
  port map(place_199_tip, place_199_rst, place_199_top, reset, clk);

  place_20 : place
  generic map(1, 1, '0')
  port map(place_20_tip, place_20_rst, place_20_top, reset, clk);

  place_200 : place
  generic map(1, 1, '0')
  port map(place_200_tip, place_200_rst, place_200_top, reset, clk);

  place_201 : place
  generic map(1, 1, '0')
  port map(place_201_tip, place_201_rst, place_201_top, reset, clk);

  place_202 : place
  generic map(1, 1, '0')
  port map(place_202_tip, place_202_rst, place_202_top, reset, clk);

  place_203 : place
  generic map(1, 1, '0')
  port map(place_203_tip, place_203_rst, place_203_top, reset, clk);

  place_204 : place
  generic map(1, 1, '0')
  port map(place_204_tip, place_204_rst, place_204_top, reset, clk);

  place_205 : place
  generic map(1, 1, '0')
  port map(place_205_tip, place_205_rst, place_205_top, reset, clk);

  place_206 : place
  generic map(1, 1, '0')
  port map(place_206_tip, place_206_rst, place_206_top, reset, clk);

  place_208 : place
  generic map(1, 1, '0')
  port map(place_208_tip, place_208_rst, place_208_top, reset, clk);

  place_209 : place
  generic map(2, 1, '0')
  port map(place_209_tip, place_209_rst, place_209_top, reset, clk);

  place_210 : place
  generic map(1, 1, '0')
  port map(place_210_tip, place_210_rst, place_210_top, reset, clk);

  place_211 : place
  generic map(1, 1, '0')
  port map(place_211_tip, place_211_rst, place_211_top, reset, clk);

  place_212 : place
  generic map(1, 1, '0')
  port map(place_212_tip, place_212_rst, place_212_top, reset, clk);

  place_213 : place
  generic map(2, 1, '0')
  port map(place_213_tip, place_213_rst, place_213_top, reset, clk);

  place_214 : place
  generic map(1, 1, '0')
  port map(place_214_tip, place_214_rst, place_214_top, reset, clk);

  place_215 : place
  generic map(1, 1, '0')
  port map(place_215_tip, place_215_rst, place_215_top, reset, clk);

  place_216 : place
  generic map(1, 1, '0')
  port map(place_216_tip, place_216_rst, place_216_top, reset, clk);

  place_217 : place
  generic map(1, 1, '0')
  port map(place_217_tip, place_217_rst, place_217_top, reset, clk);

  place_218 : place
  generic map(1, 1, '0')
  port map(place_218_tip, place_218_rst, place_218_top, reset, clk);

  place_219 : place
  generic map(1, 1, '0')
  port map(place_219_tip, place_219_rst, place_219_top, reset, clk);

  place_22 : place
  generic map(1, 1, '0')
  port map(place_22_tip, place_22_rst, place_22_top, reset, clk);

  place_220 : place
  generic map(1, 1, '0')
  port map(place_220_tip, place_220_rst, place_220_top, reset, clk);

  place_221 : place
  generic map(1, 1, '0')
  port map(place_221_tip, place_221_rst, place_221_top, reset, clk);

  place_222 : place
  generic map(1, 2, '0')
  port map(place_222_tip, place_222_rst, place_222_top, reset, clk);

  place_223 : place
  generic map(1, 1, '0')
  port map(place_223_tip, place_223_rst, place_223_top, reset, clk);

  place_224 : place
  generic map(1, 1, '0')
  port map(place_224_tip, place_224_rst, place_224_top, reset, clk);

  place_225 : place
  generic map(1, 1, '0')
  port map(place_225_tip, place_225_rst, place_225_top, reset, clk);

  place_226 : place
  generic map(1, 1, '0')
  port map(place_226_tip, place_226_rst, place_226_top, reset, clk);

  place_227 : place
  generic map(1, 1, '0')
  port map(place_227_tip, place_227_rst, place_227_top, reset, clk);

  place_228 : place
  generic map(1, 1, '0')
  port map(place_228_tip, place_228_rst, place_228_top, reset, clk);

  place_229 : place
  generic map(1, 1, '0')
  port map(place_229_tip, place_229_rst, place_229_top, reset, clk);

  place_230 : place
  generic map(1, 1, '0')
  port map(place_230_tip, place_230_rst, place_230_top, reset, clk);

  place_231 : place
  generic map(1, 1, '0')
  port map(place_231_tip, place_231_rst, place_231_top, reset, clk);

  place_232 : place
  generic map(2, 1, '0')
  port map(place_232_tip, place_232_rst, place_232_top, reset, clk);

  place_233 : place
  generic map(1, 1, '0')
  port map(place_233_tip, place_233_rst, place_233_top, reset, clk);

  place_234 : place
  generic map(1, 1, '0')
  port map(place_234_tip, place_234_rst, place_234_top, reset, clk);

  place_235 : place
  generic map(1, 1, '0')
  port map(place_235_tip, place_235_rst, place_235_top, reset, clk);

  place_236 : place
  generic map(2, 1, '0')
  port map(place_236_tip, place_236_rst, place_236_top, reset, clk);

  place_237 : place
  generic map(1, 1, '0')
  port map(place_237_tip, place_237_rst, place_237_top, reset, clk);

  place_238 : place
  generic map(1, 1, '0')
  port map(place_238_tip, place_238_rst, place_238_top, reset, clk);

  place_239 : place
  generic map(1, 1, '0')
  port map(place_239_tip, place_239_rst, place_239_top, reset, clk);

  place_24 : place
  generic map(1, 1, '0')
  port map(place_24_tip, place_24_rst, place_24_top, reset, clk);

  place_240 : place
  generic map(1, 1, '0')
  port map(place_240_tip, place_240_rst, place_240_top, reset, clk);

  place_241 : place
  generic map(1, 1, '0')
  port map(place_241_tip, place_241_rst, place_241_top, reset, clk);

  place_242 : place
  generic map(1, 1, '0')
  port map(place_242_tip, place_242_rst, place_242_top, reset, clk);

  place_243 : place
  generic map(1, 1, '0')
  port map(place_243_tip, place_243_rst, place_243_top, reset, clk);

  place_244 : place
  generic map(1, 1, '0')
  port map(place_244_tip, place_244_rst, place_244_top, reset, clk);

  place_245 : place
  generic map(1, 1, '0')
  port map(place_245_tip, place_245_rst, place_245_top, reset, clk);

  place_246 : place
  generic map(1, 1, '0')
  port map(place_246_tip, place_246_rst, place_246_top, reset, clk);

  place_247 : place
  generic map(1, 1, '0')
  port map(place_247_tip, place_247_rst, place_247_top, reset, clk);

  place_248 : place
  generic map(1, 1, '0')
  port map(place_248_tip, place_248_rst, place_248_top, reset, clk);

  place_249 : place
  generic map(1, 1, '0')
  port map(place_249_tip, place_249_rst, place_249_top, reset, clk);

  place_25 : place
  generic map(1, 1, '0')
  port map(place_25_tip, place_25_rst, place_25_top, reset, clk);

  place_250 : place
  generic map(1, 1, '0')
  port map(place_250_tip, place_250_rst, place_250_top, reset, clk);

  place_251 : place
  generic map(1, 1, '0')
  port map(place_251_tip, place_251_rst, place_251_top, reset, clk);

  place_252 : place
  generic map(1, 1, '0')
  port map(place_252_tip, place_252_rst, place_252_top, reset, clk);

  place_253 : place
  generic map(1, 1, '0')
  port map(place_253_tip, place_253_rst, place_253_top, reset, clk);

  place_254 : place
  generic map(1, 1, '0')
  port map(place_254_tip, place_254_rst, place_254_top, reset, clk);

  place_255 : place
  generic map(1, 1, '0')
  port map(place_255_tip, place_255_rst, place_255_top, reset, clk);

  place_256 : place
  generic map(1, 2, '0')
  port map(place_256_tip, place_256_rst, place_256_top, reset, clk);

  place_257 : place
  generic map(1, 1, '0')
  port map(place_257_tip, place_257_rst, place_257_top, reset, clk);

  place_258 : place
  generic map(1, 1, '0')
  port map(place_258_tip, place_258_rst, place_258_top, reset, clk);

  place_259 : place
  generic map(1, 1, '0')
  port map(place_259_tip, place_259_rst, place_259_top, reset, clk);

  place_260 : place
  generic map(1, 1, '0')
  port map(place_260_tip, place_260_rst, place_260_top, reset, clk);

  place_261 : place
  generic map(1, 1, '0')
  port map(place_261_tip, place_261_rst, place_261_top, reset, clk);

  place_262 : place
  generic map(1, 1, '0')
  port map(place_262_tip, place_262_rst, place_262_top, reset, clk);

  place_263 : place
  generic map(1, 1, '0')
  port map(place_263_tip, place_263_rst, place_263_top, reset, clk);

  place_264 : place
  generic map(1, 1, '0')
  port map(place_264_tip, place_264_rst, place_264_top, reset, clk);

  place_265 : place
  generic map(1, 2, '0')
  port map(place_265_tip, place_265_rst, place_265_top, reset, clk);

  place_268 : place
  generic map(2, 1, '0')
  port map(place_268_tip, place_268_rst, place_268_top, reset, clk);

  place_269 : place
  generic map(1, 1, '0')
  port map(place_269_tip, place_269_rst, place_269_top, reset, clk);

  place_27 : place
  generic map(1, 1, '0')
  port map(place_27_tip, place_27_rst, place_27_top, reset, clk);

  place_270 : place
  generic map(1, 1, '0')
  port map(place_270_tip, place_270_rst, place_270_top, reset, clk);

  place_273 : place
  generic map(2, 1, '0')
  port map(place_273_tip, place_273_rst, place_273_top, reset, clk);

  place_274 : place
  generic map(1, 1, '0')
  port map(place_274_tip, place_274_rst, place_274_top, reset, clk);

  place_275 : place
  generic map(1, 1, '0')
  port map(place_275_tip, place_275_rst, place_275_top, reset, clk);

  place_276 : place
  generic map(1, 1, '0')
  port map(place_276_tip, place_276_rst, place_276_top, reset, clk);

  place_277 : place
  generic map(1, 1, '0')
  port map(place_277_tip, place_277_rst, place_277_top, reset, clk);

  place_278 : place
  generic map(1, 1, '0')
  port map(place_278_tip, place_278_rst, place_278_top, reset, clk);

  place_279 : place
  generic map(1, 1, '0')
  port map(place_279_tip, place_279_rst, place_279_top, reset, clk);

  place_280 : place
  generic map(1, 1, '0')
  port map(place_280_tip, place_280_rst, place_280_top, reset, clk);

  place_281 : place
  generic map(1, 1, '0')
  port map(place_281_tip, place_281_rst, place_281_top, reset, clk);

  place_282 : place
  generic map(1, 1, '0')
  port map(place_282_tip, place_282_rst, place_282_top, reset, clk);

  place_283 : place
  generic map(1, 1, '0')
  port map(place_283_tip, place_283_rst, place_283_top, reset, clk);

  place_284 : place
  generic map(1, 1, '0')
  port map(place_284_tip, place_284_rst, place_284_top, reset, clk);

  place_285 : place
  generic map(1, 1, '0')
  port map(place_285_tip, place_285_rst, place_285_top, reset, clk);

  place_286 : place
  generic map(1, 1, '0')
  port map(place_286_tip, place_286_rst, place_286_top, reset, clk);

  place_287 : place
  generic map(1, 1, '0')
  port map(place_287_tip, place_287_rst, place_287_top, reset, clk);

  place_288 : place
  generic map(1, 1, '0')
  port map(place_288_tip, place_288_rst, place_288_top, reset, clk);

  place_289 : place
  generic map(1, 1, '0')
  port map(place_289_tip, place_289_rst, place_289_top, reset, clk);

  place_290 : place
  generic map(1, 1, '0')
  port map(place_290_tip, place_290_rst, place_290_top, reset, clk);

  place_291 : place
  generic map(1, 1, '0')
  port map(place_291_tip, place_291_rst, place_291_top, reset, clk);

  place_292 : place
  generic map(1, 1, '0')
  port map(place_292_tip, place_292_rst, place_292_top, reset, clk);

  place_293 : place
  generic map(1, 1, '0')
  port map(place_293_tip, place_293_rst, place_293_top, reset, clk);

  place_294 : place
  generic map(1, 1, '0')
  port map(place_294_tip, place_294_rst, place_294_top, reset, clk);

  place_295 : place
  generic map(1, 1, '0')
  port map(place_295_tip, place_295_rst, place_295_top, reset, clk);

  place_296 : place
  generic map(1, 1, '0')
  port map(place_296_tip, place_296_rst, place_296_top, reset, clk);

  place_297 : place
  generic map(1, 1, '0')
  port map(place_297_tip, place_297_rst, place_297_top, reset, clk);

  place_298 : place
  generic map(1, 1, '0')
  port map(place_298_tip, place_298_rst, place_298_top, reset, clk);

  place_299 : place
  generic map(1, 1, '0')
  port map(place_299_tip, place_299_rst, place_299_top, reset, clk);

  place_30 : place
  generic map(1, 1, '0')
  port map(place_30_tip, place_30_rst, place_30_top, reset, clk);

  place_300 : place
  generic map(1, 1, '0')
  port map(place_300_tip, place_300_rst, place_300_top, reset, clk);

  place_301 : place
  generic map(1, 1, '0')
  port map(place_301_tip, place_301_rst, place_301_top, reset, clk);

  place_302 : place
  generic map(1, 1, '0')
  port map(place_302_tip, place_302_rst, place_302_top, reset, clk);

  place_303 : place
  generic map(1, 1, '0')
  port map(place_303_tip, place_303_rst, place_303_top, reset, clk);

  place_304 : place
  generic map(1, 1, '0')
  port map(place_304_tip, place_304_rst, place_304_top, reset, clk);

  place_305 : place
  generic map(1, 1, '0')
  port map(place_305_tip, place_305_rst, place_305_top, reset, clk);

  place_306 : place
  generic map(1, 1, '0')
  port map(place_306_tip, place_306_rst, place_306_top, reset, clk);

  place_307 : place
  generic map(1, 1, '0')
  port map(place_307_tip, place_307_rst, place_307_top, reset, clk);

  place_308 : place
  generic map(1, 1, '0')
  port map(place_308_tip, place_308_rst, place_308_top, reset, clk);

  place_309 : place
  generic map(1, 1, '0')
  port map(place_309_tip, place_309_rst, place_309_top, reset, clk);

  place_310 : place
  generic map(1, 2, '0')
  port map(place_310_tip, place_310_rst, place_310_top, reset, clk);

  place_311 : place
  generic map(1, 1, '0')
  port map(place_311_tip, place_311_rst, place_311_top, reset, clk);

  place_312 : place
  generic map(1, 1, '0')
  port map(place_312_tip, place_312_rst, place_312_top, reset, clk);

  place_313 : place
  generic map(1, 1, '0')
  port map(place_313_tip, place_313_rst, place_313_top, reset, clk);

  place_314 : place
  generic map(1, 1, '0')
  port map(place_314_tip, place_314_rst, place_314_top, reset, clk);

  place_315 : place
  generic map(1, 1, '0')
  port map(place_315_tip, place_315_rst, place_315_top, reset, clk);

  place_316 : place
  generic map(1, 1, '0')
  port map(place_316_tip, place_316_rst, place_316_top, reset, clk);

  place_317 : place
  generic map(1, 1, '0')
  port map(place_317_tip, place_317_rst, place_317_top, reset, clk);

  place_318 : place
  generic map(1, 1, '0')
  port map(place_318_tip, place_318_rst, place_318_top, reset, clk);

  place_319 : place
  generic map(1, 1, '0')
  port map(place_319_tip, place_319_rst, place_319_top, reset, clk);

  place_32 : place
  generic map(1, 1, '0')
  port map(place_32_tip, place_32_rst, place_32_top, reset, clk);

  place_320 : place
  generic map(1, 2, '0')
  port map(place_320_tip, place_320_rst, place_320_top, reset, clk);

  place_322 : place
  generic map(1, 1, '0')
  port map(place_322_tip, place_322_rst, place_322_top, reset, clk);

  place_323 : place
  generic map(2, 1, '0')
  port map(place_323_tip, place_323_rst, place_323_top, reset, clk);

  place_324 : place
  generic map(1, 1, '0')
  port map(place_324_tip, place_324_rst, place_324_top, reset, clk);

  place_325 : place
  generic map(1, 1, '0')
  port map(place_325_tip, place_325_rst, place_325_top, reset, clk);

  place_326 : place
  generic map(1, 1, '0')
  port map(place_326_tip, place_326_rst, place_326_top, reset, clk);

  place_327 : place
  generic map(2, 1, '0')
  port map(place_327_tip, place_327_rst, place_327_top, reset, clk);

  place_328 : place
  generic map(1, 1, '0')
  port map(place_328_tip, place_328_rst, place_328_top, reset, clk);

  place_329 : place
  generic map(1, 1, '0')
  port map(place_329_tip, place_329_rst, place_329_top, reset, clk);

  place_33 : place
  generic map(1, 1, '0')
  port map(place_33_tip, place_33_rst, place_33_top, reset, clk);

  place_330 : place
  generic map(1, 1, '0')
  port map(place_330_tip, place_330_rst, place_330_top, reset, clk);

  place_331 : place
  generic map(1, 1, '0')
  port map(place_331_tip, place_331_rst, place_331_top, reset, clk);

  place_332 : place
  generic map(1, 1, '0')
  port map(place_332_tip, place_332_rst, place_332_top, reset, clk);

  place_333 : place
  generic map(1, 1, '0')
  port map(place_333_tip, place_333_rst, place_333_top, reset, clk);

  place_334 : place
  generic map(1, 1, '0')
  port map(place_334_tip, place_334_rst, place_334_top, reset, clk);

  place_335 : place
  generic map(1, 1, '0')
  port map(place_335_tip, place_335_rst, place_335_top, reset, clk);

  place_336 : place
  generic map(1, 1, '0')
  port map(place_336_tip, place_336_rst, place_336_top, reset, clk);

  place_337 : place
  generic map(1, 1, '0')
  port map(place_337_tip, place_337_rst, place_337_top, reset, clk);

  place_338 : place
  generic map(1, 1, '0')
  port map(place_338_tip, place_338_rst, place_338_top, reset, clk);

  place_339 : place
  generic map(1, 1, '0')
  port map(place_339_tip, place_339_rst, place_339_top, reset, clk);

  place_340 : place
  generic map(1, 1, '0')
  port map(place_340_tip, place_340_rst, place_340_top, reset, clk);

  place_341 : place
  generic map(1, 1, '0')
  port map(place_341_tip, place_341_rst, place_341_top, reset, clk);

  place_342 : place
  generic map(1, 1, '0')
  port map(place_342_tip, place_342_rst, place_342_top, reset, clk);

  place_343 : place
  generic map(1, 1, '0')
  port map(place_343_tip, place_343_rst, place_343_top, reset, clk);

  place_344 : place
  generic map(1, 1, '0')
  port map(place_344_tip, place_344_rst, place_344_top, reset, clk);

  place_345 : place
  generic map(1, 1, '0')
  port map(place_345_tip, place_345_rst, place_345_top, reset, clk);

  place_346 : place
  generic map(1, 1, '0')
  port map(place_346_tip, place_346_rst, place_346_top, reset, clk);

  place_347 : place
  generic map(1, 1, '0')
  port map(place_347_tip, place_347_rst, place_347_top, reset, clk);

  place_349 : place
  generic map(2, 1, '0')
  port map(place_349_tip, place_349_rst, place_349_top, reset, clk);

  place_350 : place
  generic map(1, 1, '0')
  port map(place_350_tip, place_350_rst, place_350_top, reset, clk);

  place_351 : place
  generic map(1, 1, '0')
  port map(place_351_tip, place_351_rst, place_351_top, reset, clk);

  place_352 : place
  generic map(1, 1, '0')
  port map(place_352_tip, place_352_rst, place_352_top, reset, clk);

  place_354 : place
  generic map(1, 1, '0')
  port map(place_354_tip, place_354_rst, place_354_top, reset, clk);

  place_355 : place
  generic map(1, 1, '0')
  port map(place_355_tip, place_355_rst, place_355_top, reset, clk);

  place_356 : place
  generic map(1, 1, '0')
  port map(place_356_tip, place_356_rst, place_356_top, reset, clk);

  place_357 : place
  generic map(1, 1, '0')
  port map(place_357_tip, place_357_rst, place_357_top, reset, clk);

  place_358 : place
  generic map(1, 1, '0')
  port map(place_358_tip, place_358_rst, place_358_top, reset, clk);

  place_359 : place
  generic map(1, 1, '0')
  port map(place_359_tip, place_359_rst, place_359_top, reset, clk);

  place_36 : place
  generic map(1, 1, '0')
  port map(place_36_tip, place_36_rst, place_36_top, reset, clk);

  place_360 : place
  generic map(1, 1, '0')
  port map(place_360_tip, place_360_rst, place_360_top, reset, clk);

  place_361 : place
  generic map(1, 2, '0')
  port map(place_361_tip, place_361_rst, place_361_top, reset, clk);

  place_362 : place
  generic map(1, 1, '0')
  port map(place_362_tip, place_362_rst, place_362_top, reset, clk);

  place_363 : place
  generic map(1, 1, '0')
  port map(place_363_tip, place_363_rst, place_363_top, reset, clk);

  place_364 : place
  generic map(1, 1, '0')
  port map(place_364_tip, place_364_rst, place_364_top, reset, clk);

  place_365 : place
  generic map(1, 1, '0')
  port map(place_365_tip, place_365_rst, place_365_top, reset, clk);

  place_366 : place
  generic map(1, 1, '0')
  port map(place_366_tip, place_366_rst, place_366_top, reset, clk);

  place_367 : place
  generic map(1, 1, '0')
  port map(place_367_tip, place_367_rst, place_367_top, reset, clk);

  place_368 : place
  generic map(1, 1, '0')
  port map(place_368_tip, place_368_rst, place_368_top, reset, clk);

  place_369 : place
  generic map(1, 1, '0')
  port map(place_369_tip, place_369_rst, place_369_top, reset, clk);

  place_370 : place
  generic map(1, 1, '0')
  port map(place_370_tip, place_370_rst, place_370_top, reset, clk);

  place_371 : place
  generic map(1, 1, '0')
  port map(place_371_tip, place_371_rst, place_371_top, reset, clk);

  place_372 : place
  generic map(1, 1, '0')
  port map(place_372_tip, place_372_rst, place_372_top, reset, clk);

  place_373 : place
  generic map(1, 1, '0')
  port map(place_373_tip, place_373_rst, place_373_top, reset, clk);

  place_374 : place
  generic map(1, 1, '0')
  port map(place_374_tip, place_374_rst, place_374_top, reset, clk);

  place_375 : place
  generic map(1, 1, '0')
  port map(place_375_tip, place_375_rst, place_375_top, reset, clk);

  place_376 : place
  generic map(1, 1, '0')
  port map(place_376_tip, place_376_rst, place_376_top, reset, clk);

  place_377 : place
  generic map(1, 1, '0')
  port map(place_377_tip, place_377_rst, place_377_top, reset, clk);

  place_378 : place
  generic map(1, 1, '0')
  port map(place_378_tip, place_378_rst, place_378_top, reset, clk);

  place_379 : place
  generic map(1, 1, '0')
  port map(place_379_tip, place_379_rst, place_379_top, reset, clk);

  place_38 : place
  generic map(1, 1, '0')
  port map(place_38_tip, place_38_rst, place_38_top, reset, clk);

  place_380 : place
  generic map(1, 1, '0')
  port map(place_380_tip, place_380_rst, place_380_top, reset, clk);

  place_381 : place
  generic map(1, 1, '0')
  port map(place_381_tip, place_381_rst, place_381_top, reset, clk);

  place_382 : place
  generic map(1, 1, '0')
  port map(place_382_tip, place_382_rst, place_382_top, reset, clk);

  place_383 : place
  generic map(1, 1, '0')
  port map(place_383_tip, place_383_rst, place_383_top, reset, clk);

  place_384 : place
  generic map(1, 1, '0')
  port map(place_384_tip, place_384_rst, place_384_top, reset, clk);

  place_385 : place
  generic map(1, 1, '0')
  port map(place_385_tip, place_385_rst, place_385_top, reset, clk);

  place_386 : place
  generic map(1, 1, '0')
  port map(place_386_tip, place_386_rst, place_386_top, reset, clk);

  place_387 : place
  generic map(1, 1, '0')
  port map(place_387_tip, place_387_rst, place_387_top, reset, clk);

  place_388 : place
  generic map(1, 1, '0')
  port map(place_388_tip, place_388_rst, place_388_top, reset, clk);

  place_389 : place
  generic map(1, 1, '0')
  port map(place_389_tip, place_389_rst, place_389_top, reset, clk);

  place_390 : place
  generic map(1, 1, '0')
  port map(place_390_tip, place_390_rst, place_390_top, reset, clk);

  place_391 : place
  generic map(1, 2, '0')
  port map(place_391_tip, place_391_rst, place_391_top, reset, clk);

  place_392 : place
  generic map(1, 1, '0')
  port map(place_392_tip, place_392_rst, place_392_top, reset, clk);

  place_394 : place
  generic map(1, 1, '0')
  port map(place_394_tip, place_394_rst, place_394_top, reset, clk);

  place_396 : place
  generic map(1, 1, '0')
  port map(place_396_tip, place_396_rst, place_396_top, reset, clk);

  place_399 : place
  generic map(2, 1, '0')
  port map(place_399_tip, place_399_rst, place_399_top, reset, clk);

  place_40 : place
  generic map(1, 1, '0')
  port map(place_40_tip, place_40_rst, place_40_top, reset, clk);

  place_400 : place
  generic map(1, 1, '0')
  port map(place_400_tip, place_400_rst, place_400_top, reset, clk);

  place_401 : place
  generic map(1, 1, '0')
  port map(place_401_tip, place_401_rst, place_401_top, reset, clk);

  place_402 : place
  generic map(1, 1, '0')
  port map(place_402_tip, place_402_rst, place_402_top, reset, clk);

  place_403 : place
  generic map(1, 1, '0')
  port map(place_403_tip, place_403_rst, place_403_top, reset, clk);

  place_404 : place
  generic map(1, 1, '0')
  port map(place_404_tip, place_404_rst, place_404_top, reset, clk);

  place_405 : place
  generic map(1, 1, '0')
  port map(place_405_tip, place_405_rst, place_405_top, reset, clk);

  place_406 : place
  generic map(1, 1, '0')
  port map(place_406_tip, place_406_rst, place_406_top, reset, clk);

  place_407 : place
  generic map(1, 1, '0')
  port map(place_407_tip, place_407_rst, place_407_top, reset, clk);

  place_408 : place
  generic map(1, 1, '0')
  port map(place_408_tip, place_408_rst, place_408_top, reset, clk);

  place_409 : place
  generic map(1, 1, '0')
  port map(place_409_tip, place_409_rst, place_409_top, reset, clk);

  place_410 : place
  generic map(1, 1, '0')
  port map(place_410_tip, place_410_rst, place_410_top, reset, clk);

  place_411 : place
  generic map(1, 1, '0')
  port map(place_411_tip, place_411_rst, place_411_top, reset, clk);

  place_412 : place
  generic map(1, 1, '0')
  port map(place_412_tip, place_412_rst, place_412_top, reset, clk);

  place_413 : place
  generic map(1, 1, '0')
  port map(place_413_tip, place_413_rst, place_413_top, reset, clk);

  place_414 : place
  generic map(1, 1, '0')
  port map(place_414_tip, place_414_rst, place_414_top, reset, clk);

  place_415 : place
  generic map(1, 1, '0')
  port map(place_415_tip, place_415_rst, place_415_top, reset, clk);

  place_416 : place
  generic map(1, 1, '0')
  port map(place_416_tip, place_416_rst, place_416_top, reset, clk);

  place_417 : place
  generic map(1, 1, '0')
  port map(place_417_tip, place_417_rst, place_417_top, reset, clk);

  place_418 : place
  generic map(1, 1, '0')
  port map(place_418_tip, place_418_rst, place_418_top, reset, clk);

  place_419 : place
  generic map(1, 1, '0')
  port map(place_419_tip, place_419_rst, place_419_top, reset, clk);

  place_420 : place
  generic map(1, 1, '0')
  port map(place_420_tip, place_420_rst, place_420_top, reset, clk);

  place_421 : place
  generic map(1, 1, '0')
  port map(place_421_tip, place_421_rst, place_421_top, reset, clk);

  place_422 : place
  generic map(1, 1, '0')
  port map(place_422_tip, place_422_rst, place_422_top, reset, clk);

  place_423 : place
  generic map(1, 1, '0')
  port map(place_423_tip, place_423_rst, place_423_top, reset, clk);

  place_424 : place
  generic map(1, 1, '0')
  port map(place_424_tip, place_424_rst, place_424_top, reset, clk);

  place_425 : place
  generic map(1, 1, '0')
  port map(place_425_tip, place_425_rst, place_425_top, reset, clk);

  place_426 : place
  generic map(1, 1, '0')
  port map(place_426_tip, place_426_rst, place_426_top, reset, clk);

  place_427 : place
  generic map(1, 1, '0')
  port map(place_427_tip, place_427_rst, place_427_top, reset, clk);

  place_428 : place
  generic map(1, 1, '0')
  port map(place_428_tip, place_428_rst, place_428_top, reset, clk);

  place_429 : place
  generic map(1, 1, '0')
  port map(place_429_tip, place_429_rst, place_429_top, reset, clk);

  place_430 : place
  generic map(1, 1, '0')
  port map(place_430_tip, place_430_rst, place_430_top, reset, clk);

  place_431 : place
  generic map(1, 1, '0')
  port map(place_431_tip, place_431_rst, place_431_top, reset, clk);

  place_432 : place
  generic map(1, 1, '0')
  port map(place_432_tip, place_432_rst, place_432_top, reset, clk);

  place_433 : place
  generic map(1, 1, '0')
  port map(place_433_tip, place_433_rst, place_433_top, reset, clk);

  place_434 : place
  generic map(1, 1, '0')
  port map(place_434_tip, place_434_rst, place_434_top, reset, clk);

  place_435 : place
  generic map(1, 1, '0')
  port map(place_435_tip, place_435_rst, place_435_top, reset, clk);

  place_436 : place
  generic map(1, 1, '0')
  port map(place_436_tip, place_436_rst, place_436_top, reset, clk);

  place_437 : place
  generic map(1, 1, '0')
  port map(place_437_tip, place_437_rst, place_437_top, reset, clk);

  place_438 : place
  generic map(1, 1, '0')
  port map(place_438_tip, place_438_rst, place_438_top, reset, clk);

  place_439 : place
  generic map(1, 1, '0')
  port map(place_439_tip, place_439_rst, place_439_top, reset, clk);

  place_440 : place
  generic map(1, 1, '0')
  port map(place_440_tip, place_440_rst, place_440_top, reset, clk);

  place_441 : place
  generic map(1, 1, '0')
  port map(place_441_tip, place_441_rst, place_441_top, reset, clk);

  place_442 : place
  generic map(1, 1, '0')
  port map(place_442_tip, place_442_rst, place_442_top, reset, clk);

  place_443 : place
  generic map(1, 1, '0')
  port map(place_443_tip, place_443_rst, place_443_top, reset, clk);

  place_444 : place
  generic map(1, 1, '0')
  port map(place_444_tip, place_444_rst, place_444_top, reset, clk);

  place_445 : place
  generic map(1, 1, '0')
  port map(place_445_tip, place_445_rst, place_445_top, reset, clk);

  place_446 : place
  generic map(1, 1, '0')
  port map(place_446_tip, place_446_rst, place_446_top, reset, clk);

  place_447 : place
  generic map(1, 1, '0')
  port map(place_447_tip, place_447_rst, place_447_top, reset, clk);

  place_448 : place
  generic map(1, 1, '0')
  port map(place_448_tip, place_448_rst, place_448_top, reset, clk);

  place_449 : place
  generic map(1, 2, '0')
  port map(place_449_tip, place_449_rst, place_449_top, reset, clk);

  place_450 : place
  generic map(1, 1, '0')
  port map(place_450_tip, place_450_rst, place_450_top, reset, clk);

  place_451 : place
  generic map(1, 1, '0')
  port map(place_451_tip, place_451_rst, place_451_top, reset, clk);

  place_453 : place
  generic map(1, 1, '0')
  port map(place_453_tip, place_453_rst, place_453_top, reset, clk);

  place_454 : place
  generic map(1, 2, '0')
  port map(place_454_tip, place_454_rst, place_454_top, reset, clk);

  place_457 : place
  generic map(2, 1, '0')
  port map(place_457_tip, place_457_rst, place_457_top, reset, clk);

  place_458 : place
  generic map(1, 1, '0')
  port map(place_458_tip, place_458_rst, place_458_top, reset, clk);

  place_459 : place
  generic map(1, 1, '0')
  port map(place_459_tip, place_459_rst, place_459_top, reset, clk);

  place_46 : place
  generic map(2, 1, '0')
  port map(place_46_tip, place_46_rst, place_46_top, reset, clk);

  place_460 : place
  generic map(1, 1, '0')
  port map(place_460_tip, place_460_rst, place_460_top, reset, clk);

  place_462 : place
  generic map(1, 1, '0')
  port map(place_462_tip, place_462_rst, place_462_top, reset, clk);

  place_464 : place
  generic map(2, 1, '0')
  port map(place_464_tip, place_464_rst, place_464_top, reset, clk);

  place_465 : place
  generic map(1, 1, '0')
  port map(place_465_tip, place_465_rst, place_465_top, reset, clk);

  place_467 : place
  generic map(1, 1, '0')
  port map(place_467_tip, place_467_rst, place_467_top, reset, clk);

  place_469 : place
  generic map(1, 1, '0')
  port map(place_469_tip, place_469_rst, place_469_top, reset, clk);

  place_470 : place
  generic map(1, 2, '0')
  port map(place_470_tip, place_470_rst, place_470_top, reset, clk);

  place_471 : place
  generic map(1, 1, '0')
  port map(place_471_tip, place_471_rst, place_471_top, reset, clk);

  place_472 : place
  generic map(1, 1, '0')
  port map(place_472_tip, place_472_rst, place_472_top, reset, clk);

  place_473 : place
  generic map(1, 1, '0')
  port map(place_473_tip, place_473_rst, place_473_top, reset, clk);

  place_474 : place
  generic map(1, 1, '0')
  port map(place_474_tip, place_474_rst, place_474_top, reset, clk);

  place_475 : place
  generic map(1, 1, '0')
  port map(place_475_tip, place_475_rst, place_475_top, reset, clk);

  place_476 : place
  generic map(1, 1, '0')
  port map(place_476_tip, place_476_rst, place_476_top, reset, clk);

  place_477 : place
  generic map(1, 1, '0')
  port map(place_477_tip, place_477_rst, place_477_top, reset, clk);

  place_478 : place
  generic map(1, 1, '0')
  port map(place_478_tip, place_478_rst, place_478_top, reset, clk);

  place_479 : place
  generic map(1, 1, '0')
  port map(place_479_tip, place_479_rst, place_479_top, reset, clk);

  place_48 : place
  generic map(1, 1, '0')
  port map(place_48_tip, place_48_rst, place_48_top, reset, clk);

  place_480 : place
  generic map(1, 1, '0')
  port map(place_480_tip, place_480_rst, place_480_top, reset, clk);

  place_481 : place
  generic map(1, 1, '0')
  port map(place_481_tip, place_481_rst, place_481_top, reset, clk);

  place_482 : place
  generic map(1, 1, '0')
  port map(place_482_tip, place_482_rst, place_482_top, reset, clk);

  place_483 : place
  generic map(1, 1, '0')
  port map(place_483_tip, place_483_rst, place_483_top, reset, clk);

  place_484 : place
  generic map(1, 1, '0')
  port map(place_484_tip, place_484_rst, place_484_top, reset, clk);

  place_485 : place
  generic map(1, 1, '0')
  port map(place_485_tip, place_485_rst, place_485_top, reset, clk);

  place_486 : place
  generic map(1, 1, '0')
  port map(place_486_tip, place_486_rst, place_486_top, reset, clk);

  place_487 : place
  generic map(1, 1, '0')
  port map(place_487_tip, place_487_rst, place_487_top, reset, clk);

  place_488 : place
  generic map(1, 1, '0')
  port map(place_488_tip, place_488_rst, place_488_top, reset, clk);

  place_489 : place
  generic map(1, 1, '0')
  port map(place_489_tip, place_489_rst, place_489_top, reset, clk);

  place_490 : place
  generic map(1, 1, '0')
  port map(place_490_tip, place_490_rst, place_490_top, reset, clk);

  place_491 : place
  generic map(1, 1, '0')
  port map(place_491_tip, place_491_rst, place_491_top, reset, clk);

  place_492 : place
  generic map(1, 1, '0')
  port map(place_492_tip, place_492_rst, place_492_top, reset, clk);

  place_493 : place
  generic map(1, 1, '0')
  port map(place_493_tip, place_493_rst, place_493_top, reset, clk);

  place_494 : place
  generic map(1, 1, '0')
  port map(place_494_tip, place_494_rst, place_494_top, reset, clk);

  place_495 : place
  generic map(1, 1, '0')
  port map(place_495_tip, place_495_rst, place_495_top, reset, clk);

  place_496 : place
  generic map(1, 1, '0')
  port map(place_496_tip, place_496_rst, place_496_top, reset, clk);

  place_497 : place
  generic map(1, 1, '0')
  port map(place_497_tip, place_497_rst, place_497_top, reset, clk);

  place_498 : place
  generic map(1, 1, '0')
  port map(place_498_tip, place_498_rst, place_498_top, reset, clk);

  place_499 : place
  generic map(1, 1, '0')
  port map(place_499_tip, place_499_rst, place_499_top, reset, clk);

  place_5 : place
  generic map(1, 1, '0')
  port map(place_5_tip, place_5_rst, place_5_top, reset, clk);

  place_500 : place
  generic map(1, 1, '0')
  port map(place_500_tip, place_500_rst, place_500_top, reset, clk);

  place_501 : place
  generic map(1, 1, '0')
  port map(place_501_tip, place_501_rst, place_501_top, reset, clk);

  place_502 : place
  generic map(1, 1, '0')
  port map(place_502_tip, place_502_rst, place_502_top, reset, clk);

  place_503 : place
  generic map(1, 1, '0')
  port map(place_503_tip, place_503_rst, place_503_top, reset, clk);

  place_504 : place
  generic map(1, 1, '0')
  port map(place_504_tip, place_504_rst, place_504_top, reset, clk);

  place_505 : place
  generic map(1, 1, '0')
  port map(place_505_tip, place_505_rst, place_505_top, reset, clk);

  place_506 : place
  generic map(1, 1, '0')
  port map(place_506_tip, place_506_rst, place_506_top, reset, clk);

  place_507 : place
  generic map(1, 1, '0')
  port map(place_507_tip, place_507_rst, place_507_top, reset, clk);

  place_508 : place
  generic map(1, 1, '0')
  port map(place_508_tip, place_508_rst, place_508_top, reset, clk);

  place_509 : place
  generic map(1, 1, '0')
  port map(place_509_tip, place_509_rst, place_509_top, reset, clk);

  place_510 : place
  generic map(1, 1, '0')
  port map(place_510_tip, place_510_rst, place_510_top, reset, clk);

  place_511 : place
  generic map(1, 1, '0')
  port map(place_511_tip, place_511_rst, place_511_top, reset, clk);

  place_512 : place
  generic map(1, 1, '0')
  port map(place_512_tip, place_512_rst, place_512_top, reset, clk);

  place_513 : place
  generic map(1, 1, '0')
  port map(place_513_tip, place_513_rst, place_513_top, reset, clk);

  place_514 : place
  generic map(1, 2, '0')
  port map(place_514_tip, place_514_rst, place_514_top, reset, clk);

  place_515 : place
  generic map(1, 1, '0')
  port map(place_515_tip, place_515_rst, place_515_top, reset, clk);

  place_516 : place
  generic map(1, 1, '0')
  port map(place_516_tip, place_516_rst, place_516_top, reset, clk);

  place_517 : place
  generic map(2, 1, '0')
  port map(place_517_tip, place_517_rst, place_517_top, reset, clk);

  place_518 : place
  generic map(1, 1, '0')
  port map(place_518_tip, place_518_rst, place_518_top, reset, clk);

  place_519 : place
  generic map(1, 1, '0')
  port map(place_519_tip, place_519_rst, place_519_top, reset, clk);

  place_52 : place
  generic map(1, 1, '0')
  port map(place_52_tip, place_52_rst, place_52_top, reset, clk);

  place_520 : place
  generic map(2, 1, '0')
  port map(place_520_tip, place_520_rst, place_520_top, reset, clk);

  place_521 : place
  generic map(1, 1, '0')
  port map(place_521_tip, place_521_rst, place_521_top, reset, clk);

  place_522 : place
  generic map(1, 1, '0')
  port map(place_522_tip, place_522_rst, place_522_top, reset, clk);

  place_524 : place
  generic map(1, 1, '0')
  port map(place_524_tip, place_524_rst, place_524_top, reset, clk);

  place_525 : place
  generic map(1, 1, '0')
  port map(place_525_tip, place_525_rst, place_525_top, reset, clk);

  place_526 : place
  generic map(1, 1, '0')
  port map(place_526_tip, place_526_rst, place_526_top, reset, clk);

  place_527 : place
  generic map(1, 1, '0')
  port map(place_527_tip, place_527_rst, place_527_top, reset, clk);

  place_528 : place
  generic map(1, 1, '0')
  port map(place_528_tip, place_528_rst, place_528_top, reset, clk);

  place_529 : place
  generic map(1, 1, '0')
  port map(place_529_tip, place_529_rst, place_529_top, reset, clk);

  place_530 : place
  generic map(1, 1, '0')
  port map(place_530_tip, place_530_rst, place_530_top, reset, clk);

  place_531 : place
  generic map(1, 1, '0')
  port map(place_531_tip, place_531_rst, place_531_top, reset, clk);

  place_532 : place
  generic map(1, 1, '0')
  port map(place_532_tip, place_532_rst, place_532_top, reset, clk);

  place_533 : place
  generic map(1, 1, '0')
  port map(place_533_tip, place_533_rst, place_533_top, reset, clk);

  place_534 : place
  generic map(1, 1, '0')
  port map(place_534_tip, place_534_rst, place_534_top, reset, clk);

  place_535 : place
  generic map(1, 1, '0')
  port map(place_535_tip, place_535_rst, place_535_top, reset, clk);

  place_536 : place
  generic map(1, 1, '0')
  port map(place_536_tip, place_536_rst, place_536_top, reset, clk);

  place_537 : place
  generic map(1, 2, '0')
  port map(place_537_tip, place_537_rst, place_537_top, reset, clk);

  place_538 : place
  generic map(1, 1, '0')
  port map(place_538_tip, place_538_rst, place_538_top, reset, clk);

  place_539 : place
  generic map(1, 1, '0')
  port map(place_539_tip, place_539_rst, place_539_top, reset, clk);

  place_54 : place
  generic map(1, 1, '0')
  port map(place_54_tip, place_54_rst, place_54_top, reset, clk);

  place_540 : place
  generic map(1, 1, '0')
  port map(place_540_tip, place_540_rst, place_540_top, reset, clk);

  place_541 : place
  generic map(1, 1, '0')
  port map(place_541_tip, place_541_rst, place_541_top, reset, clk);

  place_542 : place
  generic map(1, 1, '0')
  port map(place_542_tip, place_542_rst, place_542_top, reset, clk);

  place_543 : place
  generic map(1, 1, '0')
  port map(place_543_tip, place_543_rst, place_543_top, reset, clk);

  place_544 : place
  generic map(1, 1, '0')
  port map(place_544_tip, place_544_rst, place_544_top, reset, clk);

  place_545 : place
  generic map(1, 1, '0')
  port map(place_545_tip, place_545_rst, place_545_top, reset, clk);

  place_546 : place
  generic map(1, 1, '0')
  port map(place_546_tip, place_546_rst, place_546_top, reset, clk);

  place_547 : place
  generic map(1, 1, '0')
  port map(place_547_tip, place_547_rst, place_547_top, reset, clk);

  place_548 : place
  generic map(1, 1, '0')
  port map(place_548_tip, place_548_rst, place_548_top, reset, clk);

  place_549 : place
  generic map(1, 1, '0')
  port map(place_549_tip, place_549_rst, place_549_top, reset, clk);

  place_550 : place
  generic map(1, 1, '0')
  port map(place_550_tip, place_550_rst, place_550_top, reset, clk);

  place_551 : place
  generic map(1, 1, '0')
  port map(place_551_tip, place_551_rst, place_551_top, reset, clk);

  place_552 : place
  generic map(1, 1, '0')
  port map(place_552_tip, place_552_rst, place_552_top, reset, clk);

  place_553 : place
  generic map(1, 1, '0')
  port map(place_553_tip, place_553_rst, place_553_top, reset, clk);

  place_554 : place
  generic map(1, 1, '0')
  port map(place_554_tip, place_554_rst, place_554_top, reset, clk);

  place_555 : place
  generic map(1, 1, '0')
  port map(place_555_tip, place_555_rst, place_555_top, reset, clk);

  place_556 : place
  generic map(1, 1, '0')
  port map(place_556_tip, place_556_rst, place_556_top, reset, clk);

  place_557 : place
  generic map(1, 1, '0')
  port map(place_557_tip, place_557_rst, place_557_top, reset, clk);

  place_558 : place
  generic map(1, 1, '0')
  port map(place_558_tip, place_558_rst, place_558_top, reset, clk);

  place_559 : place
  generic map(1, 1, '0')
  port map(place_559_tip, place_559_rst, place_559_top, reset, clk);

  place_560 : place
  generic map(1, 1, '0')
  port map(place_560_tip, place_560_rst, place_560_top, reset, clk);

  place_561 : place
  generic map(1, 1, '0')
  port map(place_561_tip, place_561_rst, place_561_top, reset, clk);

  place_562 : place
  generic map(1, 1, '0')
  port map(place_562_tip, place_562_rst, place_562_top, reset, clk);

  place_563 : place
  generic map(1, 1, '0')
  port map(place_563_tip, place_563_rst, place_563_top, reset, clk);

  place_564 : place
  generic map(1, 1, '0')
  port map(place_564_tip, place_564_rst, place_564_top, reset, clk);

  place_565 : place
  generic map(1, 1, '0')
  port map(place_565_tip, place_565_rst, place_565_top, reset, clk);

  place_566 : place
  generic map(1, 1, '0')
  port map(place_566_tip, place_566_rst, place_566_top, reset, clk);

  place_567 : place
  generic map(1, 1, '0')
  port map(place_567_tip, place_567_rst, place_567_top, reset, clk);

  place_568 : place
  generic map(1, 1, '0')
  port map(place_568_tip, place_568_rst, place_568_top, reset, clk);

  place_569 : place
  generic map(1, 1, '0')
  port map(place_569_tip, place_569_rst, place_569_top, reset, clk);

  place_570 : place
  generic map(1, 1, '0')
  port map(place_570_tip, place_570_rst, place_570_top, reset, clk);

  place_571 : place
  generic map(1, 1, '0')
  port map(place_571_tip, place_571_rst, place_571_top, reset, clk);

  place_572 : place
  generic map(1, 2, '0')
  port map(place_572_tip, place_572_rst, place_572_top, reset, clk);

  place_573 : place
  generic map(1, 1, '0')
  port map(place_573_tip, place_573_rst, place_573_top, reset, clk);

  place_574 : place
  generic map(1, 1, '0')
  port map(place_574_tip, place_574_rst, place_574_top, reset, clk);

  place_575 : place
  generic map(1, 1, '0')
  port map(place_575_tip, place_575_rst, place_575_top, reset, clk);

  place_576 : place
  generic map(1, 1, '0')
  port map(place_576_tip, place_576_rst, place_576_top, reset, clk);

  place_577 : place
  generic map(1, 1, '0')
  port map(place_577_tip, place_577_rst, place_577_top, reset, clk);

  place_578 : place
  generic map(1, 1, '0')
  port map(place_578_tip, place_578_rst, place_578_top, reset, clk);

  place_579 : place
  generic map(1, 1, '0')
  port map(place_579_tip, place_579_rst, place_579_top, reset, clk);

  place_580 : place
  generic map(1, 1, '0')
  port map(place_580_tip, place_580_rst, place_580_top, reset, clk);

  place_581 : place
  generic map(1, 1, '0')
  port map(place_581_tip, place_581_rst, place_581_top, reset, clk);

  place_582 : place
  generic map(1, 1, '0')
  port map(place_582_tip, place_582_rst, place_582_top, reset, clk);

  place_583 : place
  generic map(1, 1, '0')
  port map(place_583_tip, place_583_rst, place_583_top, reset, clk);

  place_584 : place
  generic map(1, 1, '0')
  port map(place_584_tip, place_584_rst, place_584_top, reset, clk);

  place_585 : place
  generic map(1, 1, '0')
  port map(place_585_tip, place_585_rst, place_585_top, reset, clk);

  place_586 : place
  generic map(1, 1, '0')
  port map(place_586_tip, place_586_rst, place_586_top, reset, clk);

  place_587 : place
  generic map(1, 1, '0')
  port map(place_587_tip, place_587_rst, place_587_top, reset, clk);

  place_588 : place
  generic map(1, 1, '0')
  port map(place_588_tip, place_588_rst, place_588_top, reset, clk);

  place_589 : place
  generic map(1, 1, '0')
  port map(place_589_tip, place_589_rst, place_589_top, reset, clk);

  place_59 : place
  generic map(1, 1, '0')
  port map(place_59_tip, place_59_rst, place_59_top, reset, clk);

  place_590 : place
  generic map(1, 1, '0')
  port map(place_590_tip, place_590_rst, place_590_top, reset, clk);

  place_591 : place
  generic map(1, 1, '0')
  port map(place_591_tip, place_591_rst, place_591_top, reset, clk);

  place_592 : place
  generic map(1, 1, '0')
  port map(place_592_tip, place_592_rst, place_592_top, reset, clk);

  place_593 : place
  generic map(1, 1, '0')
  port map(place_593_tip, place_593_rst, place_593_top, reset, clk);

  place_594 : place
  generic map(1, 1, '0')
  port map(place_594_tip, place_594_rst, place_594_top, reset, clk);

  place_595 : place
  generic map(1, 1, '0')
  port map(place_595_tip, place_595_rst, place_595_top, reset, clk);

  place_596 : place
  generic map(1, 1, '0')
  port map(place_596_tip, place_596_rst, place_596_top, reset, clk);

  place_597 : place
  generic map(1, 1, '0')
  port map(place_597_tip, place_597_rst, place_597_top, reset, clk);

  place_598 : place
  generic map(1, 1, '0')
  port map(place_598_tip, place_598_rst, place_598_top, reset, clk);

  place_599 : place
  generic map(1, 1, '0')
  port map(place_599_tip, place_599_rst, place_599_top, reset, clk);

  place_600 : place
  generic map(1, 1, '0')
  port map(place_600_tip, place_600_rst, place_600_top, reset, clk);

  place_601 : place
  generic map(1, 1, '0')
  port map(place_601_tip, place_601_rst, place_601_top, reset, clk);

  place_602 : place
  generic map(1, 1, '0')
  port map(place_602_tip, place_602_rst, place_602_top, reset, clk);

  place_603 : place
  generic map(1, 1, '0')
  port map(place_603_tip, place_603_rst, place_603_top, reset, clk);

  place_604 : place
  generic map(1, 1, '0')
  port map(place_604_tip, place_604_rst, place_604_top, reset, clk);

  place_605 : place
  generic map(1, 1, '0')
  port map(place_605_tip, place_605_rst, place_605_top, reset, clk);

  place_606 : place
  generic map(1, 1, '0')
  port map(place_606_tip, place_606_rst, place_606_top, reset, clk);

  place_607 : place
  generic map(1, 1, '0')
  port map(place_607_tip, place_607_rst, place_607_top, reset, clk);

  place_608 : place
  generic map(1, 2, '0')
  port map(place_608_tip, place_608_rst, place_608_top, reset, clk);

  place_609 : place
  generic map(1, 1, '0')
  port map(place_609_tip, place_609_rst, place_609_top, reset, clk);

  place_61 : place
  generic map(1, 1, '0')
  port map(place_61_tip, place_61_rst, place_61_top, reset, clk);

  place_610 : place
  generic map(1, 1, '0')
  port map(place_610_tip, place_610_rst, place_610_top, reset, clk);

  place_612 : place
  generic map(1, 1, '0')
  port map(place_612_tip, place_612_rst, place_612_top, reset, clk);

  place_613 : place
  generic map(1, 1, '0')
  port map(place_613_tip, place_613_rst, place_613_top, reset, clk);

  place_614 : place
  generic map(1, 1, '0')
  port map(place_614_tip, place_614_rst, place_614_top, reset, clk);

  place_615 : place
  generic map(1, 2, '0')
  port map(place_615_tip, place_615_rst, place_615_top, reset, clk);

  place_617 : place
  generic map(1, 1, '0')
  port map(place_617_tip, place_617_rst, place_617_top, reset, clk);

  place_618 : place
  generic map(2, 1, '0')
  port map(place_618_tip, place_618_rst, place_618_top, reset, clk);

  place_619 : place
  generic map(1, 1, '0')
  port map(place_619_tip, place_619_rst, place_619_top, reset, clk);

  place_620 : place
  generic map(1, 1, '0')
  port map(place_620_tip, place_620_rst, place_620_top, reset, clk);

  place_621 : place
  generic map(1, 1, '0')
  port map(place_621_tip, place_621_rst, place_621_top, reset, clk);

  place_622 : place
  generic map(2, 1, '0')
  port map(place_622_tip, place_622_rst, place_622_top, reset, clk);

  place_623 : place
  generic map(1, 1, '0')
  port map(place_623_tip, place_623_rst, place_623_top, reset, clk);

  place_624 : place
  generic map(1, 1, '0')
  port map(place_624_tip, place_624_rst, place_624_top, reset, clk);

  place_625 : place
  generic map(1, 1, '0')
  port map(place_625_tip, place_625_rst, place_625_top, reset, clk);

  place_626 : place
  generic map(1, 1, '0')
  port map(place_626_tip, place_626_rst, place_626_top, reset, clk);

  place_627 : place
  generic map(1, 1, '0')
  port map(place_627_tip, place_627_rst, place_627_top, reset, clk);

  place_628 : place
  generic map(1, 1, '0')
  port map(place_628_tip, place_628_rst, place_628_top, reset, clk);

  place_629 : place
  generic map(1, 1, '0')
  port map(place_629_tip, place_629_rst, place_629_top, reset, clk);

  place_63 : place
  generic map(3, 1, '0')
  port map(place_63_tip, place_63_rst, place_63_top, reset, clk);

  place_630 : place
  generic map(1, 1, '0')
  port map(place_630_tip, place_630_rst, place_630_top, reset, clk);

  place_631 : place
  generic map(1, 1, '0')
  port map(place_631_tip, place_631_rst, place_631_top, reset, clk);

  place_632 : place
  generic map(1, 2, '0')
  port map(place_632_tip, place_632_rst, place_632_top, reset, clk);

  place_635 : place
  generic map(2, 1, '0')
  port map(place_635_tip, place_635_rst, place_635_top, reset, clk);

  place_636 : place
  generic map(1, 1, '0')
  port map(place_636_tip, place_636_rst, place_636_top, reset, clk);

  place_637 : place
  generic map(1, 1, '0')
  port map(place_637_tip, place_637_rst, place_637_top, reset, clk);

  place_638 : place
  generic map(1, 1, '0')
  port map(place_638_tip, place_638_rst, place_638_top, reset, clk);

  place_639 : place
  generic map(1, 1, '0')
  port map(place_639_tip, place_639_rst, place_639_top, reset, clk);

  place_640 : place
  generic map(1, 1, '0')
  port map(place_640_tip, place_640_rst, place_640_top, reset, clk);

  place_641 : place
  generic map(1, 1, '0')
  port map(place_641_tip, place_641_rst, place_641_top, reset, clk);

  place_642 : place
  generic map(1, 1, '0')
  port map(place_642_tip, place_642_rst, place_642_top, reset, clk);

  place_643 : place
  generic map(1, 1, '0')
  port map(place_643_tip, place_643_rst, place_643_top, reset, clk);

  place_644 : place
  generic map(1, 1, '0')
  port map(place_644_tip, place_644_rst, place_644_top, reset, clk);

  place_645 : place
  generic map(1, 1, '0')
  port map(place_645_tip, place_645_rst, place_645_top, reset, clk);

  place_646 : place
  generic map(1, 1, '0')
  port map(place_646_tip, place_646_rst, place_646_top, reset, clk);

  place_647 : place
  generic map(1, 1, '0')
  port map(place_647_tip, place_647_rst, place_647_top, reset, clk);

  place_648 : place
  generic map(1, 1, '0')
  port map(place_648_tip, place_648_rst, place_648_top, reset, clk);

  place_649 : place
  generic map(1, 1, '0')
  port map(place_649_tip, place_649_rst, place_649_top, reset, clk);

  place_65 : place
  generic map(1, 1, '0')
  port map(place_65_tip, place_65_rst, place_65_top, reset, clk);

  place_650 : place
  generic map(1, 1, '0')
  port map(place_650_tip, place_650_rst, place_650_top, reset, clk);

  place_651 : place
  generic map(1, 1, '0')
  port map(place_651_tip, place_651_rst, place_651_top, reset, clk);

  place_652 : place
  generic map(1, 1, '0')
  port map(place_652_tip, place_652_rst, place_652_top, reset, clk);

  place_653 : place
  generic map(1, 1, '0')
  port map(place_653_tip, place_653_rst, place_653_top, reset, clk);

  place_654 : place
  generic map(1, 1, '0')
  port map(place_654_tip, place_654_rst, place_654_top, reset, clk);

  place_655 : place
  generic map(1, 1, '0')
  port map(place_655_tip, place_655_rst, place_655_top, reset, clk);

  place_656 : place
  generic map(1, 1, '0')
  port map(place_656_tip, place_656_rst, place_656_top, reset, clk);

  place_657 : place
  generic map(1, 1, '0')
  port map(place_657_tip, place_657_rst, place_657_top, reset, clk);

  place_658 : place
  generic map(1, 1, '0')
  port map(place_658_tip, place_658_rst, place_658_top, reset, clk);

  place_659 : place
  generic map(1, 1, '0')
  port map(place_659_tip, place_659_rst, place_659_top, reset, clk);

  place_66 : place
  generic map(1, 1, '0')
  port map(place_66_tip, place_66_rst, place_66_top, reset, clk);

  place_660 : place
  generic map(1, 1, '0')
  port map(place_660_tip, place_660_rst, place_660_top, reset, clk);

  place_661 : place
  generic map(1, 1, '0')
  port map(place_661_tip, place_661_rst, place_661_top, reset, clk);

  place_662 : place
  generic map(1, 1, '0')
  port map(place_662_tip, place_662_rst, place_662_top, reset, clk);

  place_663 : place
  generic map(1, 1, '0')
  port map(place_663_tip, place_663_rst, place_663_top, reset, clk);

  place_664 : place
  generic map(1, 1, '0')
  port map(place_664_tip, place_664_rst, place_664_top, reset, clk);

  place_665 : place
  generic map(1, 1, '0')
  port map(place_665_tip, place_665_rst, place_665_top, reset, clk);

  place_666 : place
  generic map(1, 1, '0')
  port map(place_666_tip, place_666_rst, place_666_top, reset, clk);

  place_667 : place
  generic map(1, 2, '0')
  port map(place_667_tip, place_667_rst, place_667_top, reset, clk);

  place_668 : place
  generic map(1, 1, '0')
  port map(place_668_tip, place_668_rst, place_668_top, reset, clk);

  place_669 : place
  generic map(1, 1, '0')
  port map(place_669_tip, place_669_rst, place_669_top, reset, clk);

  place_671 : place
  generic map(1, 1, '0')
  port map(place_671_tip, place_671_rst, place_671_top, reset, clk);

  place_673 : place
  generic map(2, 1, '0')
  port map(place_673_tip, place_673_rst, place_673_top, reset, clk);

  place_674 : place
  generic map(1, 1, '0')
  port map(place_674_tip, place_674_rst, place_674_top, reset, clk);

  place_675 : place
  generic map(1, 1, '0')
  port map(place_675_tip, place_675_rst, place_675_top, reset, clk);

  place_676 : place
  generic map(1, 1, '0')
  port map(place_676_tip, place_676_rst, place_676_top, reset, clk);

  place_677 : place
  generic map(1, 1, '0')
  port map(place_677_tip, place_677_rst, place_677_top, reset, clk);

  place_678 : place
  generic map(1, 1, '0')
  port map(place_678_tip, place_678_rst, place_678_top, reset, clk);

  place_679 : place
  generic map(1, 1, '0')
  port map(place_679_tip, place_679_rst, place_679_top, reset, clk);

  place_680 : place
  generic map(1, 1, '0')
  port map(place_680_tip, place_680_rst, place_680_top, reset, clk);

  place_681 : place
  generic map(1, 1, '0')
  port map(place_681_tip, place_681_rst, place_681_top, reset, clk);

  place_682 : place
  generic map(1, 2, '0')
  port map(place_682_tip, place_682_rst, place_682_top, reset, clk);

  place_684 : place
  generic map(1, 1, '0')
  port map(place_684_tip, place_684_rst, place_684_top, reset, clk);

  place_685 : place
  generic map(2, 1, '0')
  port map(place_685_tip, place_685_rst, place_685_top, reset, clk);

  place_686 : place
  generic map(1, 1, '0')
  port map(place_686_tip, place_686_rst, place_686_top, reset, clk);

  place_687 : place
  generic map(1, 1, '0')
  port map(place_687_tip, place_687_rst, place_687_top, reset, clk);

  place_688 : place
  generic map(1, 1, '0')
  port map(place_688_tip, place_688_rst, place_688_top, reset, clk);

  place_689 : place
  generic map(2, 1, '0')
  port map(place_689_tip, place_689_rst, place_689_top, reset, clk);

  place_69 : place
  generic map(1, 1, '0')
  port map(place_69_tip, place_69_rst, place_69_top, reset, clk);

  place_690 : place
  generic map(1, 1, '0')
  port map(place_690_tip, place_690_rst, place_690_top, reset, clk);

  place_691 : place
  generic map(1, 1, '0')
  port map(place_691_tip, place_691_rst, place_691_top, reset, clk);

  place_692 : place
  generic map(1, 1, '0')
  port map(place_692_tip, place_692_rst, place_692_top, reset, clk);

  place_693 : place
  generic map(1, 1, '0')
  port map(place_693_tip, place_693_rst, place_693_top, reset, clk);

  place_694 : place
  generic map(1, 1, '0')
  port map(place_694_tip, place_694_rst, place_694_top, reset, clk);

  place_695 : place
  generic map(1, 1, '0')
  port map(place_695_tip, place_695_rst, place_695_top, reset, clk);

  place_696 : place
  generic map(1, 1, '0')
  port map(place_696_tip, place_696_rst, place_696_top, reset, clk);

  place_697 : place
  generic map(1, 1, '0')
  port map(place_697_tip, place_697_rst, place_697_top, reset, clk);

  place_698 : place
  generic map(1, 2, '0')
  port map(place_698_tip, place_698_rst, place_698_top, reset, clk);

  place_7 : place
  generic map(1, 1, '0')
  port map(place_7_tip, place_7_rst, place_7_top, reset, clk);

  place_701 : place
  generic map(2, 1, '0')
  port map(place_701_tip, place_701_rst, place_701_top, reset, clk);

  place_702 : place
  generic map(1, 1, '0')
  port map(place_702_tip, place_702_rst, place_702_top, reset, clk);

  place_703 : place
  generic map(1, 1, '0')
  port map(place_703_tip, place_703_rst, place_703_top, reset, clk);

  place_704 : place
  generic map(1, 1, '0')
  port map(place_704_tip, place_704_rst, place_704_top, reset, clk);

  place_705 : place
  generic map(1, 1, '0')
  port map(place_705_tip, place_705_rst, place_705_top, reset, clk);

  place_706 : place
  generic map(1, 1, '0')
  port map(place_706_tip, place_706_rst, place_706_top, reset, clk);

  place_707 : place
  generic map(1, 1, '0')
  port map(place_707_tip, place_707_rst, place_707_top, reset, clk);

  place_708 : place
  generic map(1, 1, '0')
  port map(place_708_tip, place_708_rst, place_708_top, reset, clk);

  place_709 : place
  generic map(1, 1, '0')
  port map(place_709_tip, place_709_rst, place_709_top, reset, clk);

  place_710 : place
  generic map(1, 1, '0')
  port map(place_710_tip, place_710_rst, place_710_top, reset, clk);

  place_711 : place
  generic map(1, 1, '0')
  port map(place_711_tip, place_711_rst, place_711_top, reset, clk);

  place_712 : place
  generic map(1, 1, '0')
  port map(place_712_tip, place_712_rst, place_712_top, reset, clk);

  place_713 : place
  generic map(1, 1, '0')
  port map(place_713_tip, place_713_rst, place_713_top, reset, clk);

  place_714 : place
  generic map(1, 1, '0')
  port map(place_714_tip, place_714_rst, place_714_top, reset, clk);

  place_715 : place
  generic map(1, 1, '0')
  port map(place_715_tip, place_715_rst, place_715_top, reset, clk);

  place_716 : place
  generic map(1, 1, '0')
  port map(place_716_tip, place_716_rst, place_716_top, reset, clk);

  place_717 : place
  generic map(1, 1, '0')
  port map(place_717_tip, place_717_rst, place_717_top, reset, clk);

  place_718 : place
  generic map(1, 1, '0')
  port map(place_718_tip, place_718_rst, place_718_top, reset, clk);

  place_719 : place
  generic map(1, 1, '0')
  port map(place_719_tip, place_719_rst, place_719_top, reset, clk);

  place_72 : place
  generic map(1, 1, '0')
  port map(place_72_tip, place_72_rst, place_72_top, reset, clk);

  place_720 : place
  generic map(1, 1, '0')
  port map(place_720_tip, place_720_rst, place_720_top, reset, clk);

  place_721 : place
  generic map(1, 1, '0')
  port map(place_721_tip, place_721_rst, place_721_top, reset, clk);

  place_722 : place
  generic map(1, 1, '0')
  port map(place_722_tip, place_722_rst, place_722_top, reset, clk);

  place_723 : place
  generic map(1, 1, '0')
  port map(place_723_tip, place_723_rst, place_723_top, reset, clk);

  place_724 : place
  generic map(1, 1, '0')
  port map(place_724_tip, place_724_rst, place_724_top, reset, clk);

  place_725 : place
  generic map(1, 1, '0')
  port map(place_725_tip, place_725_rst, place_725_top, reset, clk);

  place_726 : place
  generic map(1, 1, '0')
  port map(place_726_tip, place_726_rst, place_726_top, reset, clk);

  place_727 : place
  generic map(1, 1, '0')
  port map(place_727_tip, place_727_rst, place_727_top, reset, clk);

  place_728 : place
  generic map(1, 1, '0')
  port map(place_728_tip, place_728_rst, place_728_top, reset, clk);

  place_729 : place
  generic map(1, 1, '0')
  port map(place_729_tip, place_729_rst, place_729_top, reset, clk);

  place_730 : place
  generic map(1, 1, '0')
  port map(place_730_tip, place_730_rst, place_730_top, reset, clk);

  place_731 : place
  generic map(1, 1, '0')
  port map(place_731_tip, place_731_rst, place_731_top, reset, clk);

  place_732 : place
  generic map(1, 1, '0')
  port map(place_732_tip, place_732_rst, place_732_top, reset, clk);

  place_733 : place
  generic map(1, 1, '0')
  port map(place_733_tip, place_733_rst, place_733_top, reset, clk);

  place_734 : place
  generic map(1, 1, '0')
  port map(place_734_tip, place_734_rst, place_734_top, reset, clk);

  place_735 : place
  generic map(1, 1, '0')
  port map(place_735_tip, place_735_rst, place_735_top, reset, clk);

  place_736 : place
  generic map(1, 1, '0')
  port map(place_736_tip, place_736_rst, place_736_top, reset, clk);

  place_737 : place
  generic map(1, 1, '0')
  port map(place_737_tip, place_737_rst, place_737_top, reset, clk);

  place_738 : place
  generic map(1, 2, '0')
  port map(place_738_tip, place_738_rst, place_738_top, reset, clk);

  place_739 : place
  generic map(1, 1, '0')
  port map(place_739_tip, place_739_rst, place_739_top, reset, clk);

  place_74 : place
  generic map(1, 1, '0')
  port map(place_74_tip, place_74_rst, place_74_top, reset, clk);

  place_740 : place
  generic map(1, 1, '0')
  port map(place_740_tip, place_740_rst, place_740_top, reset, clk);

  place_742 : place
  generic map(1, 1, '0')
  port map(place_742_tip, place_742_rst, place_742_top, reset, clk);

  place_744 : place
  generic map(2, 1, '0')
  port map(place_744_tip, place_744_rst, place_744_top, reset, clk);

  place_745 : place
  generic map(1, 1, '0')
  port map(place_745_tip, place_745_rst, place_745_top, reset, clk);

  place_746 : place
  generic map(1, 1, '0')
  port map(place_746_tip, place_746_rst, place_746_top, reset, clk);

  place_747 : place
  generic map(1, 1, '0')
  port map(place_747_tip, place_747_rst, place_747_top, reset, clk);

  place_748 : place
  generic map(1, 1, '0')
  port map(place_748_tip, place_748_rst, place_748_top, reset, clk);

  place_749 : place
  generic map(1, 1, '0')
  port map(place_749_tip, place_749_rst, place_749_top, reset, clk);

  place_75 : place
  generic map(1, 1, '0')
  port map(place_75_tip, place_75_rst, place_75_top, reset, clk);

  place_750 : place
  generic map(1, 1, '0')
  port map(place_750_tip, place_750_rst, place_750_top, reset, clk);

  place_751 : place
  generic map(1, 1, '0')
  port map(place_751_tip, place_751_rst, place_751_top, reset, clk);

  place_752 : place
  generic map(1, 1, '0')
  port map(place_752_tip, place_752_rst, place_752_top, reset, clk);

  place_753 : place
  generic map(1, 2, '0')
  port map(place_753_tip, place_753_rst, place_753_top, reset, clk);

  place_77 : place
  generic map(1, 1, '0')
  port map(place_77_tip, place_77_rst, place_77_top, reset, clk);

  place_81 : place
  generic map(1, 1, '0')
  port map(place_81_tip, place_81_rst, place_81_top, reset, clk);

  place_83 : place
  generic map(1, 1, '0')
  port map(place_83_tip, place_83_rst, place_83_top, reset, clk);

  place_84 : place
  generic map(1, 1, '1')
  port map(place_84_tip, place_84_rst, place_84_top, reset, clk);

  place_86 : place
  generic map(1, 1, '0')
  port map(place_86_tip, place_86_rst, place_86_top, reset, clk);

  place_87 : place
  generic map(1, 1, '0')
  port map(place_87_tip, place_87_rst, place_87_top, reset, clk);

  place_88 : place
  generic map(1, 1, '0')
  port map(place_88_tip, place_88_rst, place_88_top, reset, clk);

  place_89 : place
  generic map(1, 1, '0')
  port map(place_89_tip, place_89_rst, place_89_top, reset, clk);

  place_9 : place
  generic map(1, 1, '0')
  port map(place_9_tip, place_9_rst, place_9_top, reset, clk);

  place_90 : place
  generic map(1, 1, '0')
  port map(place_90_tip, place_90_rst, place_90_top, reset, clk);

  place_91 : place
  generic map(1, 1, '0')
  port map(place_91_tip, place_91_rst, place_91_top, reset, clk);

  place_92 : place
  generic map(1, 1, '0')
  port map(place_92_tip, place_92_rst, place_92_top, reset, clk);

  place_93 : place
  generic map(1, 1, '0')
  port map(place_93_tip, place_93_rst, place_93_top, reset, clk);

  place_94 : place
  generic map(1, 1, '0')
  port map(place_94_tip, place_94_rst, place_94_top, reset, clk);

  place_95 : place
  generic map(1, 1, '0')
  port map(place_95_tip, place_95_rst, place_95_top, reset, clk);

  place_96 : place
  generic map(1, 1, '0')
  port map(place_96_tip, place_96_rst, place_96_top, reset, clk);

  place_97 : place
  generic map(1, 1, '0')
  port map(place_97_tip, place_97_rst, place_97_top, reset, clk);

  place_99 : place
  generic map(1, 1, '0')
  port map(place_99_tip, place_99_rst, place_99_top, reset, clk);


  cbr_10_oper_tmp_d_42_bool_d_req : transition
  generic map(2)
  port map(cbr_10_oper_tmp_d_42_bool_d_req_tip, cbr_10_oper_tmp_d_42_bool_d_req_ge, cbr_10_oper_tmp_d_42_bool_d_req_top);

  cbr_11_oper_tmp_d_54_bool_d_req : transition
  generic map(3)
  port map(cbr_11_oper_tmp_d_54_bool_d_req_tip, cbr_11_oper_tmp_d_54_bool_d_req_ge, cbr_11_oper_tmp_d_54_bool_d_req_top);

  cbr_12_oper_tmp_d_4223_bool_d_req : transition
  generic map(2)
  port map(cbr_12_oper_tmp_d_4223_bool_d_req_tip, cbr_12_oper_tmp_d_4223_bool_d_req_ge, cbr_12_oper_tmp_d_4223_bool_d_req_top);

  cbr_13_oper_exitcond128_bool_d_req : transition
  generic map(4)
  port map(cbr_13_oper_exitcond128_bool_d_req_tip, cbr_13_oper_exitcond128_bool_d_req_ge, cbr_13_oper_exitcond128_bool_d_req_top);

  cbr_14_oper_exitcond131_bool_d_req : transition
  generic map(2)
  port map(cbr_14_oper_exitcond131_bool_d_req_tip, cbr_14_oper_exitcond131_bool_d_req_ge, cbr_14_oper_exitcond131_bool_d_req_top);

  cbr_15_oper_tmp_d_92_bool_d_req : transition
  generic map(1)
  port map(cbr_15_oper_tmp_d_92_bool_d_req_tip, cbr_15_oper_tmp_d_92_bool_d_req_ge, cbr_15_oper_tmp_d_92_bool_d_req_top);

  cbr_16_oper_tmp_d_11348_bool_d_req : transition
  generic map(3)
  port map(cbr_16_oper_tmp_d_11348_bool_d_req_tip, cbr_16_oper_tmp_d_11348_bool_d_req_ge, cbr_16_oper_tmp_d_11348_bool_d_req_top);

  cbr_17_oper_tmp_d_113_bool_d_req : transition
  generic map(4)
  port map(cbr_17_oper_tmp_d_113_bool_d_req_tip, cbr_17_oper_tmp_d_113_bool_d_req_ge, cbr_17_oper_tmp_d_113_bool_d_req_top);

  cbr_18_oper_exitcond142_bool_d_req : transition
  generic map(1)
  port map(cbr_18_oper_exitcond142_bool_d_req_tip, cbr_18_oper_exitcond142_bool_d_req_ge, cbr_18_oper_exitcond142_bool_d_req_top);

  cbr_19_oper_tmp_d_149_bool_d_req : transition
  generic map(1)
  port map(cbr_19_oper_tmp_d_149_bool_d_req_tip, cbr_19_oper_tmp_d_149_bool_d_req_ge, cbr_19_oper_tmp_d_149_bool_d_req_top);

  cbr_20_oper_tmp_d_14574_bool_d_req : transition
  generic map(4)
  port map(cbr_20_oper_tmp_d_14574_bool_d_req_tip, cbr_20_oper_tmp_d_14574_bool_d_req_ge, cbr_20_oper_tmp_d_14574_bool_d_req_top);

  cbr_21_oper_tmp_d_166_bool_d_req : transition
  generic map(2)
  port map(cbr_21_oper_tmp_d_166_bool_d_req_tip, cbr_21_oper_tmp_d_166_bool_d_req_ge, cbr_21_oper_tmp_d_166_bool_d_req_top);

  cbr_22_oper_tmp_d_14578_bool_d_req : transition
  generic map(4)
  port map(cbr_22_oper_tmp_d_14578_bool_d_req_tip, cbr_22_oper_tmp_d_14578_bool_d_req_ge, cbr_22_oper_tmp_d_14578_bool_d_req_top);

  cbr_23_oper_tmp_d_14580_bool_d_req : transition
  generic map(4)
  port map(cbr_23_oper_tmp_d_14580_bool_d_req_tip, cbr_23_oper_tmp_d_14580_bool_d_req_ge, cbr_23_oper_tmp_d_14580_bool_d_req_top);

  cbr_24_oper_exitcond145_bool_d_req : transition
  generic map(1)
  port map(cbr_24_oper_exitcond145_bool_d_req_tip, cbr_24_oper_exitcond145_bool_d_req_ge, cbr_24_oper_exitcond145_bool_d_req_top);

  cbr_25_oper_tmp_d_202_bool_d_req : transition
  generic map(3)
  port map(cbr_25_oper_tmp_d_202_bool_d_req_tip, cbr_25_oper_tmp_d_202_bool_d_req_ge, cbr_25_oper_tmp_d_202_bool_d_req_top);

  cbr_26_oper_tmp_d_20299_bool_d_req : transition
  generic map(4)
  port map(cbr_26_oper_tmp_d_20299_bool_d_req_tip, cbr_26_oper_tmp_d_20299_bool_d_req_ge, cbr_26_oper_tmp_d_20299_bool_d_req_top);

  cbr_27_oper_exitcond150_bool_d_req : transition
  generic map(2)
  port map(cbr_27_oper_exitcond150_bool_d_req_tip, cbr_27_oper_exitcond150_bool_d_req_ge, cbr_27_oper_exitcond150_bool_d_req_top);

  cbr_28_oper_tmp_d_221_bool_d_req : transition
  generic map(2)
  port map(cbr_28_oper_tmp_d_221_bool_d_req_tip, cbr_28_oper_tmp_d_221_bool_d_req_ge, cbr_28_oper_tmp_d_221_bool_d_req_top);

  cbr_29_oper_tmp_d_221111_bool_d_req : transition
  generic map(4)
  port map(cbr_29_oper_tmp_d_221111_bool_d_req_tip, cbr_29_oper_tmp_d_221111_bool_d_req_ge, cbr_29_oper_tmp_d_221111_bool_d_req_top);

  cbr_30_oper_exitcond158_bool_d_req : transition
  generic map(2)
  port map(cbr_30_oper_exitcond158_bool_d_req_tip, cbr_30_oper_exitcond158_bool_d_req_ge, cbr_30_oper_exitcond158_bool_d_req_top);

  cbr_6_oper_exitcond_bool_d_req : transition
  generic map(3)
  port map(cbr_6_oper_exitcond_bool_d_req_tip, cbr_6_oper_exitcond_bool_d_req_ge, cbr_6_oper_exitcond_bool_d_req_top);

  cbr_7_oper_exitcond120_bool_d_req : transition
  generic map(1)
  port map(cbr_7_oper_exitcond120_bool_d_req_tip, cbr_7_oper_exitcond120_bool_d_req_ge, cbr_7_oper_exitcond120_bool_d_req_top);

  cbr_8_oper_tmp_d_16_bool_d_req : transition
  generic map(1)
  port map(cbr_8_oper_tmp_d_16_bool_d_req_tip, cbr_8_oper_tmp_d_16_bool_d_req_ge, cbr_8_oper_tmp_d_16_bool_d_req_top);

  cbr_9_oper_tmp_d_1614_bool_d_req : transition
  generic map(4)
  port map(cbr_9_oper_tmp_d_1614_bool_d_req_tip, cbr_9_oper_tmp_d_1614_bool_d_req_ge, cbr_9_oper_tmp_d_1614_bool_d_req_top);

  else_d_0_d_entry : transition
  generic map(1)
  port map(else_d_0_d_entry_tip, else_d_0_d_entry_ge, else_d_0_d_entry_top);

  else_d_0_to_else_d_1_src : transition
  generic map(1)
  port map(else_d_0_to_else_d_1_src_tip, else_d_0_to_else_d_1_src_ge, else_d_0_to_else_d_1_src_top);

  else_d_0_to_then_d_2_src : transition
  generic map(1)
  port map(else_d_0_to_then_d_2_src_tip, else_d_0_to_then_d_2_src_ge, else_d_0_to_then_d_2_src_top);

  else_d_1_d_entry : transition
  generic map(1)
  port map(else_d_1_d_entry_tip, else_d_1_d_entry_ge, else_d_1_d_entry_top);

  else_d_1_to_loopexit_d_10_src : transition
  generic map(1)
  port map(else_d_1_to_loopexit_d_10_src_tip, else_d_1_to_loopexit_d_10_src_ge, else_d_1_to_loopexit_d_10_src_top);

  else_d_1_to_no_exit_d_10_d_backedge_src : transition
  generic map(1)
  port map(else_d_1_to_no_exit_d_10_d_backedge_src_tip, else_d_1_to_no_exit_d_10_d_backedge_src_ge, else_d_1_to_no_exit_d_10_d_backedge_src_top);

  fin : transition
  generic map(1)
  port map(fin_tip, fin_ge, fin_top);

  indvar118_d_ph_d_ph_mux_1_d_ack : transition
  generic map(1)
  port map(indvar118_d_ph_d_ph_mux_1_d_ack_tip, indvar118_d_ph_d_ph_mux_1_d_ack_ge, indvar118_d_ph_d_ph_mux_1_d_ack_top);

  indvar118_d_ph_d_ph_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar118_d_ph_d_ph_mux_1_d_req0_tip, indvar118_d_ph_d_ph_mux_1_d_req0_ge, indvar118_d_ph_d_ph_mux_1_d_req0_top);

  indvar118_d_ph_d_ph_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar118_d_ph_d_ph_mux_1_d_req1_tip, indvar118_d_ph_d_ph_mux_1_d_req1_ge, indvar118_d_ph_d_ph_mux_1_d_req1_top);

  indvar121_mux_1_d_ack : transition
  generic map(1)
  port map(indvar121_mux_1_d_ack_tip, indvar121_mux_1_d_ack_ge, indvar121_mux_1_d_ack_top);

  indvar121_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar121_mux_1_d_req0_tip, indvar121_mux_1_d_req0_ge, indvar121_mux_1_d_req0_top);

  indvar121_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar121_mux_1_d_req1_tip, indvar121_mux_1_d_req1_ge, indvar121_mux_1_d_req1_top);

  indvar123_mux_1_d_ack : transition
  generic map(1)
  port map(indvar123_mux_1_d_ack_tip, indvar123_mux_1_d_ack_ge, indvar123_mux_1_d_ack_top);

  indvar123_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar123_mux_1_d_req0_tip, indvar123_mux_1_d_req0_ge, indvar123_mux_1_d_req0_top);

  indvar123_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar123_mux_1_d_req1_tip, indvar123_mux_1_d_req1_ge, indvar123_mux_1_d_req1_top);

  indvar126_mux_1_d_ack : transition
  generic map(1)
  port map(indvar126_mux_1_d_ack_tip, indvar126_mux_1_d_ack_ge, indvar126_mux_1_d_ack_top);

  indvar126_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar126_mux_1_d_req0_tip, indvar126_mux_1_d_req0_ge, indvar126_mux_1_d_req0_top);

  indvar126_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar126_mux_1_d_req1_tip, indvar126_mux_1_d_req1_ge, indvar126_mux_1_d_req1_top);

  indvar129_mux_1_d_ack : transition
  generic map(1)
  port map(indvar129_mux_1_d_ack_tip, indvar129_mux_1_d_ack_ge, indvar129_mux_1_d_ack_top);

  indvar129_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar129_mux_1_d_req0_tip, indvar129_mux_1_d_req0_ge, indvar129_mux_1_d_req0_top);

  indvar129_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar129_mux_1_d_req1_tip, indvar129_mux_1_d_req1_ge, indvar129_mux_1_d_req1_top);

  indvar132_mux_1_d_ack : transition
  generic map(1)
  port map(indvar132_mux_1_d_ack_tip, indvar132_mux_1_d_ack_ge, indvar132_mux_1_d_ack_top);

  indvar132_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar132_mux_1_d_req0_tip, indvar132_mux_1_d_req0_ge, indvar132_mux_1_d_req0_top);

  indvar132_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar132_mux_1_d_req1_tip, indvar132_mux_1_d_req1_ge, indvar132_mux_1_d_req1_top);

  indvar134_mux_1_d_ack : transition
  generic map(1)
  port map(indvar134_mux_1_d_ack_tip, indvar134_mux_1_d_ack_ge, indvar134_mux_1_d_ack_top);

  indvar134_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar134_mux_1_d_req0_tip, indvar134_mux_1_d_req0_ge, indvar134_mux_1_d_req0_top);

  indvar134_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar134_mux_1_d_req1_tip, indvar134_mux_1_d_req1_ge, indvar134_mux_1_d_req1_top);

  indvar138_mux_1_d_ack : transition
  generic map(1)
  port map(indvar138_mux_1_d_ack_tip, indvar138_mux_1_d_ack_ge, indvar138_mux_1_d_ack_top);

  indvar138_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar138_mux_1_d_req0_tip, indvar138_mux_1_d_req0_ge, indvar138_mux_1_d_req0_top);

  indvar138_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar138_mux_1_d_req1_tip, indvar138_mux_1_d_req1_ge, indvar138_mux_1_d_req1_top);

  indvar143_mux_1_d_ack : transition
  generic map(1)
  port map(indvar143_mux_1_d_ack_tip, indvar143_mux_1_d_ack_ge, indvar143_mux_1_d_ack_top);

  indvar143_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar143_mux_1_d_req0_tip, indvar143_mux_1_d_req0_ge, indvar143_mux_1_d_req0_top);

  indvar143_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar143_mux_1_d_req1_tip, indvar143_mux_1_d_req1_ge, indvar143_mux_1_d_req1_top);

  indvar146_mux_1_d_ack : transition
  generic map(1)
  port map(indvar146_mux_1_d_ack_tip, indvar146_mux_1_d_ack_ge, indvar146_mux_1_d_ack_top);

  indvar146_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar146_mux_1_d_req0_tip, indvar146_mux_1_d_req0_ge, indvar146_mux_1_d_req0_top);

  indvar146_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar146_mux_1_d_req1_tip, indvar146_mux_1_d_req1_ge, indvar146_mux_1_d_req1_top);

  indvar148_mux_1_d_ack : transition
  generic map(1)
  port map(indvar148_mux_1_d_ack_tip, indvar148_mux_1_d_ack_ge, indvar148_mux_1_d_ack_top);

  indvar148_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar148_mux_1_d_req0_tip, indvar148_mux_1_d_req0_ge, indvar148_mux_1_d_req0_top);

  indvar148_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar148_mux_1_d_req1_tip, indvar148_mux_1_d_req1_ge, indvar148_mux_1_d_req1_top);

  indvar151_mux_1_d_ack : transition
  generic map(1)
  port map(indvar151_mux_1_d_ack_tip, indvar151_mux_1_d_ack_ge, indvar151_mux_1_d_ack_top);

  indvar151_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar151_mux_1_d_req0_tip, indvar151_mux_1_d_req0_ge, indvar151_mux_1_d_req0_top);

  indvar151_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar151_mux_1_d_req1_tip, indvar151_mux_1_d_req1_ge, indvar151_mux_1_d_req1_top);

  indvar153_mux_1_d_ack : transition
  generic map(1)
  port map(indvar153_mux_1_d_ack_tip, indvar153_mux_1_d_ack_ge, indvar153_mux_1_d_ack_top);

  indvar153_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar153_mux_1_d_req0_tip, indvar153_mux_1_d_req0_ge, indvar153_mux_1_d_req0_top);

  indvar153_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar153_mux_1_d_req1_tip, indvar153_mux_1_d_req1_ge, indvar153_mux_1_d_req1_top);

  indvar_mux_1_d_ack : transition
  generic map(1)
  port map(indvar_mux_1_d_ack_tip, indvar_mux_1_d_ack_ge, indvar_mux_1_d_ack_top);

  indvar_mux_1_d_req0 : transition
  generic map(1)
  port map(indvar_mux_1_d_req0_tip, indvar_mux_1_d_req0_ge, indvar_mux_1_d_req0_top);

  indvar_mux_1_d_req1 : transition
  generic map(1)
  port map(indvar_mux_1_d_req1_tip, indvar_mux_1_d_req1_ge, indvar_mux_1_d_req1_top);

  init : transition
  generic map(1)
  port map(init_tip, init_ge, init_top);

  j_d_3_d_in_d_ph_mux_1_d_ack : transition
  generic map(1)
  port map(j_d_3_d_in_d_ph_mux_1_d_ack_tip, j_d_3_d_in_d_ph_mux_1_d_ack_ge, j_d_3_d_in_d_ph_mux_1_d_ack_top);

  j_d_3_d_in_d_ph_mux_1_d_req0 : transition
  generic map(1)
  port map(j_d_3_d_in_d_ph_mux_1_d_req0_tip, j_d_3_d_in_d_ph_mux_1_d_req0_ge, j_d_3_d_in_d_ph_mux_1_d_req0_top);

  j_d_3_d_in_d_ph_mux_1_d_req1 : transition
  generic map(1)
  port map(j_d_3_d_in_d_ph_mux_1_d_req1_tip, j_d_3_d_in_d_ph_mux_1_d_req1_ge, j_d_3_d_in_d_ph_mux_1_d_req1_top);

  j_d_3_d_in_mux_1_d_ack : transition
  generic map(1)
  port map(j_d_3_d_in_mux_1_d_ack_tip, j_d_3_d_in_mux_1_d_ack_ge, j_d_3_d_in_mux_1_d_ack_top);

  j_d_3_d_in_mux_1_d_req0 : transition
  generic map(1)
  port map(j_d_3_d_in_mux_1_d_req0_tip, j_d_3_d_in_mux_1_d_req0_ge, j_d_3_d_in_mux_1_d_req0_top);

  j_d_3_d_in_mux_1_d_req1 : transition
  generic map(1)
  port map(j_d_3_d_in_mux_1_d_req1_tip, j_d_3_d_in_mux_1_d_req1_ge, j_d_3_d_in_mux_1_d_req1_top);

  j_d_9_d_2_d_be_mux_1_d_ack : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_1_d_ack_tip, j_d_9_d_2_d_be_mux_1_d_ack_ge, j_d_9_d_2_d_be_mux_1_d_ack_top);

  j_d_9_d_2_d_be_mux_1_d_req0 : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_1_d_req0_tip, j_d_9_d_2_d_be_mux_1_d_req0_ge, j_d_9_d_2_d_be_mux_1_d_req0_top);

  j_d_9_d_2_d_be_mux_1_d_req1 : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_1_d_req1_tip, j_d_9_d_2_d_be_mux_1_d_req1_ge, j_d_9_d_2_d_be_mux_1_d_req1_top);

  j_d_9_d_2_d_be_mux_2_d_ack : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_2_d_ack_tip, j_d_9_d_2_d_be_mux_2_d_ack_ge, j_d_9_d_2_d_be_mux_2_d_ack_top);

  j_d_9_d_2_d_be_mux_2_d_req0 : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_2_d_req0_tip, j_d_9_d_2_d_be_mux_2_d_req0_ge, j_d_9_d_2_d_be_mux_2_d_req0_top);

  j_d_9_d_2_d_be_mux_2_d_req1 : transition
  generic map(1)
  port map(j_d_9_d_2_d_be_mux_2_d_req1_tip, j_d_9_d_2_d_be_mux_2_d_req1_ge, j_d_9_d_2_d_be_mux_2_d_req1_top);

  j_d_9_d_2_mux_1_d_ack : transition
  generic map(1)
  port map(j_d_9_d_2_mux_1_d_ack_tip, j_d_9_d_2_mux_1_d_ack_ge, j_d_9_d_2_mux_1_d_ack_top);

  j_d_9_d_2_mux_1_d_req0 : transition
  generic map(1)
  port map(j_d_9_d_2_mux_1_d_req0_tip, j_d_9_d_2_mux_1_d_req0_ge, j_d_9_d_2_mux_1_d_req0_top);

  j_d_9_d_2_mux_1_d_req1 : transition
  generic map(1)
  port map(j_d_9_d_2_mux_1_d_req1_tip, j_d_9_d_2_mux_1_d_req1_ge, j_d_9_d_2_mux_1_d_req1_top);

  k_d_1_d_in_d_ph_mux_1_d_ack : transition
  generic map(1)
  port map(k_d_1_d_in_d_ph_mux_1_d_ack_tip, k_d_1_d_in_d_ph_mux_1_d_ack_ge, k_d_1_d_in_d_ph_mux_1_d_ack_top);

  k_d_1_d_in_d_ph_mux_1_d_req0 : transition
  generic map(1)
  port map(k_d_1_d_in_d_ph_mux_1_d_req0_tip, k_d_1_d_in_d_ph_mux_1_d_req0_ge, k_d_1_d_in_d_ph_mux_1_d_req0_top);

  k_d_1_d_in_d_ph_mux_1_d_req1 : transition
  generic map(1)
  port map(k_d_1_d_in_d_ph_mux_1_d_req1_tip, k_d_1_d_in_d_ph_mux_1_d_req1_ge, k_d_1_d_in_d_ph_mux_1_d_req1_top);

  k_d_2_d_3_mux_1_d_ack : transition
  generic map(1)
  port map(k_d_2_d_3_mux_1_d_ack_tip, k_d_2_d_3_mux_1_d_ack_ge, k_d_2_d_3_mux_1_d_ack_top);

  k_d_2_d_3_mux_1_d_req0 : transition
  generic map(1)
  port map(k_d_2_d_3_mux_1_d_req0_tip, k_d_2_d_3_mux_1_d_req0_ge, k_d_2_d_3_mux_1_d_req0_top);

  k_d_2_d_3_mux_1_d_req1 : transition
  generic map(1)
  port map(k_d_2_d_3_mux_1_d_req1_tip, k_d_2_d_3_mux_1_d_req1_ge, k_d_2_d_3_mux_1_d_req1_top);

  k_d_3_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(k_d_3_d_0_mux_1_d_ack_tip, k_d_3_d_0_mux_1_d_ack_ge, k_d_3_d_0_mux_1_d_ack_top);

  k_d_3_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(k_d_3_d_0_mux_1_d_req0_tip, k_d_3_d_0_mux_1_d_req0_ge, k_d_3_d_0_mux_1_d_req0_top);

  k_d_3_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(k_d_3_d_0_mux_1_d_req1_tip, k_d_3_d_0_mux_1_d_req1_ge, k_d_3_d_0_mux_1_d_req1_top);

  k_d_4_d_3_mux_1_d_ack : transition
  generic map(1)
  port map(k_d_4_d_3_mux_1_d_ack_tip, k_d_4_d_3_mux_1_d_ack_ge, k_d_4_d_3_mux_1_d_ack_top);

  k_d_4_d_3_mux_1_d_req0 : transition
  generic map(1)
  port map(k_d_4_d_3_mux_1_d_req0_tip, k_d_4_d_3_mux_1_d_req0_ge, k_d_4_d_3_mux_1_d_req0_top);

  k_d_4_d_3_mux_1_d_req1 : transition
  generic map(1)
  port map(k_d_4_d_3_mux_1_d_req1_tip, k_d_4_d_3_mux_1_d_req1_ge, k_d_4_d_3_mux_1_d_req1_top);

  k_d_5_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(k_d_5_d_0_mux_1_d_ack_tip, k_d_5_d_0_mux_1_d_ack_ge, k_d_5_d_0_mux_1_d_ack_top);

  k_d_5_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(k_d_5_d_0_mux_1_d_req0_tip, k_d_5_d_0_mux_1_d_req0_ge, k_d_5_d_0_mux_1_d_req0_top);

  k_d_5_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(k_d_5_d_0_mux_1_d_req1_tip, k_d_5_d_0_mux_1_d_req1_ge, k_d_5_d_0_mux_1_d_req1_top);

  load_A_d_ack : transition
  generic map(1)
  port map(load_A_d_ack_tip, load_A_d_ack_ge, load_A_d_ack_top);

  load_A_d_req : transition
  generic map(1)
  port map(load_A_d_req_tip, load_A_d_req_ge, load_A_d_req_top);

  load_ccoeff_d_ack : transition
  generic map(1)
  port map(load_ccoeff_d_ack_tip, load_ccoeff_d_ack_ge, load_ccoeff_d_ack_top);

  load_ccoeff_d_req : transition
  generic map(1)
  port map(load_ccoeff_d_req_tip, load_ccoeff_d_req_ge, load_ccoeff_d_req_top);

  load_l_array_d_ack : transition
  generic map(1)
  port map(load_l_array_d_ack_tip, load_l_array_d_ack_ge, load_l_array_d_ack_top);

  load_l_array_d_req : transition
  generic map(1)
  port map(load_l_array_d_req_tip, load_l_array_d_req_ge, load_l_array_d_req_top);

  load_noofelem_d_ack : transition
  generic map(1)
  port map(load_noofelem_d_ack_tip, load_noofelem_d_ack_ge, load_noofelem_d_ack_top);

  load_noofelem_d_req : transition
  generic map(1)
  port map(load_noofelem_d_req_tip, load_noofelem_d_req_ge, load_noofelem_d_req_top);

  load_rcoeff_d_ack : transition
  generic map(1)
  port map(load_rcoeff_d_ack_tip, load_rcoeff_d_ack_ge, load_rcoeff_d_ack_top);

  load_rcoeff_d_req : transition
  generic map(1)
  port map(load_rcoeff_d_req_tip, load_rcoeff_d_req_ge, load_rcoeff_d_req_top);

  load_start_call_divide_0_return_d_ack : transition
  generic map(1)
  port map(load_start_call_divide_0_return_d_ack_tip, load_start_call_divide_0_return_d_ack_ge, load_start_call_divide_0_return_d_ack_top);

  load_start_call_divide_0_return_d_req : transition
  generic map(1)
  port map(load_start_call_divide_0_return_d_req_tip, load_start_call_divide_0_return_d_req_ge, load_start_call_divide_0_return_d_req_top);

  load_tmp_d_103_d_ack : transition
  generic map(1)
  port map(load_tmp_d_103_d_ack_tip, load_tmp_d_103_d_ack_ge, load_tmp_d_103_d_ack_top);

  load_tmp_d_103_d_req : transition
  generic map(1)
  port map(load_tmp_d_103_d_req_tip, load_tmp_d_103_d_req_ge, load_tmp_d_103_d_req_top);

  load_tmp_d_108_d_ack : transition
  generic map(1)
  port map(load_tmp_d_108_d_ack_tip, load_tmp_d_108_d_ack_ge, load_tmp_d_108_d_ack_top);

  load_tmp_d_108_d_req : transition
  generic map(2)
  port map(load_tmp_d_108_d_req_tip, load_tmp_d_108_d_req_ge, load_tmp_d_108_d_req_top);

  load_tmp_d_123_d_ack : transition
  generic map(1)
  port map(load_tmp_d_123_d_ack_tip, load_tmp_d_123_d_ack_ge, load_tmp_d_123_d_ack_top);

  load_tmp_d_123_d_req : transition
  generic map(1)
  port map(load_tmp_d_123_d_req_tip, load_tmp_d_123_d_req_ge, load_tmp_d_123_d_req_top);

  load_tmp_d_128_d_ack : transition
  generic map(1)
  port map(load_tmp_d_128_d_ack_tip, load_tmp_d_128_d_ack_ge, load_tmp_d_128_d_ack_top);

  load_tmp_d_128_d_req : transition
  generic map(2)
  port map(load_tmp_d_128_d_req_tip, load_tmp_d_128_d_req_ge, load_tmp_d_128_d_req_top);

  load_tmp_d_133_d_ack : transition
  generic map(1)
  port map(load_tmp_d_133_d_ack_tip, load_tmp_d_133_d_ack_ge, load_tmp_d_133_d_ack_top);

  load_tmp_d_133_d_req : transition
  generic map(2)
  port map(load_tmp_d_133_d_req_tip, load_tmp_d_133_d_req_ge, load_tmp_d_133_d_req_top);

  load_tmp_d_159_d_ack : transition
  generic map(1)
  port map(load_tmp_d_159_d_ack_tip, load_tmp_d_159_d_ack_ge, load_tmp_d_159_d_ack_top);

  load_tmp_d_159_d_req : transition
  generic map(1)
  port map(load_tmp_d_159_d_req_tip, load_tmp_d_159_d_req_ge, load_tmp_d_159_d_req_top);

  load_tmp_d_180_d_ack : transition
  generic map(1)
  port map(load_tmp_d_180_d_ack_tip, load_tmp_d_180_d_ack_ge, load_tmp_d_180_d_ack_top);

  load_tmp_d_180_d_req : transition
  generic map(2)
  port map(load_tmp_d_180_d_req_tip, load_tmp_d_180_d_req_ge, load_tmp_d_180_d_req_top);

  load_tmp_d_193_d_ack : transition
  generic map(1)
  port map(load_tmp_d_193_d_ack_tip, load_tmp_d_193_d_ack_ge, load_tmp_d_193_d_ack_top);

  load_tmp_d_193_d_req : transition
  generic map(2)
  port map(load_tmp_d_193_d_req_tip, load_tmp_d_193_d_req_ge, load_tmp_d_193_d_req_top);

  load_tmp_d_211_d_ack : transition
  generic map(1)
  port map(load_tmp_d_211_d_ack_tip, load_tmp_d_211_d_ack_ge, load_tmp_d_211_d_ack_top);

  load_tmp_d_211_d_req : transition
  generic map(1)
  port map(load_tmp_d_211_d_req_tip, load_tmp_d_211_d_req_ge, load_tmp_d_211_d_req_top);

  load_tmp_d_21_d_ack : transition
  generic map(1)
  port map(load_tmp_d_21_d_ack_tip, load_tmp_d_21_d_ack_ge, load_tmp_d_21_d_ack_top);

  load_tmp_d_21_d_req : transition
  generic map(1)
  port map(load_tmp_d_21_d_req_tip, load_tmp_d_21_d_req_ge, load_tmp_d_21_d_req_top);

  load_tmp_d_230_d_ack : transition
  generic map(1)
  port map(load_tmp_d_230_d_ack_tip, load_tmp_d_230_d_ack_ge, load_tmp_d_230_d_ack_top);

  load_tmp_d_230_d_req : transition
  generic map(1)
  port map(load_tmp_d_230_d_req_tip, load_tmp_d_230_d_req_ge, load_tmp_d_230_d_req_top);

  load_tmp_d_26_d_ack : transition
  generic map(1)
  port map(load_tmp_d_26_d_ack_tip, load_tmp_d_26_d_ack_ge, load_tmp_d_26_d_ack_top);

  load_tmp_d_26_d_req : transition
  generic map(2)
  port map(load_tmp_d_26_d_req_tip, load_tmp_d_26_d_req_ge, load_tmp_d_26_d_req_top);

  load_tmp_d_31_d_ack : transition
  generic map(1)
  port map(load_tmp_d_31_d_ack_tip, load_tmp_d_31_d_ack_ge, load_tmp_d_31_d_ack_top);

  load_tmp_d_31_d_req : transition
  generic map(2)
  port map(load_tmp_d_31_d_req_tip, load_tmp_d_31_d_req_ge, load_tmp_d_31_d_req_top);

  load_tmp_d_48_d_ack : transition
  generic map(1)
  port map(load_tmp_d_48_d_ack_tip, load_tmp_d_48_d_ack_ge, load_tmp_d_48_d_ack_top);

  load_tmp_d_48_d_req : transition
  generic map(1)
  port map(load_tmp_d_48_d_req_tip, load_tmp_d_48_d_req_ge, load_tmp_d_48_d_req_top);

  load_tmp_d_53_d_ack : transition
  generic map(1)
  port map(load_tmp_d_53_d_ack_tip, load_tmp_d_53_d_ack_ge, load_tmp_d_53_d_ack_top);

  load_tmp_d_53_d_req : transition
  generic map(1)
  port map(load_tmp_d_53_d_req_tip, load_tmp_d_53_d_req_ge, load_tmp_d_53_d_req_top);

  load_tmp_d_66_d_ack : transition
  generic map(1)
  port map(load_tmp_d_66_d_ack_tip, load_tmp_d_66_d_ack_ge, load_tmp_d_66_d_ack_top);

  load_tmp_d_66_d_req : transition
  generic map(1)
  port map(load_tmp_d_66_d_req_tip, load_tmp_d_66_d_req_ge, load_tmp_d_66_d_req_top);

  load_tmp_d_75_d_ack : transition
  generic map(1)
  port map(load_tmp_d_75_d_ack_tip, load_tmp_d_75_d_ack_ge, load_tmp_d_75_d_ack_top);

  load_tmp_d_75_d_req : transition
  generic map(2)
  port map(load_tmp_d_75_d_req_tip, load_tmp_d_75_d_req_ge, load_tmp_d_75_d_req_top);

  load_u_array_d_ack : transition
  generic map(1)
  port map(load_u_array_d_ack_tip, load_u_array_d_ack_ge, load_u_array_d_ack_top);

  load_u_array_d_req : transition
  generic map(1)
  port map(load_u_array_d_req_tip, load_u_array_d_req_ge, load_u_array_d_req_top);

  loopentry_d_12_d_entry : transition
  generic map(1)
  port map(loopentry_d_12_d_entry_tip, loopentry_d_12_d_entry_ge, loopentry_d_12_d_entry_top);

  loopentry_d_12_d_loopexit_to_loopentry_d_12_src : transition
  generic map(1)
  port map(loopentry_d_12_d_loopexit_to_loopentry_d_12_src_tip, loopentry_d_12_d_loopexit_to_loopentry_d_12_src_ge, loopentry_d_12_d_loopexit_to_loopentry_d_12_src_top);

  loopentry_d_12_d_pre : transition
  generic map(2)
  port map(loopentry_d_12_d_pre_tip, loopentry_d_12_d_pre_ge, loopentry_d_12_d_pre_top);

  loopentry_d_12_to_loopexit_d_12_src : transition
  generic map(1)
  port map(loopentry_d_12_to_loopexit_d_12_src_tip, loopentry_d_12_to_loopexit_d_12_src_ge, loopentry_d_12_to_loopexit_d_12_src_top);

  loopentry_d_12_to_no_exit_d_12_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_12_to_no_exit_d_12_d_preheader_src_tip, loopentry_d_12_to_no_exit_d_12_d_preheader_src_ge, loopentry_d_12_to_no_exit_d_12_d_preheader_src_top);

  loopentry_d_14_d_entry : transition
  generic map(1)
  port map(loopentry_d_14_d_entry_tip, loopentry_d_14_d_entry_ge, loopentry_d_14_d_entry_top);

  loopentry_d_14_d_loopexit_to_loopentry_d_14_src : transition
  generic map(1)
  port map(loopentry_d_14_d_loopexit_to_loopentry_d_14_src_tip, loopentry_d_14_d_loopexit_to_loopentry_d_14_src_ge, loopentry_d_14_d_loopexit_to_loopentry_d_14_src_top);

  loopentry_d_14_d_pre : transition
  generic map(2)
  port map(loopentry_d_14_d_pre_tip, loopentry_d_14_d_pre_ge, loopentry_d_14_d_pre_top);

  loopentry_d_14_to_loopexit_d_14_src : transition
  generic map(1)
  port map(loopentry_d_14_to_loopexit_d_14_src_tip, loopentry_d_14_to_loopexit_d_14_src_ge, loopentry_d_14_to_loopexit_d_14_src_top);

  loopentry_d_14_to_no_exit_d_14_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_14_to_no_exit_d_14_d_preheader_src_tip, loopentry_d_14_to_no_exit_d_14_d_preheader_src_ge, loopentry_d_14_to_no_exit_d_14_d_preheader_src_top);

  loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_tip, loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_ge, loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_top);

  loopentry_d_2_to_no_exit_d_2_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_2_to_no_exit_d_2_d_preheader_src_tip, loopentry_d_2_to_no_exit_d_2_d_preheader_src_ge, loopentry_d_2_to_no_exit_d_2_d_preheader_src_top);

  loopentry_d_4_d_entry : transition
  generic map(1)
  port map(loopentry_d_4_d_entry_tip, loopentry_d_4_d_entry_ge, loopentry_d_4_d_entry_top);

  loopentry_d_4_d_loopexit_to_loopentry_d_4_src : transition
  generic map(1)
  port map(loopentry_d_4_d_loopexit_to_loopentry_d_4_src_tip, loopentry_d_4_d_loopexit_to_loopentry_d_4_src_ge, loopentry_d_4_d_loopexit_to_loopentry_d_4_src_top);

  loopentry_d_4_d_outer_d_entry : transition
  generic map(1)
  port map(loopentry_d_4_d_outer_d_entry_tip, loopentry_d_4_d_outer_d_entry_ge, loopentry_d_4_d_outer_d_entry_top);

  loopentry_d_4_d_outer_d_pre : transition
  generic map(3)
  port map(loopentry_d_4_d_outer_d_pre_tip, loopentry_d_4_d_outer_d_pre_ge, loopentry_d_4_d_outer_d_pre_top);

  loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src : transition
  generic map(1)
  port map(loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_tip, loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_ge, loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top);

  loopentry_d_4_d_outer_to_loopentry_d_4_src : transition
  generic map(4)
  port map(loopentry_d_4_d_outer_to_loopentry_d_4_src_tip, loopentry_d_4_d_outer_to_loopentry_d_4_src_ge, loopentry_d_4_d_outer_to_loopentry_d_4_src_top);

  loopentry_d_4_d_pre : transition
  generic map(2)
  port map(loopentry_d_4_d_pre_tip, loopentry_d_4_d_pre_ge, loopentry_d_4_d_pre_top);

  loopentry_d_4_to_no_exit_d_4_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_4_to_no_exit_d_4_d_preheader_src_tip, loopentry_d_4_to_no_exit_d_4_d_preheader_src_ge, loopentry_d_4_to_no_exit_d_4_d_preheader_src_top);

  loopentry_d_4_to_no_exit_d_5_d_preheader_src : transition
  generic map(1)
  port map(loopentry_d_4_to_no_exit_d_5_d_preheader_src_tip, loopentry_d_4_to_no_exit_d_5_d_preheader_src_ge, loopentry_d_4_to_no_exit_d_5_d_preheader_src_top);

  loopentry_d_7_d_outer_d_entry : transition
  generic map(1)
  port map(loopentry_d_7_d_outer_d_entry_tip, loopentry_d_7_d_outer_d_entry_ge, loopentry_d_7_d_outer_d_entry_top);

  loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src : transition
  generic map(1)
  port map(loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_tip, loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_ge, loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_top);

  loopentry_d_7_d_outer_d_pre : transition
  generic map(2)
  port map(loopentry_d_7_d_outer_d_pre_tip, loopentry_d_7_d_outer_d_pre_ge, loopentry_d_7_d_outer_d_pre_top);

  loopentry_d_7_d_outer_to_loopentry_d_7_src : transition
  generic map(4)
  port map(loopentry_d_7_d_outer_to_loopentry_d_7_src_tip, loopentry_d_7_d_outer_to_loopentry_d_7_src_ge, loopentry_d_7_d_outer_to_loopentry_d_7_src_top);

  loopentry_d_7_to_loopexit_d_7_src : transition
  generic map(1)
  port map(loopentry_d_7_to_loopexit_d_7_src_tip, loopentry_d_7_to_loopexit_d_7_src_ge, loopentry_d_7_to_loopexit_d_7_src_top);

  loopentry_d_7_to_no_exit_d_7_src : transition
  generic map(1)
  port map(loopentry_d_7_to_no_exit_d_7_src_tip, loopentry_d_7_to_no_exit_d_7_src_ge, loopentry_d_7_to_no_exit_d_7_src_top);

  loopexit_d_10_to_loopentry_d_12_d_loopexit_src : transition
  generic map(1)
  port map(loopexit_d_10_to_loopentry_d_12_d_loopexit_src_tip, loopexit_d_10_to_loopentry_d_12_d_loopexit_src_ge, loopexit_d_10_to_loopentry_d_12_d_loopexit_src_top);

  loopexit_d_10_to_no_exit_d_10_d_outer_src : transition
  generic map(1)
  port map(loopexit_d_10_to_no_exit_d_10_d_outer_src_tip, loopexit_d_10_to_no_exit_d_10_d_outer_src_ge, loopexit_d_10_to_no_exit_d_10_d_outer_src_top);

  loopexit_d_12_d_entry : transition
  generic map(1)
  port map(loopexit_d_12_d_entry_tip, loopexit_d_12_d_entry_ge, loopexit_d_12_d_entry_top);

  loopexit_d_12_to_loopentry_d_12_src : transition
  generic map(1)
  port map(loopexit_d_12_to_loopentry_d_12_src_tip, loopexit_d_12_to_loopentry_d_12_src_ge, loopexit_d_12_to_loopentry_d_12_src_top);

  loopexit_d_12_to_loopentry_d_14_d_loopexit_src : transition
  generic map(1)
  port map(loopexit_d_12_to_loopentry_d_14_d_loopexit_src_tip, loopexit_d_12_to_loopentry_d_14_d_loopexit_src_ge, loopexit_d_12_to_loopentry_d_14_d_loopexit_src_top);

  loopexit_d_14_d_entry : transition
  generic map(1)
  port map(loopexit_d_14_d_entry_tip, loopexit_d_14_d_entry_ge, loopexit_d_14_d_entry_top);

  loopexit_d_14_to_loopentry_d_14_src : transition
  generic map(1)
  port map(loopexit_d_14_to_loopentry_d_14_src_tip, loopexit_d_14_to_loopentry_d_14_src_ge, loopexit_d_14_to_loopentry_d_14_src_top);

  loopexit_d_14_to_return_src : transition
  generic map(1)
  port map(loopexit_d_14_to_return_src_tip, loopexit_d_14_to_return_src_ge, loopexit_d_14_to_return_src_top);

  loopexit_d_1_to_loopentry_d_2_src : transition
  generic map(1)
  port map(loopexit_d_1_to_loopentry_d_2_src_tip, loopexit_d_1_to_loopentry_d_2_src_ge, loopexit_d_1_to_loopentry_d_2_src_top);

  loopexit_d_1_to_no_exit_d_1_d_outer_src : transition
  generic map(1)
  port map(loopexit_d_1_to_no_exit_d_1_d_outer_src_tip, loopexit_d_1_to_no_exit_d_1_d_outer_src_ge, loopexit_d_1_to_no_exit_d_1_d_outer_src_top);

  loopexit_d_5_d_entry : transition
  generic map(1)
  port map(loopexit_d_5_d_entry_tip, loopexit_d_5_d_entry_ge, loopexit_d_5_d_entry_top);

  loopexit_d_5_to_loopentry_d_4_d_outer_src : transition
  generic map(1)
  port map(loopexit_d_5_to_loopentry_d_4_d_outer_src_tip, loopexit_d_5_to_loopentry_d_4_d_outer_src_ge, loopexit_d_5_to_loopentry_d_4_d_outer_src_top);

  loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src : transition
  generic map(1)
  port map(loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_tip, loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_ge, loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_top);

  loopexit_d_7_to_loopentry_d_7_d_outer_src : transition
  generic map(1)
  port map(loopexit_d_7_to_loopentry_d_7_d_outer_src_tip, loopexit_d_7_to_loopentry_d_7_d_outer_src_ge, loopexit_d_7_to_loopentry_d_7_d_outer_src_top);

  loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src : transition
  generic map(1)
  port map(loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_tip, loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_ge, loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_top);

  maxcoeff_d_2_d_2_mux_1_d_ack : transition
  generic map(1)
  port map(maxcoeff_d_2_d_2_mux_1_d_ack_tip, maxcoeff_d_2_d_2_mux_1_d_ack_ge, maxcoeff_d_2_d_2_mux_1_d_ack_top);

  maxcoeff_d_2_d_2_mux_1_d_req0 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_2_mux_1_d_req0_tip, maxcoeff_d_2_d_2_mux_1_d_req0_ge, maxcoeff_d_2_d_2_mux_1_d_req0_top);

  maxcoeff_d_2_d_2_mux_1_d_req1 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_2_mux_1_d_req1_tip, maxcoeff_d_2_d_2_mux_1_d_req1_ge, maxcoeff_d_2_d_2_mux_1_d_req1_top);

  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack : transition
  generic map(1)
  port map(maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_tip, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_ge, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_top);

  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_tip, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_ge, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_top);

  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_tip, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_ge, maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_top);

  maxcoeff_d_2_d_ph_mux_1_d_ack : transition
  generic map(1)
  port map(maxcoeff_d_2_d_ph_mux_1_d_ack_tip, maxcoeff_d_2_d_ph_mux_1_d_ack_ge, maxcoeff_d_2_d_ph_mux_1_d_ack_top);

  maxcoeff_d_2_d_ph_mux_1_d_req0 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_ph_mux_1_d_req0_tip, maxcoeff_d_2_d_ph_mux_1_d_req0_ge, maxcoeff_d_2_d_ph_mux_1_d_req0_top);

  maxcoeff_d_2_d_ph_mux_1_d_req1 : transition
  generic map(1)
  port map(maxcoeff_d_2_d_ph_mux_1_d_req1_tip, maxcoeff_d_2_d_ph_mux_1_d_req1_ge, maxcoeff_d_2_d_ph_mux_1_d_req1_top);

  maxcoeff_d_2_mux_1_d_ack : transition
  generic map(1)
  port map(maxcoeff_d_2_mux_1_d_ack_tip, maxcoeff_d_2_mux_1_d_ack_ge, maxcoeff_d_2_mux_1_d_ack_top);

  maxcoeff_d_2_mux_1_d_req0 : transition
  generic map(1)
  port map(maxcoeff_d_2_mux_1_d_req0_tip, maxcoeff_d_2_mux_1_d_req0_ge, maxcoeff_d_2_mux_1_d_req0_top);

  maxcoeff_d_2_mux_1_d_req1 : transition
  generic map(1)
  port map(maxcoeff_d_2_mux_1_d_req1_tip, maxcoeff_d_2_mux_1_d_req1_ge, maxcoeff_d_2_mux_1_d_req1_top);

  no_exit_d_10_to_else_d_0_src : transition
  generic map(1)
  port map(no_exit_d_10_to_else_d_0_src_tip, no_exit_d_10_to_else_d_0_src_ge, no_exit_d_10_to_else_d_0_src_top);

  no_exit_d_10_to_then_d_1_src : transition
  generic map(1)
  port map(no_exit_d_10_to_then_d_1_src_tip, no_exit_d_10_to_then_d_1_src_ge, no_exit_d_10_to_then_d_1_src_top);

  no_exit_d_12_d_entry : transition
  generic map(1)
  port map(no_exit_d_12_d_entry_tip, no_exit_d_12_d_entry_ge, no_exit_d_12_d_entry_top);

  no_exit_d_12_to_loopexit_d_12_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_12_to_loopexit_d_12_d_loopexit_src_tip, no_exit_d_12_to_loopexit_d_12_d_loopexit_src_ge, no_exit_d_12_to_loopexit_d_12_d_loopexit_src_top);

  no_exit_d_12_to_no_exit_d_12_src : transition
  generic map(1)
  port map(no_exit_d_12_to_no_exit_d_12_src_tip, no_exit_d_12_to_no_exit_d_12_src_ge, no_exit_d_12_to_no_exit_d_12_src_top);

  no_exit_d_14_d_entry : transition
  generic map(1)
  port map(no_exit_d_14_d_entry_tip, no_exit_d_14_d_entry_ge, no_exit_d_14_d_entry_top);

  no_exit_d_14_to_loopexit_d_14_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_14_to_loopexit_d_14_d_loopexit_src_tip, no_exit_d_14_to_loopexit_d_14_d_loopexit_src_ge, no_exit_d_14_to_loopexit_d_14_d_loopexit_src_top);

  no_exit_d_14_to_no_exit_d_14_src : transition
  generic map(1)
  port map(no_exit_d_14_to_no_exit_d_14_src_tip, no_exit_d_14_to_no_exit_d_14_src_ge, no_exit_d_14_to_no_exit_d_14_src_top);

  no_exit_d_1_d_entry : transition
  generic map(1)
  port map(no_exit_d_1_d_entry_tip, no_exit_d_1_d_entry_ge, no_exit_d_1_d_entry_top);

  no_exit_d_1_to_loopexit_d_1_src : transition
  generic map(1)
  port map(no_exit_d_1_to_loopexit_d_1_src_tip, no_exit_d_1_to_loopexit_d_1_src_ge, no_exit_d_1_to_loopexit_d_1_src_top);

  no_exit_d_1_to_no_exit_d_1_src : transition
  generic map(1)
  port map(no_exit_d_1_to_no_exit_d_1_src_tip, no_exit_d_1_to_no_exit_d_1_src_ge, no_exit_d_1_to_no_exit_d_1_src_top);

  no_exit_d_2_d_entry : transition
  generic map(1)
  port map(no_exit_d_2_d_entry_tip, no_exit_d_2_d_entry_ge, no_exit_d_2_d_entry_top);

  no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_tip, no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_ge, no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_top);

  no_exit_d_2_to_no_exit_d_2_src : transition
  generic map(1)
  port map(no_exit_d_2_to_no_exit_d_2_src_tip, no_exit_d_2_to_no_exit_d_2_src_ge, no_exit_d_2_to_no_exit_d_2_src_top);

  no_exit_d_4_d_entry : transition
  generic map(1)
  port map(no_exit_d_4_d_entry_tip, no_exit_d_4_d_entry_ge, no_exit_d_4_d_entry_top);

  no_exit_d_4_d_pre : transition
  generic map(2)
  port map(no_exit_d_4_d_pre_tip, no_exit_d_4_d_pre_ge, no_exit_d_4_d_pre_top);

  no_exit_d_4_d_preheader_d_entry : transition
  generic map(1)
  port map(no_exit_d_4_d_preheader_d_entry_tip, no_exit_d_4_d_preheader_d_entry_ge, no_exit_d_4_d_preheader_d_entry_top);

  no_exit_d_4_d_preheader_to_no_exit_d_4_src : transition
  generic map(2)
  port map(no_exit_d_4_d_preheader_to_no_exit_d_4_src_tip, no_exit_d_4_d_preheader_to_no_exit_d_4_src_ge, no_exit_d_4_d_preheader_to_no_exit_d_4_src_top);

  no_exit_d_4_to_loopentry_d_4_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_4_to_loopentry_d_4_d_loopexit_src_tip, no_exit_d_4_to_loopentry_d_4_d_loopexit_src_ge, no_exit_d_4_to_loopentry_d_4_d_loopexit_src_top);

  no_exit_d_4_to_then_d_0_src : transition
  generic map(1)
  port map(no_exit_d_4_to_then_d_0_src_tip, no_exit_d_4_to_then_d_0_src_ge, no_exit_d_4_to_then_d_0_src_top);

  no_exit_d_5_d_entry : transition
  generic map(1)
  port map(no_exit_d_5_d_entry_tip, no_exit_d_5_d_entry_ge, no_exit_d_5_d_entry_top);

  no_exit_d_5_to_loopexit_d_5_src : transition
  generic map(1)
  port map(no_exit_d_5_to_loopexit_d_5_src_tip, no_exit_d_5_to_loopexit_d_5_src_ge, no_exit_d_5_to_loopexit_d_5_src_top);

  no_exit_d_5_to_no_exit_d_5_src : transition
  generic map(1)
  port map(no_exit_d_5_to_no_exit_d_5_src_tip, no_exit_d_5_to_no_exit_d_5_src_ge, no_exit_d_5_to_no_exit_d_5_src_top);

  no_exit_d_7_d_entry : transition
  generic map(1)
  port map(no_exit_d_7_d_entry_tip, no_exit_d_7_d_entry_ge, no_exit_d_7_d_entry_top);

  no_exit_d_7_to_loopentry_d_7_d_backedge_src : transition
  generic map(1)
  port map(no_exit_d_7_to_loopentry_d_7_d_backedge_src_tip, no_exit_d_7_to_loopentry_d_7_d_backedge_src_ge, no_exit_d_7_to_loopentry_d_7_d_backedge_src_top);

  no_exit_d_7_to_no_exit_d_8_d_preheader_src : transition
  generic map(1)
  port map(no_exit_d_7_to_no_exit_d_8_d_preheader_src_tip, no_exit_d_7_to_no_exit_d_8_d_preheader_src_ge, no_exit_d_7_to_no_exit_d_8_d_preheader_src_top);

  no_exit_d_8_d_entry : transition
  generic map(1)
  port map(no_exit_d_8_d_entry_tip, no_exit_d_8_d_entry_ge, no_exit_d_8_d_entry_top);

  no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src : transition
  generic map(1)
  port map(no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_tip, no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_ge, no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_top);

  no_exit_d_8_to_no_exit_d_8_src : transition
  generic map(1)
  port map(no_exit_d_8_to_no_exit_d_8_src_tip, no_exit_d_8_to_no_exit_d_8_src_ge, no_exit_d_8_to_no_exit_d_8_src_top);

  oper_exitcond120_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond120_bool_d_ack_tip, oper_exitcond120_bool_d_ack_ge, oper_exitcond120_bool_d_ack_top);

  oper_exitcond120_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond120_bool_d_req_tip, oper_exitcond120_bool_d_req_ge, oper_exitcond120_bool_d_req_top);

  oper_exitcond128_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond128_bool_d_ack_tip, oper_exitcond128_bool_d_ack_ge, oper_exitcond128_bool_d_ack_top);

  oper_exitcond128_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond128_bool_d_req_tip, oper_exitcond128_bool_d_req_ge, oper_exitcond128_bool_d_req_top);

  oper_exitcond131_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond131_bool_d_ack_tip, oper_exitcond131_bool_d_ack_ge, oper_exitcond131_bool_d_ack_top);

  oper_exitcond131_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond131_bool_d_req_tip, oper_exitcond131_bool_d_req_ge, oper_exitcond131_bool_d_req_top);

  oper_exitcond142_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond142_bool_d_ack_tip, oper_exitcond142_bool_d_ack_ge, oper_exitcond142_bool_d_ack_top);

  oper_exitcond142_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond142_bool_d_req_tip, oper_exitcond142_bool_d_req_ge, oper_exitcond142_bool_d_req_top);

  oper_exitcond145_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond145_bool_d_ack_tip, oper_exitcond145_bool_d_ack_ge, oper_exitcond145_bool_d_ack_top);

  oper_exitcond145_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond145_bool_d_req_tip, oper_exitcond145_bool_d_req_ge, oper_exitcond145_bool_d_req_top);

  oper_exitcond150_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond150_bool_d_ack_tip, oper_exitcond150_bool_d_ack_ge, oper_exitcond150_bool_d_ack_top);

  oper_exitcond150_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond150_bool_d_req_tip, oper_exitcond150_bool_d_req_ge, oper_exitcond150_bool_d_req_top);

  oper_exitcond158_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond158_bool_d_ack_tip, oper_exitcond158_bool_d_ack_ge, oper_exitcond158_bool_d_ack_top);

  oper_exitcond158_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond158_bool_d_req_tip, oper_exitcond158_bool_d_req_ge, oper_exitcond158_bool_d_req_top);

  oper_exitcond_bool_d_ack : transition
  generic map(1)
  port map(oper_exitcond_bool_d_ack_tip, oper_exitcond_bool_d_ack_ge, oper_exitcond_bool_d_ack_top);

  oper_exitcond_bool_d_req : transition
  generic map(1)
  port map(oper_exitcond_bool_d_req_tip, oper_exitcond_bool_d_req_ge, oper_exitcond_bool_d_req_top);

  oper_inc_d_11_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_11_int_d_ack_tip, oper_inc_d_11_int_d_ack_ge, oper_inc_d_11_int_d_ack_top);

  oper_inc_d_11_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_11_int_d_req_tip, oper_inc_d_11_int_d_req_ge, oper_inc_d_11_int_d_req_top);

  oper_inc_d_12_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_12_int_d_ack_tip, oper_inc_d_12_int_d_ack_ge, oper_inc_d_12_int_d_ack_top);

  oper_inc_d_12_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_12_int_d_req_tip, oper_inc_d_12_int_d_req_ge, oper_inc_d_12_int_d_req_top);

  oper_inc_d_14_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_14_int_d_ack_tip, oper_inc_d_14_int_d_ack_ge, oper_inc_d_14_int_d_ack_top);

  oper_inc_d_14_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_14_int_d_req_tip, oper_inc_d_14_int_d_req_ge, oper_inc_d_14_int_d_req_top);

  oper_inc_d_15_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_15_int_d_ack_tip, oper_inc_d_15_int_d_ack_ge, oper_inc_d_15_int_d_ack_top);

  oper_inc_d_15_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_15_int_d_req_tip, oper_inc_d_15_int_d_req_ge, oper_inc_d_15_int_d_req_top);

  oper_inc_d_2_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_2_int_d_ack_tip, oper_inc_d_2_int_d_ack_ge, oper_inc_d_2_int_d_ack_top);

  oper_inc_d_2_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_2_int_d_req_tip, oper_inc_d_2_int_d_req_ge, oper_inc_d_2_int_d_req_top);

  oper_inc_d_5_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_5_int_d_ack_tip, oper_inc_d_5_int_d_ack_ge, oper_inc_d_5_int_d_ack_top);

  oper_inc_d_5_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_5_int_d_req_tip, oper_inc_d_5_int_d_req_ge, oper_inc_d_5_int_d_req_top);

  oper_inc_d_960_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_960_int_d_ack_tip, oper_inc_d_960_int_d_ack_ge, oper_inc_d_960_int_d_ack_top);

  oper_inc_d_960_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_960_int_d_req_tip, oper_inc_d_960_int_d_req_ge, oper_inc_d_960_int_d_req_top);

  oper_inc_d_976_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_976_int_d_ack_tip, oper_inc_d_976_int_d_ack_ge, oper_inc_d_976_int_d_ack_top);

  oper_inc_d_976_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_976_int_d_req_tip, oper_inc_d_976_int_d_req_ge, oper_inc_d_976_int_d_req_top);

  oper_inc_d_9_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_9_int_d_ack_tip, oper_inc_d_9_int_d_ack_ge, oper_inc_d_9_int_d_ack_top);

  oper_inc_d_9_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_9_int_d_req_tip, oper_inc_d_9_int_d_req_ge, oper_inc_d_9_int_d_req_top);

  oper_indvar_d_next119_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next119_uint_d_ack_tip, oper_indvar_d_next119_uint_d_ack_ge, oper_indvar_d_next119_uint_d_ack_top);

  oper_indvar_d_next119_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next119_uint_d_req_tip, oper_indvar_d_next119_uint_d_req_ge, oper_indvar_d_next119_uint_d_req_top);

  oper_indvar_d_next122_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next122_uint_d_ack_tip, oper_indvar_d_next122_uint_d_ack_ge, oper_indvar_d_next122_uint_d_ack_top);

  oper_indvar_d_next122_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next122_uint_d_req_tip, oper_indvar_d_next122_uint_d_req_ge, oper_indvar_d_next122_uint_d_req_top);

  oper_indvar_d_next124_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next124_uint_d_ack_tip, oper_indvar_d_next124_uint_d_ack_ge, oper_indvar_d_next124_uint_d_ack_top);

  oper_indvar_d_next124_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next124_uint_d_req_tip, oper_indvar_d_next124_uint_d_req_ge, oper_indvar_d_next124_uint_d_req_top);

  oper_indvar_d_next127_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next127_uint_d_ack_tip, oper_indvar_d_next127_uint_d_ack_ge, oper_indvar_d_next127_uint_d_ack_top);

  oper_indvar_d_next127_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next127_uint_d_req_tip, oper_indvar_d_next127_uint_d_req_ge, oper_indvar_d_next127_uint_d_req_top);

  oper_indvar_d_next130_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next130_uint_d_ack_tip, oper_indvar_d_next130_uint_d_ack_ge, oper_indvar_d_next130_uint_d_ack_top);

  oper_indvar_d_next130_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next130_uint_d_req_tip, oper_indvar_d_next130_uint_d_req_ge, oper_indvar_d_next130_uint_d_req_top);

  oper_indvar_d_next133_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next133_uint_d_ack_tip, oper_indvar_d_next133_uint_d_ack_ge, oper_indvar_d_next133_uint_d_ack_top);

  oper_indvar_d_next133_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next133_uint_d_req_tip, oper_indvar_d_next133_uint_d_req_ge, oper_indvar_d_next133_uint_d_req_top);

  oper_indvar_d_next139_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next139_uint_d_ack_tip, oper_indvar_d_next139_uint_d_ack_ge, oper_indvar_d_next139_uint_d_ack_top);

  oper_indvar_d_next139_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next139_uint_d_req_tip, oper_indvar_d_next139_uint_d_req_ge, oper_indvar_d_next139_uint_d_req_top);

  oper_indvar_d_next144_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next144_uint_d_ack_tip, oper_indvar_d_next144_uint_d_ack_ge, oper_indvar_d_next144_uint_d_ack_top);

  oper_indvar_d_next144_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next144_uint_d_req_tip, oper_indvar_d_next144_uint_d_req_ge, oper_indvar_d_next144_uint_d_req_top);

  oper_indvar_d_next147_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next147_uint_d_ack_tip, oper_indvar_d_next147_uint_d_ack_ge, oper_indvar_d_next147_uint_d_ack_top);

  oper_indvar_d_next147_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next147_uint_d_req_tip, oper_indvar_d_next147_uint_d_req_ge, oper_indvar_d_next147_uint_d_req_top);

  oper_indvar_d_next149_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next149_uint_d_ack_tip, oper_indvar_d_next149_uint_d_ack_ge, oper_indvar_d_next149_uint_d_ack_top);

  oper_indvar_d_next149_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next149_uint_d_req_tip, oper_indvar_d_next149_uint_d_req_ge, oper_indvar_d_next149_uint_d_req_top);

  oper_indvar_d_next152_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next152_uint_d_ack_tip, oper_indvar_d_next152_uint_d_ack_ge, oper_indvar_d_next152_uint_d_ack_top);

  oper_indvar_d_next152_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next152_uint_d_req_tip, oper_indvar_d_next152_uint_d_req_ge, oper_indvar_d_next152_uint_d_req_top);

  oper_indvar_d_next157_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next157_uint_d_ack_tip, oper_indvar_d_next157_uint_d_ack_ge, oper_indvar_d_next157_uint_d_ack_top);

  oper_indvar_d_next157_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next157_uint_d_req_tip, oper_indvar_d_next157_uint_d_req_ge, oper_indvar_d_next157_uint_d_req_top);

  oper_indvar_d_next_uint_d_ack : transition
  generic map(1)
  port map(oper_indvar_d_next_uint_d_ack_tip, oper_indvar_d_next_uint_d_ack_ge, oper_indvar_d_next_uint_d_ack_top);

  oper_indvar_d_next_uint_d_req : transition
  generic map(1)
  port map(oper_indvar_d_next_uint_d_req_tip, oper_indvar_d_next_uint_d_req_ge, oper_indvar_d_next_uint_d_req_top);

  oper_j_d_321_int_d_ack : transition
  generic map(1)
  port map(oper_j_d_321_int_d_ack_tip, oper_j_d_321_int_d_ack_ge, oper_j_d_321_int_d_ack_top);

  oper_j_d_321_int_d_req : transition
  generic map(1)
  port map(oper_j_d_321_int_d_req_tip, oper_j_d_321_int_d_req_ge, oper_j_d_321_int_d_req_top);

  oper_j_d_3_int_d_ack : transition
  generic map(1)
  port map(oper_j_d_3_int_d_ack_tip, oper_j_d_3_int_d_ack_ge, oper_j_d_3_int_d_ack_top);

  oper_j_d_3_int_d_req : transition
  generic map(1)
  port map(oper_j_d_3_int_d_req_tip, oper_j_d_3_int_d_req_ge, oper_j_d_3_int_d_req_top);

  oper_j_d_746_int_d_ack : transition
  generic map(1)
  port map(oper_j_d_746_int_d_ack_tip, oper_j_d_746_int_d_ack_ge, oper_j_d_746_int_d_ack_top);

  oper_j_d_746_int_d_req : transition
  generic map(1)
  port map(oper_j_d_746_int_d_req_tip, oper_j_d_746_int_d_req_ge, oper_j_d_746_int_d_req_top);

  oper_j_d_7_int_d_ack : transition
  generic map(1)
  port map(oper_j_d_7_int_d_ack_tip, oper_j_d_7_int_d_ack_ge, oper_j_d_7_int_d_ack_top);

  oper_j_d_7_int_d_req : transition
  generic map(1)
  port map(oper_j_d_7_int_d_req_tip, oper_j_d_7_int_d_req_ge, oper_j_d_7_int_d_req_top);

  oper_k_d_1_d_in_int_d_ack : transition
  generic map(1)
  port map(oper_k_d_1_d_in_int_d_ack_tip, oper_k_d_1_d_in_int_d_ack_ge, oper_k_d_1_d_in_int_d_ack_top);

  oper_k_d_1_d_in_int_d_req : transition
  generic map(1)
  port map(oper_k_d_1_d_in_int_d_req_tip, oper_k_d_1_d_in_int_d_req_ge, oper_k_d_1_d_in_int_d_req_top);

  oper_k_d_1_int_d_ack : transition
  generic map(1)
  port map(oper_k_d_1_int_d_ack_tip, oper_k_d_1_int_d_ack_ge, oper_k_d_1_int_d_ack_top);

  oper_k_d_1_int_d_req : transition
  generic map(1)
  port map(oper_k_d_1_int_d_req_tip, oper_k_d_1_int_d_req_ge, oper_k_d_1_int_d_req_top);

  oper_k_d_2_d_2_int_d_ack : transition
  generic map(1)
  port map(oper_k_d_2_d_2_int_d_ack_tip, oper_k_d_2_d_2_int_d_ack_ge, oper_k_d_2_d_2_int_d_ack_top);

  oper_k_d_2_d_2_int_d_req : transition
  generic map(1)
  port map(oper_k_d_2_d_2_int_d_req_tip, oper_k_d_2_d_2_int_d_req_ge, oper_k_d_2_d_2_int_d_req_top);

  oper_k_d_4_d_2_int_d_ack : transition
  generic map(1)
  port map(oper_k_d_4_d_2_int_d_ack_tip, oper_k_d_4_d_2_int_d_ack_ge, oper_k_d_4_d_2_int_d_ack_top);

  oper_k_d_4_d_2_int_d_req : transition
  generic map(1)
  port map(oper_k_d_4_d_2_int_d_req_tip, oper_k_d_4_d_2_int_d_req_ge, oper_k_d_4_d_2_int_d_req_top);

  oper_tmp_d_107_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_107_d_id_d_1_uint_d_ack_tip, oper_tmp_d_107_d_id_d_1_uint_d_ack_ge, oper_tmp_d_107_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_107_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_107_d_id_d_1_uint_d_req_tip, oper_tmp_d_107_d_id_d_1_uint_d_req_ge, oper_tmp_d_107_d_id_d_1_uint_d_req_top);

  oper_tmp_d_107_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_107_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_107_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_107_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_107_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_107_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_107_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_107_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_107_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_107_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_107_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_107_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_107_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_107_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_107_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_107_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_11348_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11348_bool_d_ack_tip, oper_tmp_d_11348_bool_d_ack_ge, oper_tmp_d_11348_bool_d_ack_top);

  oper_tmp_d_11348_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11348_bool_d_req_tip, oper_tmp_d_11348_bool_d_req_ge, oper_tmp_d_11348_bool_d_req_top);

  oper_tmp_d_113_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_113_bool_d_ack_tip, oper_tmp_d_113_bool_d_ack_ge, oper_tmp_d_113_bool_d_ack_top);

  oper_tmp_d_113_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_113_bool_d_req_tip, oper_tmp_d_113_bool_d_req_ge, oper_tmp_d_113_bool_d_req_top);

  oper_tmp_d_118_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_118_d_id_d_1_uint_d_ack_tip, oper_tmp_d_118_d_id_d_1_uint_d_ack_ge, oper_tmp_d_118_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_118_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_118_d_id_d_1_uint_d_req_tip, oper_tmp_d_118_d_id_d_1_uint_d_req_ge, oper_tmp_d_118_d_id_d_1_uint_d_req_top);

  oper_tmp_d_118_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_118_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_118_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_118_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_118_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_118_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_118_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_118_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_118_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_118_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_118_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_118_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_118_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_118_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_118_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_118_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_11_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11_d_id_d_1_uint_d_ack_tip, oper_tmp_d_11_d_id_d_1_uint_d_ack_ge, oper_tmp_d_11_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_11_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11_d_id_d_1_uint_d_req_tip, oper_tmp_d_11_d_id_d_1_uint_d_req_ge, oper_tmp_d_11_d_id_d_1_uint_d_req_top);

  oper_tmp_d_11_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_11_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_11_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_11_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_11_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_11_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_11_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_11_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_11_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_11_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_11_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_11_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_125_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_125_uint_d_ack_tip, oper_tmp_d_125_uint_d_ack_ge, oper_tmp_d_125_uint_d_ack_top);

  oper_tmp_d_125_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_125_uint_d_req_tip, oper_tmp_d_125_uint_d_req_ge, oper_tmp_d_125_uint_d_req_top);

  oper_tmp_d_132_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_132_d_id_d_1_uint_d_ack_tip, oper_tmp_d_132_d_id_d_1_uint_d_ack_ge, oper_tmp_d_132_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_132_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_132_d_id_d_1_uint_d_req_tip, oper_tmp_d_132_d_id_d_1_uint_d_req_ge, oper_tmp_d_132_d_id_d_1_uint_d_req_top);

  oper_tmp_d_132_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_132_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_132_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_132_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_132_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_132_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_132_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_132_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_132_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_132_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_132_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_132_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_132_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_132_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_132_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_132_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_134_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_134_float_d_ack_tip, oper_tmp_d_134_float_d_ack_ge, oper_tmp_d_134_float_d_ack_top);

  oper_tmp_d_134_float_d_req : transition
  generic map(2)
  port map(oper_tmp_d_134_float_d_req_tip, oper_tmp_d_134_float_d_req_ge, oper_tmp_d_134_float_d_req_top);

  oper_tmp_d_135_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_135_float_d_ack_tip, oper_tmp_d_135_float_d_ack_ge, oper_tmp_d_135_float_d_ack_top);

  oper_tmp_d_135_float_d_req : transition
  generic map(2)
  port map(oper_tmp_d_135_float_d_req_tip, oper_tmp_d_135_float_d_req_ge, oper_tmp_d_135_float_d_req_top);

  oper_tmp_d_136_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_136_uint_d_ack_tip, oper_tmp_d_136_uint_d_ack_ge, oper_tmp_d_136_uint_d_ack_top);

  oper_tmp_d_136_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_136_uint_d_req_tip, oper_tmp_d_136_uint_d_req_ge, oper_tmp_d_136_uint_d_req_top);

  oper_tmp_d_137_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_137_uint_d_ack_tip, oper_tmp_d_137_uint_d_ack_ge, oper_tmp_d_137_uint_d_ack_top);

  oper_tmp_d_137_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_137_uint_d_req_tip, oper_tmp_d_137_uint_d_req_ge, oper_tmp_d_137_uint_d_req_top);

  oper_tmp_d_14574_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_14574_bool_d_ack_tip, oper_tmp_d_14574_bool_d_ack_ge, oper_tmp_d_14574_bool_d_ack_top);

  oper_tmp_d_14574_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_14574_bool_d_req_tip, oper_tmp_d_14574_bool_d_req_ge, oper_tmp_d_14574_bool_d_req_top);

  oper_tmp_d_14578_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_14578_bool_d_ack_tip, oper_tmp_d_14578_bool_d_ack_ge, oper_tmp_d_14578_bool_d_ack_top);

  oper_tmp_d_14578_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_14578_bool_d_req_tip, oper_tmp_d_14578_bool_d_req_ge, oper_tmp_d_14578_bool_d_req_top);

  oper_tmp_d_14580_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_14580_bool_d_ack_tip, oper_tmp_d_14580_bool_d_ack_ge, oper_tmp_d_14580_bool_d_ack_top);

  oper_tmp_d_14580_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_14580_bool_d_req_tip, oper_tmp_d_14580_bool_d_req_ge, oper_tmp_d_14580_bool_d_req_top);

  oper_tmp_d_149_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_149_bool_d_ack_tip, oper_tmp_d_149_bool_d_ack_ge, oper_tmp_d_149_bool_d_ack_top);

  oper_tmp_d_149_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_149_bool_d_req_tip, oper_tmp_d_149_bool_d_req_ge, oper_tmp_d_149_bool_d_req_top);

  oper_tmp_d_154_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_154_d_id_d_1_uint_d_ack_tip, oper_tmp_d_154_d_id_d_1_uint_d_ack_ge, oper_tmp_d_154_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_154_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_154_d_id_d_1_uint_d_req_tip, oper_tmp_d_154_d_id_d_1_uint_d_req_ge, oper_tmp_d_154_d_id_d_1_uint_d_req_top);

  oper_tmp_d_154_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_154_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_154_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_154_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_154_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_154_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_154_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_154_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_154_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_154_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_154_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_154_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_154_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_154_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_154_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_154_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_155_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_155_uint_d_ack_tip, oper_tmp_d_155_uint_d_ack_ge, oper_tmp_d_155_uint_d_ack_top);

  oper_tmp_d_155_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_155_uint_d_req_tip, oper_tmp_d_155_uint_d_req_ge, oper_tmp_d_155_uint_d_req_top);

  oper_tmp_d_158_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_158_d_id_d_1_uint_d_ack_tip, oper_tmp_d_158_d_id_d_1_uint_d_ack_ge, oper_tmp_d_158_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_158_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_158_d_id_d_1_uint_d_req_tip, oper_tmp_d_158_d_id_d_1_uint_d_req_ge, oper_tmp_d_158_d_id_d_1_uint_d_req_top);

  oper_tmp_d_158_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_158_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_158_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_158_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_158_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_158_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_158_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_158_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_158_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_158_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_158_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_158_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_158_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_158_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_158_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_158_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_1614_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_1614_bool_d_ack_tip, oper_tmp_d_1614_bool_d_ack_ge, oper_tmp_d_1614_bool_d_ack_top);

  oper_tmp_d_1614_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_1614_bool_d_req_tip, oper_tmp_d_1614_bool_d_req_ge, oper_tmp_d_1614_bool_d_req_top);

  oper_tmp_d_163_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_163_d_id_d_1_uint_d_ack_tip, oper_tmp_d_163_d_id_d_1_uint_d_ack_ge, oper_tmp_d_163_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_163_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_163_d_id_d_1_uint_d_req_tip, oper_tmp_d_163_d_id_d_1_uint_d_req_ge, oper_tmp_d_163_d_id_d_1_uint_d_req_top);

  oper_tmp_d_163_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_163_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_163_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_163_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_163_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_163_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_163_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_163_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_163_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_163_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_163_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_163_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_163_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_163_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_163_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_163_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_166_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_166_bool_d_ack_tip, oper_tmp_d_166_bool_d_ack_ge, oper_tmp_d_166_bool_d_ack_top);

  oper_tmp_d_166_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_166_bool_d_req_tip, oper_tmp_d_166_bool_d_req_ge, oper_tmp_d_166_bool_d_req_top);

  oper_tmp_d_16_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_16_bool_d_ack_tip, oper_tmp_d_16_bool_d_ack_ge, oper_tmp_d_16_bool_d_ack_top);

  oper_tmp_d_16_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_16_bool_d_req_tip, oper_tmp_d_16_bool_d_req_ge, oper_tmp_d_16_bool_d_req_top);

  oper_tmp_d_171_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_171_d_id_d_1_uint_d_ack_tip, oper_tmp_d_171_d_id_d_1_uint_d_ack_ge, oper_tmp_d_171_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_171_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_171_d_id_d_1_uint_d_req_tip, oper_tmp_d_171_d_id_d_1_uint_d_req_ge, oper_tmp_d_171_d_id_d_1_uint_d_req_top);

  oper_tmp_d_171_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_171_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_171_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_171_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_171_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_171_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_171_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_171_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_171_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_171_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_171_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_171_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_171_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_171_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_171_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_171_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_175_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_175_d_id_d_1_uint_d_ack_tip, oper_tmp_d_175_d_id_d_1_uint_d_ack_ge, oper_tmp_d_175_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_175_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_175_d_id_d_1_uint_d_req_tip, oper_tmp_d_175_d_id_d_1_uint_d_req_ge, oper_tmp_d_175_d_id_d_1_uint_d_req_top);

  oper_tmp_d_175_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_175_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_175_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_175_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_175_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_175_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_175_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_175_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_175_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_175_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_175_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_175_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_175_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_175_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_175_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_175_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_179_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_179_d_id_d_1_uint_d_ack_tip, oper_tmp_d_179_d_id_d_1_uint_d_ack_ge, oper_tmp_d_179_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_179_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_179_d_id_d_1_uint_d_req_tip, oper_tmp_d_179_d_id_d_1_uint_d_req_ge, oper_tmp_d_179_d_id_d_1_uint_d_req_top);

  oper_tmp_d_179_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_179_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_179_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_179_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_179_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_179_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_179_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_179_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_179_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_179_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_179_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_179_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_179_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_179_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_179_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_179_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_188_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_188_d_id_d_1_uint_d_ack_tip, oper_tmp_d_188_d_id_d_1_uint_d_ack_ge, oper_tmp_d_188_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_188_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_188_d_id_d_1_uint_d_req_tip, oper_tmp_d_188_d_id_d_1_uint_d_req_ge, oper_tmp_d_188_d_id_d_1_uint_d_req_top);

  oper_tmp_d_188_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_188_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_188_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_188_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_188_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_188_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_188_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_188_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_188_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_188_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_188_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_188_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_188_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_188_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_188_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_188_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_192_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_192_d_id_d_1_uint_d_ack_tip, oper_tmp_d_192_d_id_d_1_uint_d_ack_ge, oper_tmp_d_192_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_192_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_192_d_id_d_1_uint_d_req_tip, oper_tmp_d_192_d_id_d_1_uint_d_req_ge, oper_tmp_d_192_d_id_d_1_uint_d_req_top);

  oper_tmp_d_192_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_192_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_192_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_192_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_192_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_192_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_192_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_192_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_192_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_192_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_192_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_192_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_192_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_192_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_192_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_192_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_20299_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_20299_bool_d_ack_tip, oper_tmp_d_20299_bool_d_ack_ge, oper_tmp_d_20299_bool_d_ack_top);

  oper_tmp_d_20299_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_20299_bool_d_req_tip, oper_tmp_d_20299_bool_d_req_ge, oper_tmp_d_20299_bool_d_req_top);

  oper_tmp_d_202_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_202_bool_d_ack_tip, oper_tmp_d_202_bool_d_ack_ge, oper_tmp_d_202_bool_d_ack_top);

  oper_tmp_d_202_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_202_bool_d_req_tip, oper_tmp_d_202_bool_d_req_ge, oper_tmp_d_202_bool_d_req_top);

  oper_tmp_d_206_d_lvl_d_0_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_206_d_lvl_d_0_uint_d_ack_tip, oper_tmp_d_206_d_lvl_d_0_uint_d_ack_ge, oper_tmp_d_206_d_lvl_d_0_uint_d_ack_top);

  oper_tmp_d_206_d_lvl_d_0_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_206_d_lvl_d_0_uint_d_req_tip, oper_tmp_d_206_d_lvl_d_0_uint_d_req_ge, oper_tmp_d_206_d_lvl_d_0_uint_d_req_top);

  oper_tmp_d_20_d_lvl_d_0_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_20_d_lvl_d_0_uint_d_ack_tip, oper_tmp_d_20_d_lvl_d_0_uint_d_ack_ge, oper_tmp_d_20_d_lvl_d_0_uint_d_ack_top);

  oper_tmp_d_20_d_lvl_d_0_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_20_d_lvl_d_0_uint_d_req_tip, oper_tmp_d_20_d_lvl_d_0_uint_d_req_ge, oper_tmp_d_20_d_lvl_d_0_uint_d_req_top);

  oper_tmp_d_210_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_210_d_id_d_1_uint_d_ack_tip, oper_tmp_d_210_d_id_d_1_uint_d_ack_ge, oper_tmp_d_210_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_210_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_210_d_id_d_1_uint_d_req_tip, oper_tmp_d_210_d_id_d_1_uint_d_req_ge, oper_tmp_d_210_d_id_d_1_uint_d_req_top);

  oper_tmp_d_210_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_210_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_210_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_210_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_210_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_210_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_210_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_210_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_210_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_210_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_210_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_210_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_210_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_210_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_210_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_210_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_221111_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_221111_bool_d_ack_tip, oper_tmp_d_221111_bool_d_ack_ge, oper_tmp_d_221111_bool_d_ack_top);

  oper_tmp_d_221111_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_221111_bool_d_req_tip, oper_tmp_d_221111_bool_d_req_ge, oper_tmp_d_221111_bool_d_req_top);

  oper_tmp_d_221_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_221_bool_d_ack_tip, oper_tmp_d_221_bool_d_ack_ge, oper_tmp_d_221_bool_d_ack_top);

  oper_tmp_d_221_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_221_bool_d_req_tip, oper_tmp_d_221_bool_d_req_ge, oper_tmp_d_221_bool_d_req_top);

  oper_tmp_d_225_d_lvl_d_0_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_225_d_lvl_d_0_uint_d_ack_tip, oper_tmp_d_225_d_lvl_d_0_uint_d_ack_ge, oper_tmp_d_225_d_lvl_d_0_uint_d_ack_top);

  oper_tmp_d_225_d_lvl_d_0_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_225_d_lvl_d_0_uint_d_req_tip, oper_tmp_d_225_d_lvl_d_0_uint_d_req_ge, oper_tmp_d_225_d_lvl_d_0_uint_d_req_top);

  oper_tmp_d_229_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_229_d_id_d_1_uint_d_ack_tip, oper_tmp_d_229_d_id_d_1_uint_d_ack_ge, oper_tmp_d_229_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_229_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_229_d_id_d_1_uint_d_req_tip, oper_tmp_d_229_d_id_d_1_uint_d_req_ge, oper_tmp_d_229_d_id_d_1_uint_d_req_top);

  oper_tmp_d_229_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_229_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_229_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_229_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_229_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_229_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_229_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_229_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_229_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_229_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_229_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_229_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_229_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_229_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_229_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_229_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_25_d_lvl_d_0_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_25_d_lvl_d_0_uint_d_ack_tip, oper_tmp_d_25_d_lvl_d_0_uint_d_ack_ge, oper_tmp_d_25_d_lvl_d_0_uint_d_ack_top);

  oper_tmp_d_25_d_lvl_d_0_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_25_d_lvl_d_0_uint_d_req_tip, oper_tmp_d_25_d_lvl_d_0_uint_d_req_ge, oper_tmp_d_25_d_lvl_d_0_uint_d_req_top);

  oper_tmp_d_27_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_27_d_id_d_1_uint_d_ack_tip, oper_tmp_d_27_d_id_d_1_uint_d_ack_ge, oper_tmp_d_27_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_27_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_27_d_id_d_1_uint_d_req_tip, oper_tmp_d_27_d_id_d_1_uint_d_req_ge, oper_tmp_d_27_d_id_d_1_uint_d_req_top);

  oper_tmp_d_27_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_27_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_27_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_27_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_27_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_27_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_27_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_27_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_27_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_27_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_27_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_27_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_27_d_lvl_d_2_uint_d_req : transition
  generic map(2)
  port map(oper_tmp_d_27_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_27_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_27_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_30_d_lvl_d_0_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_30_d_lvl_d_0_uint_d_ack_tip, oper_tmp_d_30_d_lvl_d_0_uint_d_ack_ge, oper_tmp_d_30_d_lvl_d_0_uint_d_ack_top);

  oper_tmp_d_30_d_lvl_d_0_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_30_d_lvl_d_0_uint_d_req_tip, oper_tmp_d_30_d_lvl_d_0_uint_d_req_ge, oper_tmp_d_30_d_lvl_d_0_uint_d_req_top);

  oper_tmp_d_4223_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_4223_bool_d_ack_tip, oper_tmp_d_4223_bool_d_ack_ge, oper_tmp_d_4223_bool_d_ack_top);

  oper_tmp_d_4223_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_4223_bool_d_req_tip, oper_tmp_d_4223_bool_d_req_ge, oper_tmp_d_4223_bool_d_req_top);

  oper_tmp_d_42_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_42_bool_d_ack_tip, oper_tmp_d_42_bool_d_ack_ge, oper_tmp_d_42_bool_d_ack_top);

  oper_tmp_d_42_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_42_bool_d_req_tip, oper_tmp_d_42_bool_d_req_ge, oper_tmp_d_42_bool_d_req_top);

  oper_tmp_d_47_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_47_d_id_d_1_uint_d_ack_tip, oper_tmp_d_47_d_id_d_1_uint_d_ack_ge, oper_tmp_d_47_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_47_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_47_d_id_d_1_uint_d_req_tip, oper_tmp_d_47_d_id_d_1_uint_d_req_ge, oper_tmp_d_47_d_id_d_1_uint_d_req_top);

  oper_tmp_d_47_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_47_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_47_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_47_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_47_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_47_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_47_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_47_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_47_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_47_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_47_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_47_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_47_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_47_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_47_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_47_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_52_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_52_d_id_d_1_uint_d_ack_tip, oper_tmp_d_52_d_id_d_1_uint_d_ack_ge, oper_tmp_d_52_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_52_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_52_d_id_d_1_uint_d_req_tip, oper_tmp_d_52_d_id_d_1_uint_d_req_ge, oper_tmp_d_52_d_id_d_1_uint_d_req_top);

  oper_tmp_d_52_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_52_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_52_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_52_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_52_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_52_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_52_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_52_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_52_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_52_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_52_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_52_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_52_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_52_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_52_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_52_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_54_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_54_bool_d_ack_tip, oper_tmp_d_54_bool_d_ack_ge, oper_tmp_d_54_bool_d_ack_top);

  oper_tmp_d_54_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_54_bool_d_req_tip, oper_tmp_d_54_bool_d_req_ge, oper_tmp_d_54_bool_d_req_top);

  oper_tmp_d_65_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_65_d_id_d_1_uint_d_ack_tip, oper_tmp_d_65_d_id_d_1_uint_d_ack_ge, oper_tmp_d_65_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_65_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_65_d_id_d_1_uint_d_req_tip, oper_tmp_d_65_d_id_d_1_uint_d_req_ge, oper_tmp_d_65_d_id_d_1_uint_d_req_top);

  oper_tmp_d_65_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_65_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_65_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_65_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_65_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_65_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_65_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_65_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_65_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_65_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_65_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_65_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_65_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_65_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_65_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_65_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_74_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_74_d_id_d_1_uint_d_ack_tip, oper_tmp_d_74_d_id_d_1_uint_d_ack_ge, oper_tmp_d_74_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_74_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_74_d_id_d_1_uint_d_req_tip, oper_tmp_d_74_d_id_d_1_uint_d_req_ge, oper_tmp_d_74_d_id_d_1_uint_d_req_top);

  oper_tmp_d_74_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_74_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_74_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_74_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_74_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_74_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_74_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_74_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_74_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_74_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_74_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_74_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_74_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_74_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_74_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_74_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_92_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_92_bool_d_ack_tip, oper_tmp_d_92_bool_d_ack_ge, oper_tmp_d_92_bool_d_ack_top);

  oper_tmp_d_92_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_92_bool_d_req_tip, oper_tmp_d_92_bool_d_req_ge, oper_tmp_d_92_bool_d_req_top);

  oper_tmp_d_97_d_id_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_97_d_id_d_1_uint_d_ack_tip, oper_tmp_d_97_d_id_d_1_uint_d_ack_ge, oper_tmp_d_97_d_id_d_1_uint_d_ack_top);

  oper_tmp_d_97_d_id_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_97_d_id_d_1_uint_d_req_tip, oper_tmp_d_97_d_id_d_1_uint_d_req_ge, oper_tmp_d_97_d_id_d_1_uint_d_req_top);

  oper_tmp_d_97_d_lvl_d_1_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_97_d_lvl_d_1_uint_d_ack_tip, oper_tmp_d_97_d_lvl_d_1_uint_d_ack_ge, oper_tmp_d_97_d_lvl_d_1_uint_d_ack_top);

  oper_tmp_d_97_d_lvl_d_1_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_97_d_lvl_d_1_uint_d_req_tip, oper_tmp_d_97_d_lvl_d_1_uint_d_req_ge, oper_tmp_d_97_d_lvl_d_1_uint_d_req_top);

  oper_tmp_d_97_d_lvl_d_2_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_97_d_lvl_d_2_uint_d_ack_tip, oper_tmp_d_97_d_lvl_d_2_uint_d_ack_ge, oper_tmp_d_97_d_lvl_d_2_uint_d_ack_top);

  oper_tmp_d_97_d_lvl_d_2_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_97_d_lvl_d_2_uint_d_req_tip, oper_tmp_d_97_d_lvl_d_2_uint_d_req_ge, oper_tmp_d_97_d_lvl_d_2_uint_d_req_top);

  oper_tmp_d_uint_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_uint_d_ack_tip, oper_tmp_d_uint_d_ack_ge, oper_tmp_d_uint_d_ack_top);

  oper_tmp_d_uint_d_req : transition
  generic map(1)
  port map(oper_tmp_d_uint_d_req_tip, oper_tmp_d_uint_d_req_ge, oper_tmp_d_uint_d_req_top);

  start_call_divide_0_actual_0_wr_d_ack : transition
  generic map(1)
  port map(start_call_divide_0_actual_0_wr_d_ack_tip, start_call_divide_0_actual_0_wr_d_ack_ge, start_call_divide_0_actual_0_wr_d_ack_top);

  start_call_divide_0_actual_0_wr_d_req : transition
  generic map(2)
  port map(start_call_divide_0_actual_0_wr_d_req_tip, start_call_divide_0_actual_0_wr_d_req_ge, start_call_divide_0_actual_0_wr_d_req_top);

  start_call_divide_0_actual_1_wr_d_ack : transition
  generic map(1)
  port map(start_call_divide_0_actual_1_wr_d_ack_tip, start_call_divide_0_actual_1_wr_d_ack_ge, start_call_divide_0_actual_1_wr_d_ack_top);

  start_call_divide_0_actual_1_wr_d_req : transition
  generic map(2)
  port map(start_call_divide_0_actual_1_wr_d_req_tip, start_call_divide_0_actual_1_wr_d_req_ge, start_call_divide_0_actual_1_wr_d_req_top);

  start_call_divide_0_d_ack : transition
  generic map(1)
  port map(start_call_divide_0_d_ack_tip, start_call_divide_0_d_ack_ge, start_call_divide_0_d_ack_top);

  start_call_divide_0_d_req : transition
  generic map(1)
  port map(start_call_divide_0_d_req_tip, start_call_divide_0_d_req_ge, start_call_divide_0_d_req_top);

  store_0_d_ack : transition
  generic map(1)
  port map(store_0_d_ack_tip, store_0_d_ack_ge, store_0_d_ack_top);

  store_0_d_req : transition
  generic map(1)
  port map(store_0_d_req_tip, store_0_d_req_ge, store_0_d_req_top);

  store_10_d_ack : transition
  generic map(1)
  port map(store_10_d_ack_tip, store_10_d_ack_ge, store_10_d_ack_top);

  store_10_d_req : transition
  generic map(1)
  port map(store_10_d_req_tip, store_10_d_req_ge, store_10_d_req_top);

  store_11_d_ack : transition
  generic map(1)
  port map(store_11_d_ack_tip, store_11_d_ack_ge, store_11_d_ack_top);

  store_11_d_req : transition
  generic map(3)
  port map(store_11_d_req_tip, store_11_d_req_ge, store_11_d_req_top);

  store_12_d_ack : transition
  generic map(1)
  port map(store_12_d_ack_tip, store_12_d_ack_ge, store_12_d_ack_top);

  store_12_d_req : transition
  generic map(3)
  port map(store_12_d_req_tip, store_12_d_req_ge, store_12_d_req_top);

  store_13_d_ack : transition
  generic map(1)
  port map(store_13_d_ack_tip, store_13_d_ack_ge, store_13_d_ack_top);

  store_13_d_req : transition
  generic map(3)
  port map(store_13_d_req_tip, store_13_d_req_ge, store_13_d_req_top);

  store_1_d_ack : transition
  generic map(1)
  port map(store_1_d_ack_tip, store_1_d_ack_ge, store_1_d_ack_top);

  store_1_d_req : transition
  generic map(3)
  port map(store_1_d_req_tip, store_1_d_req_ge, store_1_d_req_top);

  store_2_d_ack : transition
  generic map(1)
  port map(store_2_d_ack_tip, store_2_d_ack_ge, store_2_d_ack_top);

  store_2_d_req : transition
  generic map(3)
  port map(store_2_d_req_tip, store_2_d_req_ge, store_2_d_req_top);

  store_3_d_ack : transition
  generic map(1)
  port map(store_3_d_ack_tip, store_3_d_ack_ge, store_3_d_ack_top);

  store_3_d_req : transition
  generic map(3)
  port map(store_3_d_req_tip, store_3_d_req_ge, store_3_d_req_top);

  store_4_d_ack : transition
  generic map(1)
  port map(store_4_d_ack_tip, store_4_d_ack_ge, store_4_d_ack_top);

  store_4_d_req : transition
  generic map(3)
  port map(store_4_d_req_tip, store_4_d_req_ge, store_4_d_req_top);

  store_5_d_ack : transition
  generic map(1)
  port map(store_5_d_ack_tip, store_5_d_ack_ge, store_5_d_ack_top);

  store_5_d_req : transition
  generic map(3)
  port map(store_5_d_req_tip, store_5_d_req_ge, store_5_d_req_top);

  store_6_d_ack : transition
  generic map(1)
  port map(store_6_d_ack_tip, store_6_d_ack_ge, store_6_d_ack_top);

  store_6_d_req : transition
  generic map(3)
  port map(store_6_d_req_tip, store_6_d_req_ge, store_6_d_req_top);

  store_7_d_ack : transition
  generic map(1)
  port map(store_7_d_ack_tip, store_7_d_ack_ge, store_7_d_ack_top);

  store_7_d_req : transition
  generic map(2)
  port map(store_7_d_req_tip, store_7_d_req_ge, store_7_d_req_top);

  store_8_d_ack : transition
  generic map(1)
  port map(store_8_d_ack_tip, store_8_d_ack_ge, store_8_d_ack_top);

  store_8_d_req : transition
  generic map(1)
  port map(store_8_d_req_tip, store_8_d_req_ge, store_8_d_req_top);

  store_9_d_ack : transition
  generic map(1)
  port map(store_9_d_ack_tip, store_9_d_ack_ge, store_9_d_ack_top);

  store_9_d_req : transition
  generic map(3)
  port map(store_9_d_req_tip, store_9_d_req_ge, store_9_d_req_top);

  tc_i_d_1_d_0_d_ack : transition
  generic map(1)
  port map(tc_i_d_1_d_0_d_ack_tip, tc_i_d_1_d_0_d_ack_ge, tc_i_d_1_d_0_d_ack_top);

  tc_i_d_1_d_0_d_req : transition
  generic map(1)
  port map(tc_i_d_1_d_0_d_req_tip, tc_i_d_1_d_0_d_req_ge, tc_i_d_1_d_0_d_req_top);

  tc_i_d_2_d_0_d_ph_d_ack : transition
  generic map(1)
  port map(tc_i_d_2_d_0_d_ph_d_ack_tip, tc_i_d_2_d_0_d_ph_d_ack_ge, tc_i_d_2_d_0_d_ph_d_ack_top);

  tc_i_d_2_d_0_d_ph_d_req : transition
  generic map(1)
  port map(tc_i_d_2_d_0_d_ph_d_req_tip, tc_i_d_2_d_0_d_ph_d_req_ge, tc_i_d_2_d_0_d_ph_d_req_top);

  tc_i_d_3_d_0_d_ph_d_ack : transition
  generic map(1)
  port map(tc_i_d_3_d_0_d_ph_d_ack_tip, tc_i_d_3_d_0_d_ph_d_ack_ge, tc_i_d_3_d_0_d_ph_d_ack_top);

  tc_i_d_3_d_0_d_ph_d_req : transition
  generic map(1)
  port map(tc_i_d_3_d_0_d_ph_d_req_tip, tc_i_d_3_d_0_d_ph_d_req_ge, tc_i_d_3_d_0_d_ph_d_req_top);

  tc_i_d_4_d_0_d_ack : transition
  generic map(1)
  port map(tc_i_d_4_d_0_d_ack_tip, tc_i_d_4_d_0_d_ack_ge, tc_i_d_4_d_0_d_ack_top);

  tc_i_d_4_d_0_d_req : transition
  generic map(1)
  port map(tc_i_d_4_d_0_d_req_tip, tc_i_d_4_d_0_d_req_ge, tc_i_d_4_d_0_d_req_top);

  tc_i_d_5_d_0_d_ack : transition
  generic map(1)
  port map(tc_i_d_5_d_0_d_ack_tip, tc_i_d_5_d_0_d_ack_ge, tc_i_d_5_d_0_d_ack_top);

  tc_i_d_5_d_0_d_req : transition
  generic map(1)
  port map(tc_i_d_5_d_0_d_req_tip, tc_i_d_5_d_0_d_req_ge, tc_i_d_5_d_0_d_req_top);

  tc_indvar138_d_ack : transition
  generic map(1)
  port map(tc_indvar138_d_ack_tip, tc_indvar138_d_ack_ge, tc_indvar138_d_ack_top);

  tc_indvar138_d_req : transition
  generic map(1)
  port map(tc_indvar138_d_req_tip, tc_indvar138_d_req_ge, tc_indvar138_d_req_top);

  tc_indvar151_d_ack : transition
  generic map(1)
  port map(tc_indvar151_d_ack_tip, tc_indvar151_d_ack_ge, tc_indvar151_d_ack_top);

  tc_indvar151_d_req : transition
  generic map(1)
  port map(tc_indvar151_d_req_tip, tc_indvar151_d_req_ge, tc_indvar151_d_req_top);

  tc_j_d_11_d_2_d_ack : transition
  generic map(1)
  port map(tc_j_d_11_d_2_d_ack_tip, tc_j_d_11_d_2_d_ack_ge, tc_j_d_11_d_2_d_ack_top);

  tc_j_d_11_d_2_d_req : transition
  generic map(1)
  port map(tc_j_d_11_d_2_d_req_tip, tc_j_d_11_d_2_d_req_ge, tc_j_d_11_d_2_d_req_top);

  tc_j_d_13_d_2_d_ack : transition
  generic map(1)
  port map(tc_j_d_13_d_2_d_ack_tip, tc_j_d_13_d_2_d_ack_ge, tc_j_d_13_d_2_d_ack_top);

  tc_j_d_13_d_2_d_req : transition
  generic map(1)
  port map(tc_j_d_13_d_2_d_req_tip, tc_j_d_13_d_2_d_req_ge, tc_j_d_13_d_2_d_req_top);

  tc_j_d_3_d_2_d_ack : transition
  generic map(1)
  port map(tc_j_d_3_d_2_d_ack_tip, tc_j_d_3_d_2_d_ack_ge, tc_j_d_3_d_2_d_ack_top);

  tc_j_d_3_d_2_d_req : transition
  generic map(1)
  port map(tc_j_d_3_d_2_d_req_tip, tc_j_d_3_d_2_d_req_ge, tc_j_d_3_d_2_d_req_top);

  tc_j_d_3_d_in_d_ack : transition
  generic map(1)
  port map(tc_j_d_3_d_in_d_ack_tip, tc_j_d_3_d_in_d_ack_ge, tc_j_d_3_d_in_d_ack_top);

  tc_j_d_3_d_in_d_req : transition
  generic map(1)
  port map(tc_j_d_3_d_in_d_req_tip, tc_j_d_3_d_in_d_req_ge, tc_j_d_3_d_in_d_req_top);

  tc_j_d_7_d_1_d_ack : transition
  generic map(1)
  port map(tc_j_d_7_d_1_d_ack_tip, tc_j_d_7_d_1_d_ack_ge, tc_j_d_7_d_1_d_ack_top);

  tc_j_d_7_d_1_d_req : transition
  generic map(1)
  port map(tc_j_d_7_d_1_d_req_tip, tc_j_d_7_d_1_d_req_ge, tc_j_d_7_d_1_d_req_top);

  tc_p_d_0_d_0_d_ph_d_ack : transition
  generic map(1)
  port map(tc_p_d_0_d_0_d_ph_d_ack_tip, tc_p_d_0_d_0_d_ph_d_ack_ge, tc_p_d_0_d_0_d_ph_d_ack_top);

  tc_p_d_0_d_0_d_ph_d_req : transition
  generic map(1)
  port map(tc_p_d_0_d_0_d_ph_d_req_tip, tc_p_d_0_d_0_d_ph_d_req_ge, tc_p_d_0_d_0_d_ph_d_req_top);

  tc_tmp_d_118_d_id_d_1_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_118_d_id_d_1_d_cast_d_ack_tip, tc_tmp_d_118_d_id_d_1_d_cast_d_ack_ge, tc_tmp_d_118_d_id_d_1_d_cast_d_ack_top);

  tc_tmp_d_118_d_id_d_1_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_118_d_id_d_1_d_cast_d_req_tip, tc_tmp_d_118_d_id_d_1_d_cast_d_req_ge, tc_tmp_d_118_d_id_d_1_d_cast_d_req_top);

  tc_tmp_d_154_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_154_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_154_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_154_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_154_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_154_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_154_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_154_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_158_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_158_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_158_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_158_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_158_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_158_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_158_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_158_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_163_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_163_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_163_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_163_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_163_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_163_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_163_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_163_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_171_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_171_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_171_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_171_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_171_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_171_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_171_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_171_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_175_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_175_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_175_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_175_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_175_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_175_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_175_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_175_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_179_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_179_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_179_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_179_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_179_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_179_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_179_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_179_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_188_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_188_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_188_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_188_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_188_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_188_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_188_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_188_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_192_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_192_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_192_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_192_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_192_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_192_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_192_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_192_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_206_d_id_d_0_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_206_d_id_d_0_d_cast_d_ack_tip, tc_tmp_d_206_d_id_d_0_d_cast_d_ack_ge, tc_tmp_d_206_d_id_d_0_d_cast_d_ack_top);

  tc_tmp_d_206_d_id_d_0_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_206_d_id_d_0_d_cast_d_req_tip, tc_tmp_d_206_d_id_d_0_d_cast_d_req_ge, tc_tmp_d_206_d_id_d_0_d_cast_d_req_top);

  tc_tmp_d_225_d_id_d_0_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_225_d_id_d_0_d_cast_d_ack_tip, tc_tmp_d_225_d_id_d_0_d_cast_d_ack_ge, tc_tmp_d_225_d_id_d_0_d_cast_d_ack_top);

  tc_tmp_d_225_d_id_d_0_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_225_d_id_d_0_d_cast_d_req_tip, tc_tmp_d_225_d_id_d_0_d_cast_d_req_ge, tc_tmp_d_225_d_id_d_0_d_cast_d_req_top);

  tc_tmp_d_27_d_id_d_1_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_27_d_id_d_1_d_cast_d_ack_tip, tc_tmp_d_27_d_id_d_1_d_cast_d_ack_ge, tc_tmp_d_27_d_id_d_1_d_cast_d_ack_top);

  tc_tmp_d_27_d_id_d_1_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_27_d_id_d_1_d_cast_d_req_tip, tc_tmp_d_27_d_id_d_1_d_cast_d_req_ge, tc_tmp_d_27_d_id_d_1_d_cast_d_req_top);

  tc_tmp_d_27_d_id_d_2_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_27_d_id_d_2_d_cast_d_ack_tip, tc_tmp_d_27_d_id_d_2_d_cast_d_ack_ge, tc_tmp_d_27_d_id_d_2_d_cast_d_ack_top);

  tc_tmp_d_27_d_id_d_2_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_27_d_id_d_2_d_cast_d_req_tip, tc_tmp_d_27_d_id_d_2_d_cast_d_req_ge, tc_tmp_d_27_d_id_d_2_d_cast_d_req_top);

  tc_tmp_d_74_d_id_d_1_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_74_d_id_d_1_d_cast_d_ack_tip, tc_tmp_d_74_d_id_d_1_d_cast_d_ack_ge, tc_tmp_d_74_d_id_d_1_d_cast_d_ack_top);

  tc_tmp_d_74_d_id_d_1_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_74_d_id_d_1_d_cast_d_req_tip, tc_tmp_d_74_d_id_d_1_d_cast_d_req_ge, tc_tmp_d_74_d_id_d_1_d_cast_d_req_top);

  tc_tmp_d_97_d_id_d_1_d_cast_d_ack : transition
  generic map(1)
  port map(tc_tmp_d_97_d_id_d_1_d_cast_d_ack_tip, tc_tmp_d_97_d_id_d_1_d_cast_d_ack_ge, tc_tmp_d_97_d_id_d_1_d_cast_d_ack_top);

  tc_tmp_d_97_d_id_d_1_d_cast_d_req : transition
  generic map(1)
  port map(tc_tmp_d_97_d_id_d_1_d_cast_d_req_tip, tc_tmp_d_97_d_id_d_1_d_cast_d_req_ge, tc_tmp_d_97_d_id_d_1_d_cast_d_req_top);

  then_d_0_d_entry : transition
  generic map(1)
  port map(then_d_0_d_entry_tip, then_d_0_d_entry_ge, then_d_0_d_entry_top);

  then_d_0_to_no_exit_d_4_src : transition
  generic map(1)
  port map(then_d_0_to_no_exit_d_4_src_tip, then_d_0_to_no_exit_d_4_src_ge, then_d_0_to_no_exit_d_4_src_top);

  then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src : transition
  generic map(1)
  port map(then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_tip, then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_ge, then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_top);

  then_d_1_d_entry : transition
  generic map(1)
  port map(then_d_1_d_entry_tip, then_d_1_d_entry_ge, then_d_1_d_entry_top);

  then_d_1_to_loopexit_d_10_src : transition
  generic map(1)
  port map(then_d_1_to_loopexit_d_10_src_tip, then_d_1_to_loopexit_d_10_src_ge, then_d_1_to_loopexit_d_10_src_top);

  then_d_1_to_no_exit_d_10_d_backedge_src : transition
  generic map(1)
  port map(then_d_1_to_no_exit_d_10_d_backedge_src_tip, then_d_1_to_no_exit_d_10_d_backedge_src_ge, then_d_1_to_no_exit_d_10_d_backedge_src_top);

  then_d_2_d_entry : transition
  generic map(1)
  port map(then_d_2_d_entry_tip, then_d_2_d_entry_ge, then_d_2_d_entry_top);

  then_d_2_to_loopexit_d_10_src : transition
  generic map(1)
  port map(then_d_2_to_loopexit_d_10_src_tip, then_d_2_to_loopexit_d_10_src_ge, then_d_2_to_loopexit_d_10_src_top);

  then_d_2_to_no_exit_d_10_d_backedge_src : transition
  generic map(1)
  port map(then_d_2_to_no_exit_d_10_d_backedge_src_tip, then_d_2_to_no_exit_d_10_d_backedge_src_ge, then_d_2_to_no_exit_d_10_d_backedge_src_top);

  place_1_tip(0) <= load_u_array_d_ack_top;
  place_1_rst(0) <= indvar118_d_ph_d_ph_mux_1_d_req0_top;
  place_100_tip(0) <= indvar118_d_ph_d_ph_mux_1_d_req0_top;
  place_100_tip(1) <= indvar118_d_ph_d_ph_mux_1_d_req1_top;
  place_100_rst(0) <= indvar118_d_ph_d_ph_mux_1_d_ack_top;
  place_101_tip(0) <= indvar118_d_ph_d_ph_mux_1_d_ack_top;
  place_101_rst(0) <= indvar_mux_1_d_req1_top;
  place_105_tip(0) <= indvar_mux_1_d_req0_top;
  place_105_tip(1) <= indvar_mux_1_d_req1_top;
  place_105_rst(0) <= indvar_mux_1_d_ack_top;
  place_106_tip(0) <= indvar_mux_1_d_ack_top;
  place_106_rst(0) <= no_exit_d_1_d_entry_top;
  place_107_tip(0) <= no_exit_d_1_to_no_exit_d_1_src_top;
  place_107_rst(0) <= indvar_mux_1_d_req0_top;
  place_108_tip(0) <= oper_tmp_d_11_d_id_d_1_uint_d_req_top;
  place_108_rst(0) <= oper_tmp_d_11_d_id_d_1_uint_d_ack_top;
  place_109_tip(0) <= no_exit_d_1_d_entry_top;
  place_109_rst(0) <= oper_tmp_d_11_d_id_d_1_uint_d_req_top;
  place_110_tip(0) <= oper_tmp_d_11_d_lvl_d_1_uint_d_req_top;
  place_110_rst(0) <= oper_tmp_d_11_d_lvl_d_1_uint_d_ack_top;
  place_111_tip(0) <= oper_tmp_d_11_d_id_d_1_uint_d_ack_top;
  place_111_rst(0) <= oper_tmp_d_11_d_lvl_d_1_uint_d_req_top;
  place_112_tip(0) <= oper_tmp_d_11_d_lvl_d_2_uint_d_req_top;
  place_112_rst(0) <= oper_tmp_d_11_d_lvl_d_2_uint_d_ack_top;
  place_113_tip(0) <= oper_tmp_d_11_d_lvl_d_1_uint_d_ack_top;
  place_113_rst(0) <= oper_tmp_d_11_d_lvl_d_2_uint_d_req_top;
  place_114_tip(0) <= store_0_d_req_top;
  place_114_rst(0) <= store_0_d_ack_top;
  place_115_tip(0) <= oper_tmp_d_11_d_lvl_d_2_uint_d_ack_top;
  place_115_rst(0) <= store_0_d_req_top;
  place_116_tip(0) <= store_0_d_ack_top;
  place_116_rst(0) <= cbr_6_oper_exitcond_bool_d_req_top;
  place_117_tip(0) <= oper_indvar_d_next_uint_d_req_top;
  place_117_rst(0) <= oper_indvar_d_next_uint_d_ack_top;
  place_118_tip(0) <= no_exit_d_1_d_entry_top;
  place_118_rst(0) <= oper_indvar_d_next_uint_d_req_top;
  place_119_tip(0) <= oper_exitcond_bool_d_req_top;
  place_119_rst(0) <= oper_exitcond_bool_d_ack_top;
  place_120_tip(0) <= oper_indvar_d_next_uint_d_ack_top;
  place_120_rst(0) <= oper_exitcond_bool_d_req_top;
  place_121_tip(0) <= oper_exitcond_bool_d_ack_top;
  place_121_rst(0) <= cbr_6_oper_exitcond_bool_d_req_top;
  place_122_tip(0) <= cbr_6_oper_exitcond_bool_d_req_top;
  place_122_rst(0) <= no_exit_d_1_to_loopexit_d_1_src_top;
  place_122_rst(1) <= no_exit_d_1_to_no_exit_d_1_src_top;
  place_123_tip(0) <= store_0_d_ack_top;
  place_123_rst(0) <= cbr_6_oper_exitcond_bool_d_req_top;
  place_124_tip(0) <= oper_indvar_d_next119_uint_d_req_top;
  place_124_rst(0) <= oper_indvar_d_next119_uint_d_ack_top;
  place_126_tip(0) <= oper_exitcond120_bool_d_req_top;
  place_126_rst(0) <= oper_exitcond120_bool_d_ack_top;
  place_127_tip(0) <= oper_indvar_d_next119_uint_d_ack_top;
  place_127_rst(0) <= oper_exitcond120_bool_d_req_top;
  place_128_tip(0) <= oper_exitcond120_bool_d_ack_top;
  place_128_rst(0) <= cbr_7_oper_exitcond120_bool_d_req_top;
  place_129_tip(0) <= cbr_7_oper_exitcond120_bool_d_req_top;
  place_129_rst(0) <= loopexit_d_1_to_loopentry_d_2_src_top;
  place_129_rst(1) <= loopexit_d_1_to_no_exit_d_1_d_outer_src_top;
  place_130_tip(0) <= oper_tmp_d_16_bool_d_req_top;
  place_130_rst(0) <= oper_tmp_d_16_bool_d_ack_top;
  place_132_tip(0) <= oper_tmp_d_16_bool_d_ack_top;
  place_132_rst(0) <= cbr_8_oper_tmp_d_16_bool_d_req_top;
  place_133_tip(0) <= cbr_8_oper_tmp_d_16_bool_d_req_top;
  place_133_rst(0) <= loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_top;
  place_133_rst(1) <= loopentry_d_2_to_no_exit_d_2_d_preheader_src_top;
  place_136_tip(0) <= indvar121_mux_1_d_req0_top;
  place_136_tip(1) <= indvar121_mux_1_d_req1_top;
  place_136_rst(0) <= indvar121_mux_1_d_ack_top;
  place_137_tip(0) <= indvar121_mux_1_d_ack_top;
  place_137_rst(0) <= no_exit_d_2_d_entry_top;
  place_138_tip(0) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_138_rst(0) <= indvar121_mux_1_d_req0_top;
  place_139_tip(0) <= tc_i_d_1_d_0_d_req_top;
  place_139_rst(0) <= tc_i_d_1_d_0_d_ack_top;
  place_14_tip(0) <= loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_top;
  place_14_tip(1) <= no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_top;
  place_14_rst(0) <= loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top;
  place_140_tip(0) <= no_exit_d_2_d_entry_top;
  place_140_rst(0) <= tc_i_d_1_d_0_d_req_top;
  place_141_tip(0) <= oper_tmp_d_20_d_lvl_d_0_uint_d_req_top;
  place_141_rst(0) <= oper_tmp_d_20_d_lvl_d_0_uint_d_ack_top;
  place_142_tip(0) <= no_exit_d_2_d_entry_top;
  place_142_rst(0) <= oper_tmp_d_20_d_lvl_d_0_uint_d_req_top;
  place_143_tip(0) <= load_tmp_d_21_d_req_top;
  place_143_rst(0) <= load_tmp_d_21_d_ack_top;
  place_144_tip(0) <= oper_tmp_d_20_d_lvl_d_0_uint_d_ack_top;
  place_144_rst(0) <= load_tmp_d_21_d_req_top;
  place_145_tip(0) <= oper_tmp_d_25_d_lvl_d_0_uint_d_req_top;
  place_145_rst(0) <= oper_tmp_d_25_d_lvl_d_0_uint_d_ack_top;
  place_146_tip(0) <= no_exit_d_2_d_entry_top;
  place_146_rst(0) <= oper_tmp_d_25_d_lvl_d_0_uint_d_req_top;
  place_147_tip(0) <= load_tmp_d_26_d_req_top;
  place_147_rst(0) <= load_tmp_d_26_d_ack_top;
  place_148_tip(0) <= oper_tmp_d_25_d_lvl_d_0_uint_d_ack_top;
  place_148_rst(0) <= load_tmp_d_26_d_req_top;
  place_149_tip(0) <= load_tmp_d_21_d_ack_top;
  place_149_rst(0) <= load_tmp_d_26_d_req_top;
  place_150_tip(0) <= tc_tmp_d_27_d_id_d_1_d_cast_d_req_top;
  place_150_rst(0) <= tc_tmp_d_27_d_id_d_1_d_cast_d_ack_top;
  place_151_tip(0) <= load_tmp_d_21_d_ack_top;
  place_151_rst(0) <= tc_tmp_d_27_d_id_d_1_d_cast_d_req_top;
  place_152_tip(0) <= oper_tmp_d_27_d_id_d_1_uint_d_req_top;
  place_152_rst(0) <= oper_tmp_d_27_d_id_d_1_uint_d_ack_top;
  place_153_tip(0) <= tc_tmp_d_27_d_id_d_1_d_cast_d_ack_top;
  place_153_rst(0) <= oper_tmp_d_27_d_id_d_1_uint_d_req_top;
  place_154_tip(0) <= oper_tmp_d_27_d_lvl_d_1_uint_d_req_top;
  place_154_rst(0) <= oper_tmp_d_27_d_lvl_d_1_uint_d_ack_top;
  place_155_tip(0) <= oper_tmp_d_27_d_id_d_1_uint_d_ack_top;
  place_155_rst(0) <= oper_tmp_d_27_d_lvl_d_1_uint_d_req_top;
  place_156_tip(0) <= tc_tmp_d_27_d_id_d_2_d_cast_d_req_top;
  place_156_rst(0) <= tc_tmp_d_27_d_id_d_2_d_cast_d_ack_top;
  place_157_tip(0) <= load_tmp_d_26_d_ack_top;
  place_157_rst(0) <= tc_tmp_d_27_d_id_d_2_d_cast_d_req_top;
  place_158_tip(0) <= oper_tmp_d_27_d_lvl_d_2_uint_d_req_top;
  place_158_rst(0) <= oper_tmp_d_27_d_lvl_d_2_uint_d_ack_top;
  place_159_tip(0) <= oper_tmp_d_27_d_lvl_d_1_uint_d_ack_top;
  place_159_rst(0) <= oper_tmp_d_27_d_lvl_d_2_uint_d_req_top;
  place_16_tip(0) <= loopentry_d_4_d_outer_d_pre_top;
  place_16_rst(0) <= loopentry_d_4_d_outer_d_entry_top;
  place_160_tip(0) <= tc_tmp_d_27_d_id_d_2_d_cast_d_ack_top;
  place_160_rst(0) <= oper_tmp_d_27_d_lvl_d_2_uint_d_req_top;
  place_161_tip(0) <= oper_tmp_d_30_d_lvl_d_0_uint_d_req_top;
  place_161_rst(0) <= oper_tmp_d_30_d_lvl_d_0_uint_d_ack_top;
  place_162_tip(0) <= no_exit_d_2_d_entry_top;
  place_162_rst(0) <= oper_tmp_d_30_d_lvl_d_0_uint_d_req_top;
  place_163_tip(0) <= load_tmp_d_31_d_req_top;
  place_163_rst(0) <= load_tmp_d_31_d_ack_top;
  place_164_tip(0) <= oper_tmp_d_30_d_lvl_d_0_uint_d_ack_top;
  place_164_rst(0) <= load_tmp_d_31_d_req_top;
  place_165_tip(0) <= load_tmp_d_26_d_ack_top;
  place_165_rst(0) <= load_tmp_d_31_d_req_top;
  place_166_tip(0) <= store_1_d_req_top;
  place_166_rst(0) <= store_1_d_ack_top;
  place_167_tip(0) <= oper_tmp_d_27_d_lvl_d_2_uint_d_ack_top;
  place_167_rst(0) <= store_1_d_req_top;
  place_168_tip(0) <= load_tmp_d_31_d_ack_top;
  place_168_rst(0) <= store_1_d_req_top;
  place_169_tip(0) <= load_tmp_d_31_d_ack_top;
  place_169_rst(0) <= store_1_d_req_top;
  place_17_tip(0) <= loopentry_d_4_d_pre_top;
  place_17_rst(0) <= loopentry_d_4_d_entry_top;
  place_170_tip(0) <= store_1_d_ack_top;
  place_170_rst(0) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  place_171_tip(0) <= oper_inc_d_2_int_d_req_top;
  place_171_rst(0) <= oper_inc_d_2_int_d_ack_top;
  place_172_tip(0) <= tc_i_d_1_d_0_d_ack_top;
  place_172_rst(0) <= oper_inc_d_2_int_d_req_top;
  place_173_tip(0) <= oper_tmp_d_1614_bool_d_req_top;
  place_173_rst(0) <= oper_tmp_d_1614_bool_d_ack_top;
  place_174_tip(0) <= oper_inc_d_2_int_d_ack_top;
  place_174_rst(0) <= oper_tmp_d_1614_bool_d_req_top;
  place_175_tip(0) <= oper_indvar_d_next122_uint_d_req_top;
  place_175_rst(0) <= oper_indvar_d_next122_uint_d_ack_top;
  place_176_tip(0) <= no_exit_d_2_d_entry_top;
  place_176_rst(0) <= oper_indvar_d_next122_uint_d_req_top;
  place_177_tip(0) <= oper_indvar_d_next122_uint_d_ack_top;
  place_177_rst(0) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  place_178_tip(0) <= oper_tmp_d_1614_bool_d_ack_top;
  place_178_rst(0) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  place_179_tip(0) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  place_179_rst(0) <= no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_top;
  place_179_rst(1) <= no_exit_d_2_to_no_exit_d_2_src_top;
  place_180_tip(0) <= store_1_d_ack_top;
  place_180_rst(0) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  place_183_tip(0) <= loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top;
  place_183_rst(0) <= indvar129_mux_1_d_req1_top;
  place_184_tip(0) <= indvar129_mux_1_d_req0_top;
  place_184_tip(1) <= indvar129_mux_1_d_req1_top;
  place_184_rst(0) <= indvar129_mux_1_d_ack_top;
  place_185_tip(0) <= indvar129_mux_1_d_ack_top;
  place_185_rst(0) <= loopentry_d_4_d_outer_d_pre_top;
  place_186_tip(0) <= loopexit_d_5_to_loopentry_d_4_d_outer_src_top;
  place_186_rst(0) <= indvar129_mux_1_d_req0_top;
  place_187_tip(0) <= loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top;
  place_187_rst(0) <= j_d_3_d_in_d_ph_mux_1_d_req1_top;
  place_188_tip(0) <= j_d_3_d_in_d_ph_mux_1_d_req0_top;
  place_188_tip(1) <= j_d_3_d_in_d_ph_mux_1_d_req1_top;
  place_188_rst(0) <= j_d_3_d_in_d_ph_mux_1_d_ack_top;
  place_189_tip(0) <= j_d_3_d_in_d_ph_mux_1_d_ack_top;
  place_189_rst(0) <= loopentry_d_4_d_outer_d_pre_top;
  place_190_tip(0) <= loopexit_d_5_to_loopentry_d_4_d_outer_src_top;
  place_190_rst(0) <= j_d_3_d_in_d_ph_mux_1_d_req0_top;
  place_191_tip(0) <= loopentry_d_4_d_outer_d_entry_top;
  place_191_rst(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_192_tip(0) <= loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_top;
  place_192_rst(0) <= maxcoeff_d_2_d_ph_mux_1_d_req1_top;
  place_193_tip(0) <= maxcoeff_d_2_d_ph_mux_1_d_req0_top;
  place_193_tip(1) <= maxcoeff_d_2_d_ph_mux_1_d_req1_top;
  place_193_rst(0) <= maxcoeff_d_2_d_ph_mux_1_d_ack_top;
  place_194_tip(0) <= maxcoeff_d_2_d_ph_mux_1_d_ack_top;
  place_194_rst(0) <= loopentry_d_4_d_outer_d_pre_top;
  place_195_tip(0) <= loopexit_d_5_to_loopentry_d_4_d_outer_src_top;
  place_195_rst(0) <= maxcoeff_d_2_d_ph_mux_1_d_req0_top;
  place_196_tip(0) <= loopentry_d_4_d_outer_d_entry_top;
  place_196_rst(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_197_tip(0) <= tc_i_d_2_d_0_d_ph_d_req_top;
  place_197_rst(0) <= tc_i_d_2_d_0_d_ph_d_ack_top;
  place_198_tip(0) <= loopentry_d_4_d_outer_d_entry_top;
  place_198_rst(0) <= tc_i_d_2_d_0_d_ph_d_req_top;
  place_199_tip(0) <= tc_i_d_2_d_0_d_ph_d_ack_top;
  place_199_rst(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_20_tip(0) <= loopentry_d_4_to_no_exit_d_4_d_preheader_src_top;
  place_20_rst(0) <= no_exit_d_4_d_preheader_d_entry_top;
  place_200_tip(0) <= oper_tmp_d_52_d_id_d_1_uint_d_req_top;
  place_200_rst(0) <= oper_tmp_d_52_d_id_d_1_uint_d_ack_top;
  place_201_tip(0) <= loopentry_d_4_d_outer_d_entry_top;
  place_201_rst(0) <= oper_tmp_d_52_d_id_d_1_uint_d_req_top;
  place_202_tip(0) <= oper_tmp_d_52_d_lvl_d_1_uint_d_req_top;
  place_202_rst(0) <= oper_tmp_d_52_d_lvl_d_1_uint_d_ack_top;
  place_203_tip(0) <= oper_tmp_d_52_d_id_d_1_uint_d_ack_top;
  place_203_rst(0) <= oper_tmp_d_52_d_lvl_d_1_uint_d_req_top;
  place_204_tip(0) <= oper_tmp_d_52_d_lvl_d_2_uint_d_req_top;
  place_204_rst(0) <= oper_tmp_d_52_d_lvl_d_2_uint_d_ack_top;
  place_205_tip(0) <= oper_tmp_d_52_d_lvl_d_1_uint_d_ack_top;
  place_205_rst(0) <= oper_tmp_d_52_d_lvl_d_2_uint_d_req_top;
  place_206_tip(0) <= oper_tmp_d_52_d_lvl_d_2_uint_d_ack_top;
  place_206_rst(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_208_tip(0) <= loopentry_d_4_d_loopexit_to_loopentry_d_4_src_top;
  place_208_rst(0) <= j_d_3_d_in_mux_1_d_req1_top;
  place_209_tip(0) <= j_d_3_d_in_mux_1_d_req0_top;
  place_209_tip(1) <= j_d_3_d_in_mux_1_d_req1_top;
  place_209_rst(0) <= j_d_3_d_in_mux_1_d_ack_top;
  place_210_tip(0) <= j_d_3_d_in_mux_1_d_ack_top;
  place_210_rst(0) <= loopentry_d_4_d_pre_top;
  place_211_tip(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_211_rst(0) <= j_d_3_d_in_mux_1_d_req0_top;
  place_212_tip(0) <= loopentry_d_4_d_loopexit_to_loopentry_d_4_src_top;
  place_212_rst(0) <= maxcoeff_d_2_mux_1_d_req1_top;
  place_213_tip(0) <= maxcoeff_d_2_mux_1_d_req0_top;
  place_213_tip(1) <= maxcoeff_d_2_mux_1_d_req1_top;
  place_213_rst(0) <= maxcoeff_d_2_mux_1_d_ack_top;
  place_214_tip(0) <= maxcoeff_d_2_mux_1_d_ack_top;
  place_214_rst(0) <= loopentry_d_4_d_pre_top;
  place_215_tip(0) <= loopentry_d_4_d_outer_to_loopentry_d_4_src_top;
  place_215_rst(0) <= maxcoeff_d_2_mux_1_d_req0_top;
  place_216_tip(0) <= loopentry_d_4_d_entry_top;
  place_216_rst(0) <= cbr_10_oper_tmp_d_42_bool_d_req_top;
  place_217_tip(0) <= oper_j_d_3_int_d_req_top;
  place_217_rst(0) <= oper_j_d_3_int_d_ack_top;
  place_218_tip(0) <= loopentry_d_4_d_entry_top;
  place_218_rst(0) <= oper_j_d_3_int_d_req_top;
  place_219_tip(0) <= oper_tmp_d_42_bool_d_req_top;
  place_219_rst(0) <= oper_tmp_d_42_bool_d_ack_top;
  place_22_tip(0) <= no_exit_d_4_d_pre_top;
  place_22_rst(0) <= no_exit_d_4_d_entry_top;
  place_220_tip(0) <= oper_j_d_3_int_d_ack_top;
  place_220_rst(0) <= oper_tmp_d_42_bool_d_req_top;
  place_221_tip(0) <= oper_tmp_d_42_bool_d_ack_top;
  place_221_rst(0) <= cbr_10_oper_tmp_d_42_bool_d_req_top;
  place_222_tip(0) <= cbr_10_oper_tmp_d_42_bool_d_req_top;
  place_222_rst(0) <= loopentry_d_4_to_no_exit_d_4_d_preheader_src_top;
  place_222_rst(1) <= loopentry_d_4_to_no_exit_d_5_d_preheader_src_top;
  place_223_tip(0) <= tc_j_d_3_d_in_d_req_top;
  place_223_rst(0) <= tc_j_d_3_d_in_d_ack_top;
  place_224_tip(0) <= no_exit_d_4_d_preheader_d_entry_top;
  place_224_rst(0) <= tc_j_d_3_d_in_d_req_top;
  place_225_tip(0) <= load_tmp_d_53_d_req_top;
  place_225_rst(0) <= load_tmp_d_53_d_ack_top;
  place_226_tip(0) <= no_exit_d_4_d_preheader_d_entry_top;
  place_226_rst(0) <= load_tmp_d_53_d_req_top;
  place_227_tip(0) <= load_tmp_d_53_d_ack_top;
  place_227_rst(0) <= no_exit_d_4_d_preheader_to_no_exit_d_4_src_top;
  place_228_tip(0) <= oper_tmp_d_uint_d_req_top;
  place_228_rst(0) <= oper_tmp_d_uint_d_ack_top;
  place_229_tip(0) <= tc_j_d_3_d_in_d_ack_top;
  place_229_rst(0) <= oper_tmp_d_uint_d_req_top;
  place_230_tip(0) <= oper_tmp_d_uint_d_ack_top;
  place_230_rst(0) <= no_exit_d_4_d_preheader_to_no_exit_d_4_src_top;
  place_231_tip(0) <= then_d_0_to_no_exit_d_4_src_top;
  place_231_rst(0) <= indvar123_mux_1_d_req1_top;
  place_232_tip(0) <= indvar123_mux_1_d_req0_top;
  place_232_tip(1) <= indvar123_mux_1_d_req1_top;
  place_232_rst(0) <= indvar123_mux_1_d_ack_top;
  place_233_tip(0) <= indvar123_mux_1_d_ack_top;
  place_233_rst(0) <= no_exit_d_4_d_pre_top;
  place_234_tip(0) <= no_exit_d_4_d_preheader_to_no_exit_d_4_src_top;
  place_234_rst(0) <= indvar123_mux_1_d_req0_top;
  place_235_tip(0) <= then_d_0_to_no_exit_d_4_src_top;
  place_235_rst(0) <= maxcoeff_d_2_d_2_mux_1_d_req1_top;
  place_236_tip(0) <= maxcoeff_d_2_d_2_mux_1_d_req0_top;
  place_236_tip(1) <= maxcoeff_d_2_d_2_mux_1_d_req1_top;
  place_236_rst(0) <= maxcoeff_d_2_d_2_mux_1_d_ack_top;
  place_237_tip(0) <= maxcoeff_d_2_d_2_mux_1_d_ack_top;
  place_237_rst(0) <= no_exit_d_4_d_pre_top;
  place_238_tip(0) <= no_exit_d_4_d_preheader_to_no_exit_d_4_src_top;
  place_238_rst(0) <= maxcoeff_d_2_d_2_mux_1_d_req0_top;
  place_239_tip(0) <= no_exit_d_4_d_entry_top;
  place_239_rst(0) <= cbr_11_oper_tmp_d_54_bool_d_req_top;
  place_24_tip(0) <= no_exit_d_4_to_then_d_0_src_top;
  place_24_rst(0) <= then_d_0_d_entry_top;
  place_240_tip(0) <= oper_tmp_d_125_uint_d_req_top;
  place_240_rst(0) <= oper_tmp_d_125_uint_d_ack_top;
  place_241_tip(0) <= no_exit_d_4_d_entry_top;
  place_241_rst(0) <= oper_tmp_d_125_uint_d_req_top;
  place_242_tip(0) <= tc_j_d_3_d_2_d_req_top;
  place_242_rst(0) <= tc_j_d_3_d_2_d_ack_top;
  place_243_tip(0) <= oper_tmp_d_125_uint_d_ack_top;
  place_243_rst(0) <= tc_j_d_3_d_2_d_req_top;
  place_244_tip(0) <= tc_j_d_3_d_2_d_ack_top;
  place_244_rst(0) <= cbr_11_oper_tmp_d_54_bool_d_req_top;
  place_245_tip(0) <= oper_tmp_d_47_d_id_d_1_uint_d_req_top;
  place_245_rst(0) <= oper_tmp_d_47_d_id_d_1_uint_d_ack_top;
  place_246_tip(0) <= oper_tmp_d_125_uint_d_ack_top;
  place_246_rst(0) <= oper_tmp_d_47_d_id_d_1_uint_d_req_top;
  place_247_tip(0) <= oper_tmp_d_47_d_lvl_d_1_uint_d_req_top;
  place_247_rst(0) <= oper_tmp_d_47_d_lvl_d_1_uint_d_ack_top;
  place_248_tip(0) <= oper_tmp_d_47_d_id_d_1_uint_d_ack_top;
  place_248_rst(0) <= oper_tmp_d_47_d_lvl_d_1_uint_d_req_top;
  place_249_tip(0) <= oper_tmp_d_47_d_lvl_d_2_uint_d_req_top;
  place_249_rst(0) <= oper_tmp_d_47_d_lvl_d_2_uint_d_ack_top;
  place_25_tip(0) <= no_exit_d_4_to_loopentry_d_4_d_loopexit_src_top;
  place_25_rst(0) <= loopentry_d_4_d_loopexit_to_loopentry_d_4_src_top;
  place_250_tip(0) <= oper_tmp_d_47_d_lvl_d_1_uint_d_ack_top;
  place_250_rst(0) <= oper_tmp_d_47_d_lvl_d_2_uint_d_req_top;
  place_251_tip(0) <= load_tmp_d_48_d_req_top;
  place_251_rst(0) <= load_tmp_d_48_d_ack_top;
  place_252_tip(0) <= oper_tmp_d_47_d_lvl_d_2_uint_d_ack_top;
  place_252_rst(0) <= load_tmp_d_48_d_req_top;
  place_253_tip(0) <= oper_tmp_d_54_bool_d_req_top;
  place_253_rst(0) <= oper_tmp_d_54_bool_d_ack_top;
  place_254_tip(0) <= load_tmp_d_48_d_ack_top;
  place_254_rst(0) <= oper_tmp_d_54_bool_d_req_top;
  place_255_tip(0) <= oper_tmp_d_54_bool_d_ack_top;
  place_255_rst(0) <= cbr_11_oper_tmp_d_54_bool_d_req_top;
  place_256_tip(0) <= cbr_11_oper_tmp_d_54_bool_d_req_top;
  place_256_rst(0) <= no_exit_d_4_to_loopentry_d_4_d_loopexit_src_top;
  place_256_rst(1) <= no_exit_d_4_to_then_d_0_src_top;
  place_257_tip(0) <= oper_j_d_321_int_d_req_top;
  place_257_rst(0) <= oper_j_d_321_int_d_ack_top;
  place_258_tip(0) <= then_d_0_d_entry_top;
  place_258_rst(0) <= oper_j_d_321_int_d_req_top;
  place_259_tip(0) <= oper_tmp_d_4223_bool_d_req_top;
  place_259_rst(0) <= oper_tmp_d_4223_bool_d_ack_top;
  place_260_tip(0) <= oper_j_d_321_int_d_ack_top;
  place_260_rst(0) <= oper_tmp_d_4223_bool_d_req_top;
  place_261_tip(0) <= oper_indvar_d_next124_uint_d_req_top;
  place_261_rst(0) <= oper_indvar_d_next124_uint_d_ack_top;
  place_262_tip(0) <= then_d_0_d_entry_top;
  place_262_rst(0) <= oper_indvar_d_next124_uint_d_req_top;
  place_263_tip(0) <= oper_indvar_d_next124_uint_d_ack_top;
  place_263_rst(0) <= cbr_12_oper_tmp_d_4223_bool_d_req_top;
  place_264_tip(0) <= oper_tmp_d_4223_bool_d_ack_top;
  place_264_rst(0) <= cbr_12_oper_tmp_d_4223_bool_d_req_top;
  place_265_tip(0) <= cbr_12_oper_tmp_d_4223_bool_d_req_top;
  place_265_rst(0) <= then_d_0_to_no_exit_d_4_src_top;
  place_265_rst(1) <= then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_top;
  place_268_tip(0) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_top;
  place_268_tip(1) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_top;
  place_268_rst(0) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_top;
  place_269_tip(0) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_top;
  place_269_rst(0) <= indvar126_mux_1_d_req1_top;
  place_27_tip(0) <= then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_top;
  place_27_rst(0) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_top;
  place_270_tip(0) <= loopentry_d_4_to_no_exit_d_5_d_preheader_src_top;
  place_270_rst(0) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_top;
  place_273_tip(0) <= indvar126_mux_1_d_req0_top;
  place_273_tip(1) <= indvar126_mux_1_d_req1_top;
  place_273_rst(0) <= indvar126_mux_1_d_ack_top;
  place_274_tip(0) <= indvar126_mux_1_d_ack_top;
  place_274_rst(0) <= no_exit_d_5_d_entry_top;
  place_275_tip(0) <= no_exit_d_5_to_no_exit_d_5_src_top;
  place_275_rst(0) <= indvar126_mux_1_d_req0_top;
  place_276_tip(0) <= oper_tmp_d_65_d_id_d_1_uint_d_req_top;
  place_276_rst(0) <= oper_tmp_d_65_d_id_d_1_uint_d_ack_top;
  place_277_tip(0) <= no_exit_d_5_d_entry_top;
  place_277_rst(0) <= oper_tmp_d_65_d_id_d_1_uint_d_req_top;
  place_278_tip(0) <= oper_tmp_d_65_d_lvl_d_1_uint_d_req_top;
  place_278_rst(0) <= oper_tmp_d_65_d_lvl_d_1_uint_d_ack_top;
  place_279_tip(0) <= oper_tmp_d_65_d_id_d_1_uint_d_ack_top;
  place_279_rst(0) <= oper_tmp_d_65_d_lvl_d_1_uint_d_req_top;
  place_280_tip(0) <= oper_tmp_d_65_d_lvl_d_2_uint_d_req_top;
  place_280_rst(0) <= oper_tmp_d_65_d_lvl_d_2_uint_d_ack_top;
  place_281_tip(0) <= oper_tmp_d_65_d_lvl_d_1_uint_d_ack_top;
  place_281_rst(0) <= oper_tmp_d_65_d_lvl_d_2_uint_d_req_top;
  place_282_tip(0) <= load_tmp_d_66_d_req_top;
  place_282_rst(0) <= load_tmp_d_66_d_ack_top;
  place_283_tip(0) <= oper_tmp_d_65_d_lvl_d_2_uint_d_ack_top;
  place_283_rst(0) <= load_tmp_d_66_d_req_top;
  place_284_tip(0) <= tc_tmp_d_74_d_id_d_1_d_cast_d_req_top;
  place_284_rst(0) <= tc_tmp_d_74_d_id_d_1_d_cast_d_ack_top;
  place_285_tip(0) <= no_exit_d_5_d_entry_top;
  place_285_rst(0) <= tc_tmp_d_74_d_id_d_1_d_cast_d_req_top;
  place_286_tip(0) <= oper_tmp_d_74_d_id_d_1_uint_d_req_top;
  place_286_rst(0) <= oper_tmp_d_74_d_id_d_1_uint_d_ack_top;
  place_287_tip(0) <= tc_tmp_d_74_d_id_d_1_d_cast_d_ack_top;
  place_287_rst(0) <= oper_tmp_d_74_d_id_d_1_uint_d_req_top;
  place_288_tip(0) <= oper_tmp_d_74_d_lvl_d_1_uint_d_req_top;
  place_288_rst(0) <= oper_tmp_d_74_d_lvl_d_1_uint_d_ack_top;
  place_289_tip(0) <= oper_tmp_d_74_d_id_d_1_uint_d_ack_top;
  place_289_rst(0) <= oper_tmp_d_74_d_lvl_d_1_uint_d_req_top;
  place_290_tip(0) <= oper_tmp_d_74_d_lvl_d_2_uint_d_req_top;
  place_290_rst(0) <= oper_tmp_d_74_d_lvl_d_2_uint_d_ack_top;
  place_291_tip(0) <= oper_tmp_d_74_d_lvl_d_1_uint_d_ack_top;
  place_291_rst(0) <= oper_tmp_d_74_d_lvl_d_2_uint_d_req_top;
  place_292_tip(0) <= load_tmp_d_75_d_req_top;
  place_292_rst(0) <= load_tmp_d_75_d_ack_top;
  place_293_tip(0) <= oper_tmp_d_74_d_lvl_d_2_uint_d_ack_top;
  place_293_rst(0) <= load_tmp_d_75_d_req_top;
  place_294_tip(0) <= load_tmp_d_66_d_ack_top;
  place_294_rst(0) <= load_tmp_d_75_d_req_top;
  place_295_tip(0) <= store_2_d_req_top;
  place_295_rst(0) <= store_2_d_ack_top;
  place_296_tip(0) <= oper_tmp_d_65_d_lvl_d_2_uint_d_ack_top;
  place_296_rst(0) <= store_2_d_req_top;
  place_297_tip(0) <= load_tmp_d_75_d_ack_top;
  place_297_rst(0) <= store_2_d_req_top;
  place_298_tip(0) <= load_tmp_d_75_d_ack_top;
  place_298_rst(0) <= store_2_d_req_top;
  place_299_tip(0) <= store_2_d_ack_top;
  place_299_rst(0) <= cbr_13_oper_exitcond128_bool_d_req_top;
  place_30_tip(0) <= no_exit_d_5_to_loopexit_d_5_src_top;
  place_30_rst(0) <= loopexit_d_5_d_entry_top;
  place_300_tip(0) <= store_3_d_req_top;
  place_300_rst(0) <= store_3_d_ack_top;
  place_301_tip(0) <= oper_tmp_d_74_d_lvl_d_2_uint_d_ack_top;
  place_301_rst(0) <= store_3_d_req_top;
  place_302_tip(0) <= load_tmp_d_66_d_ack_top;
  place_302_rst(0) <= store_3_d_req_top;
  place_303_tip(0) <= store_2_d_ack_top;
  place_303_rst(0) <= store_3_d_req_top;
  place_304_tip(0) <= store_3_d_ack_top;
  place_304_rst(0) <= cbr_13_oper_exitcond128_bool_d_req_top;
  place_305_tip(0) <= oper_indvar_d_next127_uint_d_req_top;
  place_305_rst(0) <= oper_indvar_d_next127_uint_d_ack_top;
  place_306_tip(0) <= no_exit_d_5_d_entry_top;
  place_306_rst(0) <= oper_indvar_d_next127_uint_d_req_top;
  place_307_tip(0) <= oper_exitcond128_bool_d_req_top;
  place_307_rst(0) <= oper_exitcond128_bool_d_ack_top;
  place_308_tip(0) <= oper_indvar_d_next127_uint_d_ack_top;
  place_308_rst(0) <= oper_exitcond128_bool_d_req_top;
  place_309_tip(0) <= oper_exitcond128_bool_d_ack_top;
  place_309_rst(0) <= cbr_13_oper_exitcond128_bool_d_req_top;
  place_310_tip(0) <= cbr_13_oper_exitcond128_bool_d_req_top;
  place_310_rst(0) <= no_exit_d_5_to_loopexit_d_5_src_top;
  place_310_rst(1) <= no_exit_d_5_to_no_exit_d_5_src_top;
  place_311_tip(0) <= store_3_d_ack_top;
  place_311_rst(0) <= cbr_13_oper_exitcond128_bool_d_req_top;
  place_312_tip(0) <= oper_inc_d_5_int_d_req_top;
  place_312_rst(0) <= oper_inc_d_5_int_d_ack_top;
  place_313_tip(0) <= loopexit_d_5_d_entry_top;
  place_313_rst(0) <= oper_inc_d_5_int_d_req_top;
  place_314_tip(0) <= oper_inc_d_5_int_d_ack_top;
  place_314_rst(0) <= cbr_14_oper_exitcond131_bool_d_req_top;
  place_315_tip(0) <= oper_indvar_d_next130_uint_d_req_top;
  place_315_rst(0) <= oper_indvar_d_next130_uint_d_ack_top;
  place_316_tip(0) <= loopexit_d_5_d_entry_top;
  place_316_rst(0) <= oper_indvar_d_next130_uint_d_req_top;
  place_317_tip(0) <= oper_exitcond131_bool_d_req_top;
  place_317_rst(0) <= oper_exitcond131_bool_d_ack_top;
  place_318_tip(0) <= oper_indvar_d_next130_uint_d_ack_top;
  place_318_rst(0) <= oper_exitcond131_bool_d_req_top;
  place_319_tip(0) <= oper_exitcond131_bool_d_ack_top;
  place_319_rst(0) <= cbr_14_oper_exitcond131_bool_d_req_top;
  place_32_tip(0) <= loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_top;
  place_32_rst(0) <= loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_top;
  place_320_tip(0) <= cbr_14_oper_exitcond131_bool_d_req_top;
  place_320_rst(0) <= loopexit_d_5_to_loopentry_d_4_d_outer_src_top;
  place_320_rst(1) <= loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_top;
  place_322_tip(0) <= loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_top;
  place_322_rst(0) <= indvar134_mux_1_d_req1_top;
  place_323_tip(0) <= indvar134_mux_1_d_req0_top;
  place_323_tip(1) <= indvar134_mux_1_d_req1_top;
  place_323_rst(0) <= indvar134_mux_1_d_ack_top;
  place_324_tip(0) <= indvar134_mux_1_d_ack_top;
  place_324_rst(0) <= loopentry_d_7_d_outer_d_pre_top;
  place_325_tip(0) <= loopexit_d_7_to_loopentry_d_7_d_outer_src_top;
  place_325_rst(0) <= indvar134_mux_1_d_req0_top;
  place_326_tip(0) <= loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_top;
  place_326_rst(0) <= k_d_1_d_in_d_ph_mux_1_d_req1_top;
  place_327_tip(0) <= k_d_1_d_in_d_ph_mux_1_d_req0_top;
  place_327_tip(1) <= k_d_1_d_in_d_ph_mux_1_d_req1_top;
  place_327_rst(0) <= k_d_1_d_in_d_ph_mux_1_d_ack_top;
  place_328_tip(0) <= k_d_1_d_in_d_ph_mux_1_d_ack_top;
  place_328_rst(0) <= loopentry_d_7_d_outer_d_pre_top;
  place_329_tip(0) <= loopexit_d_7_to_loopentry_d_7_d_outer_src_top;
  place_329_rst(0) <= k_d_1_d_in_d_ph_mux_1_d_req0_top;
  place_33_tip(0) <= loopentry_d_7_d_outer_d_pre_top;
  place_33_rst(0) <= loopentry_d_7_d_outer_d_entry_top;
  place_330_tip(0) <= loopentry_d_7_d_outer_d_entry_top;
  place_330_rst(0) <= loopentry_d_7_d_outer_to_loopentry_d_7_src_top;
  place_331_tip(0) <= tc_p_d_0_d_0_d_ph_d_req_top;
  place_331_rst(0) <= tc_p_d_0_d_0_d_ph_d_ack_top;
  place_332_tip(0) <= loopentry_d_7_d_outer_d_entry_top;
  place_332_rst(0) <= tc_p_d_0_d_0_d_ph_d_req_top;
  place_333_tip(0) <= oper_tmp_d_107_d_id_d_1_uint_d_req_top;
  place_333_rst(0) <= oper_tmp_d_107_d_id_d_1_uint_d_ack_top;
  place_334_tip(0) <= loopentry_d_7_d_outer_d_entry_top;
  place_334_rst(0) <= oper_tmp_d_107_d_id_d_1_uint_d_req_top;
  place_335_tip(0) <= oper_tmp_d_107_d_lvl_d_1_uint_d_req_top;
  place_335_rst(0) <= oper_tmp_d_107_d_lvl_d_1_uint_d_ack_top;
  place_336_tip(0) <= oper_tmp_d_107_d_id_d_1_uint_d_ack_top;
  place_336_rst(0) <= oper_tmp_d_107_d_lvl_d_1_uint_d_req_top;
  place_337_tip(0) <= oper_tmp_d_107_d_lvl_d_2_uint_d_req_top;
  place_337_rst(0) <= oper_tmp_d_107_d_lvl_d_2_uint_d_ack_top;
  place_338_tip(0) <= oper_tmp_d_107_d_lvl_d_1_uint_d_ack_top;
  place_338_rst(0) <= oper_tmp_d_107_d_lvl_d_2_uint_d_req_top;
  place_339_tip(0) <= oper_tmp_d_107_d_lvl_d_2_uint_d_ack_top;
  place_339_rst(0) <= loopentry_d_7_d_outer_to_loopentry_d_7_src_top;
  place_340_tip(0) <= oper_j_d_746_int_d_req_top;
  place_340_rst(0) <= oper_j_d_746_int_d_ack_top;
  place_341_tip(0) <= tc_p_d_0_d_0_d_ph_d_ack_top;
  place_341_rst(0) <= oper_j_d_746_int_d_req_top;
  place_342_tip(0) <= oper_tmp_d_11348_bool_d_req_top;
  place_342_rst(0) <= oper_tmp_d_11348_bool_d_ack_top;
  place_343_tip(0) <= oper_j_d_746_int_d_ack_top;
  place_343_rst(0) <= oper_tmp_d_11348_bool_d_req_top;
  place_344_tip(0) <= oper_tmp_d_11348_bool_d_ack_top;
  place_344_rst(0) <= loopentry_d_7_d_outer_to_loopentry_d_7_src_top;
  place_345_tip(0) <= oper_tmp_d_136_uint_d_req_top;
  place_345_rst(0) <= oper_tmp_d_136_uint_d_ack_top;
  place_346_tip(0) <= loopentry_d_7_d_outer_d_entry_top;
  place_346_rst(0) <= oper_tmp_d_136_uint_d_req_top;
  place_347_tip(0) <= oper_tmp_d_136_uint_d_ack_top;
  place_347_rst(0) <= loopentry_d_7_d_outer_to_loopentry_d_7_src_top;
  place_349_tip(0) <= indvar138_mux_1_d_req0_top;
  place_349_tip(1) <= indvar138_mux_1_d_req1_top;
  place_349_rst(0) <= indvar138_mux_1_d_ack_top;
  place_350_tip(0) <= indvar138_mux_1_d_ack_top;
  place_350_rst(0) <= tc_indvar138_d_req_top;
  place_351_tip(0) <= loopentry_d_7_d_outer_to_loopentry_d_7_src_top;
  place_351_rst(0) <= indvar138_mux_1_d_req0_top;
  place_352_tip(0) <= tc_indvar138_d_req_top;
  place_352_rst(0) <= tc_indvar138_d_ack_top;
  place_354_tip(0) <= oper_k_d_1_d_in_int_d_req_top;
  place_354_rst(0) <= oper_k_d_1_d_in_int_d_ack_top;
  place_355_tip(0) <= tc_indvar138_d_ack_top;
  place_355_rst(0) <= oper_k_d_1_d_in_int_d_req_top;
  place_356_tip(0) <= oper_k_d_1_int_d_req_top;
  place_356_rst(0) <= oper_k_d_1_int_d_ack_top;
  place_357_tip(0) <= oper_k_d_1_d_in_int_d_ack_top;
  place_357_rst(0) <= oper_k_d_1_int_d_req_top;
  place_358_tip(0) <= oper_tmp_d_92_bool_d_req_top;
  place_358_rst(0) <= oper_tmp_d_92_bool_d_ack_top;
  place_359_tip(0) <= oper_k_d_1_int_d_ack_top;
  place_359_rst(0) <= oper_tmp_d_92_bool_d_req_top;
  place_36_tip(0) <= loopentry_d_7_to_no_exit_d_7_src_top;
  place_36_rst(0) <= no_exit_d_7_d_entry_top;
  place_360_tip(0) <= oper_tmp_d_92_bool_d_ack_top;
  place_360_rst(0) <= cbr_15_oper_tmp_d_92_bool_d_req_top;
  place_361_tip(0) <= cbr_15_oper_tmp_d_92_bool_d_req_top;
  place_361_rst(0) <= loopentry_d_7_to_loopexit_d_7_src_top;
  place_361_rst(1) <= loopentry_d_7_to_no_exit_d_7_src_top;
  place_362_tip(0) <= tc_tmp_d_97_d_id_d_1_d_cast_d_req_top;
  place_362_rst(0) <= tc_tmp_d_97_d_id_d_1_d_cast_d_ack_top;
  place_363_tip(0) <= no_exit_d_7_d_entry_top;
  place_363_rst(0) <= tc_tmp_d_97_d_id_d_1_d_cast_d_req_top;
  place_364_tip(0) <= oper_tmp_d_97_d_id_d_1_uint_d_req_top;
  place_364_rst(0) <= oper_tmp_d_97_d_id_d_1_uint_d_ack_top;
  place_365_tip(0) <= tc_tmp_d_97_d_id_d_1_d_cast_d_ack_top;
  place_365_rst(0) <= oper_tmp_d_97_d_id_d_1_uint_d_req_top;
  place_366_tip(0) <= oper_tmp_d_97_d_lvl_d_1_uint_d_req_top;
  place_366_rst(0) <= oper_tmp_d_97_d_lvl_d_1_uint_d_ack_top;
  place_367_tip(0) <= oper_tmp_d_97_d_id_d_1_uint_d_ack_top;
  place_367_rst(0) <= oper_tmp_d_97_d_lvl_d_1_uint_d_req_top;
  place_368_tip(0) <= oper_tmp_d_97_d_lvl_d_2_uint_d_req_top;
  place_368_rst(0) <= oper_tmp_d_97_d_lvl_d_2_uint_d_ack_top;
  place_369_tip(0) <= oper_tmp_d_97_d_lvl_d_1_uint_d_ack_top;
  place_369_rst(0) <= oper_tmp_d_97_d_lvl_d_2_uint_d_req_top;
  place_370_tip(0) <= load_tmp_d_103_d_req_top;
  place_370_rst(0) <= load_tmp_d_103_d_ack_top;
  place_371_tip(0) <= oper_tmp_d_97_d_lvl_d_2_uint_d_ack_top;
  place_371_rst(0) <= load_tmp_d_103_d_req_top;
  place_372_tip(0) <= load_tmp_d_108_d_req_top;
  place_372_rst(0) <= load_tmp_d_108_d_ack_top;
  place_373_tip(0) <= load_tmp_d_103_d_ack_top;
  place_373_rst(0) <= load_tmp_d_108_d_req_top;
  place_374_tip(0) <= no_exit_d_7_d_entry_top;
  place_374_rst(0) <= load_tmp_d_108_d_req_top;
  place_375_tip(0) <= start_call_divide_0_d_req_top;
  place_375_rst(0) <= start_call_divide_0_d_ack_top;
  place_376_tip(0) <= load_tmp_d_103_d_ack_top;
  place_376_rst(0) <= start_call_divide_0_actual_0_wr_d_req_top;
  place_377_tip(0) <= load_tmp_d_108_d_ack_top;
  place_377_rst(0) <= start_call_divide_0_actual_0_wr_d_req_top;
  place_378_tip(0) <= start_call_divide_0_actual_0_wr_d_req_top;
  place_378_rst(0) <= start_call_divide_0_actual_0_wr_d_ack_top;
  place_379_tip(0) <= load_tmp_d_108_d_ack_top;
  place_379_rst(0) <= start_call_divide_0_actual_1_wr_d_req_top;
  place_38_tip(0) <= loopentry_d_7_to_loopexit_d_7_src_top;
  place_38_rst(0) <= oper_exitcond142_bool_d_req_top;
  place_380_tip(0) <= start_call_divide_0_actual_0_wr_d_ack_top;
  place_380_rst(0) <= start_call_divide_0_actual_1_wr_d_req_top;
  place_381_tip(0) <= start_call_divide_0_actual_1_wr_d_req_top;
  place_381_rst(0) <= start_call_divide_0_actual_1_wr_d_ack_top;
  place_382_tip(0) <= start_call_divide_0_actual_1_wr_d_ack_top;
  place_382_rst(0) <= start_call_divide_0_d_req_top;
  place_383_tip(0) <= start_call_divide_0_d_ack_top;
  place_383_rst(0) <= load_start_call_divide_0_return_d_req_top;
  place_384_tip(0) <= load_start_call_divide_0_return_d_req_top;
  place_384_rst(0) <= load_start_call_divide_0_return_d_ack_top;
  place_385_tip(0) <= store_4_d_req_top;
  place_385_rst(0) <= store_4_d_ack_top;
  place_386_tip(0) <= oper_tmp_d_97_d_lvl_d_2_uint_d_ack_top;
  place_386_rst(0) <= store_4_d_req_top;
  place_387_tip(0) <= load_start_call_divide_0_return_d_ack_top;
  place_387_rst(0) <= store_4_d_req_top;
  place_388_tip(0) <= load_start_call_divide_0_return_d_ack_top;
  place_388_rst(0) <= store_4_d_req_top;
  place_389_tip(0) <= store_4_d_ack_top;
  place_389_rst(0) <= cbr_16_oper_tmp_d_11348_bool_d_req_top;
  place_390_tip(0) <= no_exit_d_7_d_entry_top;
  place_390_rst(0) <= cbr_16_oper_tmp_d_11348_bool_d_req_top;
  place_391_tip(0) <= cbr_16_oper_tmp_d_11348_bool_d_req_top;
  place_391_rst(0) <= no_exit_d_7_to_loopentry_d_7_d_backedge_src_top;
  place_391_rst(1) <= no_exit_d_7_to_no_exit_d_8_d_preheader_src_top;
  place_392_tip(0) <= store_4_d_ack_top;
  place_392_rst(0) <= cbr_16_oper_tmp_d_11348_bool_d_req_top;
  place_394_tip(0) <= oper_indvar_d_next139_uint_d_req_top;
  place_394_rst(0) <= oper_indvar_d_next139_uint_d_ack_top;
  place_396_tip(0) <= oper_indvar_d_next139_uint_d_ack_top;
  place_396_rst(0) <= indvar138_mux_1_d_req1_top;
  place_399_tip(0) <= indvar132_mux_1_d_req0_top;
  place_399_tip(1) <= indvar132_mux_1_d_req1_top;
  place_399_rst(0) <= indvar132_mux_1_d_ack_top;
  place_40_tip(0) <= no_exit_d_7_to_no_exit_d_8_d_preheader_src_top;
  place_40_rst(0) <= indvar132_mux_1_d_req1_top;
  place_400_tip(0) <= indvar132_mux_1_d_ack_top;
  place_400_rst(0) <= no_exit_d_8_d_entry_top;
  place_401_tip(0) <= no_exit_d_8_to_no_exit_d_8_src_top;
  place_401_rst(0) <= indvar132_mux_1_d_req0_top;
  place_402_tip(0) <= oper_tmp_d_137_uint_d_req_top;
  place_402_rst(0) <= oper_tmp_d_137_uint_d_ack_top;
  place_403_tip(0) <= no_exit_d_8_d_entry_top;
  place_403_rst(0) <= oper_tmp_d_137_uint_d_req_top;
  place_404_tip(0) <= tc_j_d_7_d_1_d_req_top;
  place_404_rst(0) <= tc_j_d_7_d_1_d_ack_top;
  place_405_tip(0) <= oper_tmp_d_137_uint_d_ack_top;
  place_405_rst(0) <= tc_j_d_7_d_1_d_req_top;
  place_406_tip(0) <= tc_tmp_d_118_d_id_d_1_d_cast_d_req_top;
  place_406_rst(0) <= tc_tmp_d_118_d_id_d_1_d_cast_d_ack_top;
  place_407_tip(0) <= no_exit_d_8_d_entry_top;
  place_407_rst(0) <= tc_tmp_d_118_d_id_d_1_d_cast_d_req_top;
  place_408_tip(0) <= oper_tmp_d_118_d_id_d_1_uint_d_req_top;
  place_408_rst(0) <= oper_tmp_d_118_d_id_d_1_uint_d_ack_top;
  place_409_tip(0) <= tc_tmp_d_118_d_id_d_1_d_cast_d_ack_top;
  place_409_rst(0) <= oper_tmp_d_118_d_id_d_1_uint_d_req_top;
  place_410_tip(0) <= oper_tmp_d_118_d_lvl_d_1_uint_d_req_top;
  place_410_rst(0) <= oper_tmp_d_118_d_lvl_d_1_uint_d_ack_top;
  place_411_tip(0) <= oper_tmp_d_118_d_id_d_1_uint_d_ack_top;
  place_411_rst(0) <= oper_tmp_d_118_d_lvl_d_1_uint_d_req_top;
  place_412_tip(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_req_top;
  place_412_rst(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_ack_top;
  place_413_tip(0) <= oper_tmp_d_118_d_lvl_d_1_uint_d_ack_top;
  place_413_rst(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_req_top;
  place_414_tip(0) <= oper_tmp_d_137_uint_d_ack_top;
  place_414_rst(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_req_top;
  place_415_tip(0) <= load_tmp_d_123_d_req_top;
  place_415_rst(0) <= load_tmp_d_123_d_ack_top;
  place_416_tip(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_ack_top;
  place_416_rst(0) <= load_tmp_d_123_d_req_top;
  place_417_tip(0) <= load_tmp_d_128_d_req_top;
  place_417_rst(0) <= load_tmp_d_128_d_ack_top;
  place_418_tip(0) <= load_tmp_d_123_d_ack_top;
  place_418_rst(0) <= load_tmp_d_128_d_req_top;
  place_419_tip(0) <= no_exit_d_8_d_entry_top;
  place_419_rst(0) <= load_tmp_d_128_d_req_top;
  place_420_tip(0) <= oper_tmp_d_132_d_id_d_1_uint_d_req_top;
  place_420_rst(0) <= oper_tmp_d_132_d_id_d_1_uint_d_ack_top;
  place_421_tip(0) <= no_exit_d_8_d_entry_top;
  place_421_rst(0) <= oper_tmp_d_132_d_id_d_1_uint_d_req_top;
  place_422_tip(0) <= oper_tmp_d_132_d_lvl_d_1_uint_d_req_top;
  place_422_rst(0) <= oper_tmp_d_132_d_lvl_d_1_uint_d_ack_top;
  place_423_tip(0) <= oper_tmp_d_132_d_id_d_1_uint_d_ack_top;
  place_423_rst(0) <= oper_tmp_d_132_d_lvl_d_1_uint_d_req_top;
  place_424_tip(0) <= oper_tmp_d_132_d_lvl_d_2_uint_d_req_top;
  place_424_rst(0) <= oper_tmp_d_132_d_lvl_d_2_uint_d_ack_top;
  place_425_tip(0) <= oper_tmp_d_132_d_lvl_d_1_uint_d_ack_top;
  place_425_rst(0) <= oper_tmp_d_132_d_lvl_d_2_uint_d_req_top;
  place_426_tip(0) <= oper_tmp_d_137_uint_d_ack_top;
  place_426_rst(0) <= oper_tmp_d_132_d_lvl_d_2_uint_d_req_top;
  place_427_tip(0) <= load_tmp_d_133_d_req_top;
  place_427_rst(0) <= load_tmp_d_133_d_ack_top;
  place_428_tip(0) <= oper_tmp_d_132_d_lvl_d_2_uint_d_ack_top;
  place_428_rst(0) <= load_tmp_d_133_d_req_top;
  place_429_tip(0) <= load_tmp_d_128_d_ack_top;
  place_429_rst(0) <= load_tmp_d_133_d_req_top;
  place_430_tip(0) <= oper_tmp_d_134_float_d_req_top;
  place_430_rst(0) <= oper_tmp_d_134_float_d_ack_top;
  place_431_tip(0) <= load_tmp_d_128_d_ack_top;
  place_431_rst(0) <= oper_tmp_d_134_float_d_req_top;
  place_432_tip(0) <= load_tmp_d_133_d_ack_top;
  place_432_rst(0) <= oper_tmp_d_134_float_d_req_top;
  place_433_tip(0) <= oper_tmp_d_135_float_d_req_top;
  place_433_rst(0) <= oper_tmp_d_135_float_d_ack_top;
  place_434_tip(0) <= load_tmp_d_123_d_ack_top;
  place_434_rst(0) <= oper_tmp_d_135_float_d_req_top;
  place_435_tip(0) <= oper_tmp_d_134_float_d_ack_top;
  place_435_rst(0) <= oper_tmp_d_135_float_d_req_top;
  place_436_tip(0) <= store_5_d_req_top;
  place_436_rst(0) <= store_5_d_ack_top;
  place_437_tip(0) <= oper_tmp_d_118_d_lvl_d_2_uint_d_ack_top;
  place_437_rst(0) <= store_5_d_req_top;
  place_438_tip(0) <= oper_tmp_d_135_float_d_ack_top;
  place_438_rst(0) <= store_5_d_req_top;
  place_439_tip(0) <= load_tmp_d_133_d_ack_top;
  place_439_rst(0) <= store_5_d_req_top;
  place_440_tip(0) <= store_5_d_ack_top;
  place_440_rst(0) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  place_441_tip(0) <= oper_j_d_7_int_d_req_top;
  place_441_rst(0) <= oper_j_d_7_int_d_ack_top;
  place_442_tip(0) <= tc_j_d_7_d_1_d_ack_top;
  place_442_rst(0) <= oper_j_d_7_int_d_req_top;
  place_443_tip(0) <= oper_tmp_d_113_bool_d_req_top;
  place_443_rst(0) <= oper_tmp_d_113_bool_d_ack_top;
  place_444_tip(0) <= oper_j_d_7_int_d_ack_top;
  place_444_rst(0) <= oper_tmp_d_113_bool_d_req_top;
  place_445_tip(0) <= oper_indvar_d_next133_uint_d_req_top;
  place_445_rst(0) <= oper_indvar_d_next133_uint_d_ack_top;
  place_446_tip(0) <= no_exit_d_8_d_entry_top;
  place_446_rst(0) <= oper_indvar_d_next133_uint_d_req_top;
  place_447_tip(0) <= oper_indvar_d_next133_uint_d_ack_top;
  place_447_rst(0) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  place_448_tip(0) <= oper_tmp_d_113_bool_d_ack_top;
  place_448_rst(0) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  place_449_tip(0) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  place_449_rst(0) <= no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_top;
  place_449_rst(1) <= no_exit_d_8_to_no_exit_d_8_src_top;
  place_450_tip(0) <= store_5_d_ack_top;
  place_450_rst(0) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  place_451_tip(0) <= oper_exitcond142_bool_d_req_top;
  place_451_rst(0) <= oper_exitcond142_bool_d_ack_top;
  place_453_tip(0) <= oper_exitcond142_bool_d_ack_top;
  place_453_rst(0) <= cbr_18_oper_exitcond142_bool_d_req_top;
  place_454_tip(0) <= cbr_18_oper_exitcond142_bool_d_req_top;
  place_454_rst(0) <= loopexit_d_7_to_loopentry_d_7_d_outer_src_top;
  place_454_rst(1) <= loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_top;
  place_457_tip(0) <= indvar143_mux_1_d_req0_top;
  place_457_tip(1) <= indvar143_mux_1_d_req1_top;
  place_457_rst(0) <= indvar143_mux_1_d_ack_top;
  place_458_tip(0) <= indvar143_mux_1_d_ack_top;
  place_458_rst(0) <= tc_i_d_3_d_0_d_ph_d_req_top;
  place_459_tip(0) <= loopexit_d_10_to_no_exit_d_10_d_outer_src_top;
  place_459_rst(0) <= indvar143_mux_1_d_req0_top;
  place_46_tip(0) <= no_exit_d_7_to_loopentry_d_7_d_backedge_src_top;
  place_46_tip(1) <= no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_top;
  place_46_rst(0) <= oper_indvar_d_next139_uint_d_req_top;
  place_460_tip(0) <= tc_i_d_3_d_0_d_ph_d_req_top;
  place_460_rst(0) <= tc_i_d_3_d_0_d_ph_d_ack_top;
  place_462_tip(0) <= tc_i_d_3_d_0_d_ph_d_ack_top;
  place_462_rst(0) <= j_d_9_d_2_mux_1_d_req0_top;
  place_464_tip(0) <= j_d_9_d_2_mux_1_d_req0_top;
  place_464_tip(1) <= j_d_9_d_2_mux_1_d_req1_top;
  place_464_rst(0) <= j_d_9_d_2_mux_1_d_ack_top;
  place_465_tip(0) <= j_d_9_d_2_mux_1_d_ack_top;
  place_465_rst(0) <= oper_tmp_d_149_bool_d_req_top;
  place_467_tip(0) <= oper_tmp_d_149_bool_d_req_top;
  place_467_rst(0) <= oper_tmp_d_149_bool_d_ack_top;
  place_469_tip(0) <= oper_tmp_d_149_bool_d_ack_top;
  place_469_rst(0) <= cbr_19_oper_tmp_d_149_bool_d_req_top;
  place_470_tip(0) <= cbr_19_oper_tmp_d_149_bool_d_req_top;
  place_470_rst(0) <= no_exit_d_10_to_else_d_0_src_top;
  place_470_rst(1) <= no_exit_d_10_to_then_d_1_src_top;
  place_471_tip(0) <= oper_tmp_d_154_d_id_d_1_uint_d_req_top;
  place_471_rst(0) <= oper_tmp_d_154_d_id_d_1_uint_d_ack_top;
  place_472_tip(0) <= then_d_1_d_entry_top;
  place_472_rst(0) <= oper_tmp_d_154_d_id_d_1_uint_d_req_top;
  place_473_tip(0) <= oper_tmp_d_154_d_lvl_d_1_uint_d_req_top;
  place_473_rst(0) <= oper_tmp_d_154_d_lvl_d_1_uint_d_ack_top;
  place_474_tip(0) <= oper_tmp_d_154_d_id_d_1_uint_d_ack_top;
  place_474_rst(0) <= oper_tmp_d_154_d_lvl_d_1_uint_d_req_top;
  place_475_tip(0) <= tc_tmp_d_154_d_id_d_2_d_cast_d_req_top;
  place_475_rst(0) <= tc_tmp_d_154_d_id_d_2_d_cast_d_ack_top;
  place_476_tip(0) <= then_d_1_d_entry_top;
  place_476_rst(0) <= tc_tmp_d_154_d_id_d_2_d_cast_d_req_top;
  place_477_tip(0) <= oper_tmp_d_154_d_lvl_d_2_uint_d_req_top;
  place_477_rst(0) <= oper_tmp_d_154_d_lvl_d_2_uint_d_ack_top;
  place_478_tip(0) <= oper_tmp_d_154_d_lvl_d_1_uint_d_ack_top;
  place_478_rst(0) <= oper_tmp_d_154_d_lvl_d_2_uint_d_req_top;
  place_479_tip(0) <= tc_tmp_d_154_d_id_d_2_d_cast_d_ack_top;
  place_479_rst(0) <= oper_tmp_d_154_d_lvl_d_2_uint_d_req_top;
  place_48_tip(0) <= loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_top;
  place_48_rst(0) <= indvar143_mux_1_d_req1_top;
  place_480_tip(0) <= oper_tmp_d_158_d_id_d_1_uint_d_req_top;
  place_480_rst(0) <= oper_tmp_d_158_d_id_d_1_uint_d_ack_top;
  place_481_tip(0) <= then_d_1_d_entry_top;
  place_481_rst(0) <= oper_tmp_d_158_d_id_d_1_uint_d_req_top;
  place_482_tip(0) <= oper_tmp_d_158_d_lvl_d_1_uint_d_req_top;
  place_482_rst(0) <= oper_tmp_d_158_d_lvl_d_1_uint_d_ack_top;
  place_483_tip(0) <= oper_tmp_d_158_d_id_d_1_uint_d_ack_top;
  place_483_rst(0) <= oper_tmp_d_158_d_lvl_d_1_uint_d_req_top;
  place_484_tip(0) <= tc_tmp_d_158_d_id_d_2_d_cast_d_req_top;
  place_484_rst(0) <= tc_tmp_d_158_d_id_d_2_d_cast_d_ack_top;
  place_485_tip(0) <= then_d_1_d_entry_top;
  place_485_rst(0) <= tc_tmp_d_158_d_id_d_2_d_cast_d_req_top;
  place_486_tip(0) <= oper_tmp_d_158_d_lvl_d_2_uint_d_req_top;
  place_486_rst(0) <= oper_tmp_d_158_d_lvl_d_2_uint_d_ack_top;
  place_487_tip(0) <= oper_tmp_d_158_d_lvl_d_1_uint_d_ack_top;
  place_487_rst(0) <= oper_tmp_d_158_d_lvl_d_2_uint_d_req_top;
  place_488_tip(0) <= tc_tmp_d_158_d_id_d_2_d_cast_d_ack_top;
  place_488_rst(0) <= oper_tmp_d_158_d_lvl_d_2_uint_d_req_top;
  place_489_tip(0) <= load_tmp_d_159_d_req_top;
  place_489_rst(0) <= load_tmp_d_159_d_ack_top;
  place_490_tip(0) <= oper_tmp_d_158_d_lvl_d_2_uint_d_ack_top;
  place_490_rst(0) <= load_tmp_d_159_d_req_top;
  place_491_tip(0) <= store_6_d_req_top;
  place_491_rst(0) <= store_6_d_ack_top;
  place_492_tip(0) <= oper_tmp_d_154_d_lvl_d_2_uint_d_ack_top;
  place_492_rst(0) <= store_6_d_req_top;
  place_493_tip(0) <= load_tmp_d_159_d_ack_top;
  place_493_rst(0) <= store_6_d_req_top;
  place_494_tip(0) <= load_tmp_d_159_d_ack_top;
  place_494_rst(0) <= store_6_d_req_top;
  place_495_tip(0) <= store_6_d_ack_top;
  place_495_rst(0) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  place_496_tip(0) <= oper_tmp_d_163_d_id_d_1_uint_d_req_top;
  place_496_rst(0) <= oper_tmp_d_163_d_id_d_1_uint_d_ack_top;
  place_497_tip(0) <= then_d_1_d_entry_top;
  place_497_rst(0) <= oper_tmp_d_163_d_id_d_1_uint_d_req_top;
  place_498_tip(0) <= oper_tmp_d_163_d_lvl_d_1_uint_d_req_top;
  place_498_rst(0) <= oper_tmp_d_163_d_lvl_d_1_uint_d_ack_top;
  place_499_tip(0) <= oper_tmp_d_163_d_id_d_1_uint_d_ack_top;
  place_499_rst(0) <= oper_tmp_d_163_d_lvl_d_1_uint_d_req_top;
  place_5_tip(0) <= no_exit_d_1_to_loopexit_d_1_src_top;
  place_5_rst(0) <= oper_indvar_d_next119_uint_d_req_top;
  place_500_tip(0) <= tc_tmp_d_163_d_id_d_2_d_cast_d_req_top;
  place_500_rst(0) <= tc_tmp_d_163_d_id_d_2_d_cast_d_ack_top;
  place_501_tip(0) <= then_d_1_d_entry_top;
  place_501_rst(0) <= tc_tmp_d_163_d_id_d_2_d_cast_d_req_top;
  place_502_tip(0) <= oper_tmp_d_163_d_lvl_d_2_uint_d_req_top;
  place_502_rst(0) <= oper_tmp_d_163_d_lvl_d_2_uint_d_ack_top;
  place_503_tip(0) <= oper_tmp_d_163_d_lvl_d_1_uint_d_ack_top;
  place_503_rst(0) <= oper_tmp_d_163_d_lvl_d_2_uint_d_req_top;
  place_504_tip(0) <= tc_tmp_d_163_d_id_d_2_d_cast_d_ack_top;
  place_504_rst(0) <= oper_tmp_d_163_d_lvl_d_2_uint_d_req_top;
  place_505_tip(0) <= store_7_d_req_top;
  place_505_rst(0) <= store_7_d_ack_top;
  place_506_tip(0) <= oper_tmp_d_163_d_lvl_d_2_uint_d_ack_top;
  place_506_rst(0) <= store_7_d_req_top;
  place_507_tip(0) <= store_6_d_ack_top;
  place_507_rst(0) <= store_7_d_req_top;
  place_508_tip(0) <= store_7_d_ack_top;
  place_508_rst(0) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  place_509_tip(0) <= oper_inc_d_960_int_d_req_top;
  place_509_rst(0) <= oper_inc_d_960_int_d_ack_top;
  place_510_tip(0) <= then_d_1_d_entry_top;
  place_510_rst(0) <= oper_inc_d_960_int_d_req_top;
  place_511_tip(0) <= oper_tmp_d_14574_bool_d_req_top;
  place_511_rst(0) <= oper_tmp_d_14574_bool_d_ack_top;
  place_512_tip(0) <= oper_inc_d_960_int_d_ack_top;
  place_512_rst(0) <= oper_tmp_d_14574_bool_d_req_top;
  place_513_tip(0) <= oper_tmp_d_14574_bool_d_ack_top;
  place_513_rst(0) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  place_514_tip(0) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  place_514_rst(0) <= then_d_1_to_loopexit_d_10_src_top;
  place_514_rst(1) <= then_d_1_to_no_exit_d_10_d_backedge_src_top;
  place_515_tip(0) <= store_7_d_ack_top;
  place_515_rst(0) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  place_516_tip(0) <= else_d_1_to_no_exit_d_10_d_backedge_src_top;
  place_516_rst(0) <= j_d_9_d_2_d_be_mux_2_d_req1_top;
  place_517_tip(0) <= j_d_9_d_2_d_be_mux_2_d_req0_top;
  place_517_tip(1) <= j_d_9_d_2_d_be_mux_2_d_req1_top;
  place_517_rst(0) <= j_d_9_d_2_d_be_mux_2_d_ack_top;
  place_518_tip(0) <= j_d_9_d_2_d_be_mux_2_d_ack_top;
  place_518_rst(0) <= j_d_9_d_2_mux_1_d_req1_top;
  place_519_tip(0) <= then_d_2_to_no_exit_d_10_d_backedge_src_top;
  place_519_rst(0) <= j_d_9_d_2_d_be_mux_1_d_req1_top;
  place_52_tip(0) <= no_exit_d_10_to_then_d_1_src_top;
  place_52_rst(0) <= then_d_1_d_entry_top;
  place_520_tip(0) <= j_d_9_d_2_d_be_mux_1_d_req0_top;
  place_520_tip(1) <= j_d_9_d_2_d_be_mux_1_d_req1_top;
  place_520_rst(0) <= j_d_9_d_2_d_be_mux_1_d_ack_top;
  place_521_tip(0) <= j_d_9_d_2_d_be_mux_1_d_ack_top;
  place_521_rst(0) <= j_d_9_d_2_d_be_mux_2_d_req0_top;
  place_522_tip(0) <= then_d_1_to_no_exit_d_10_d_backedge_src_top;
  place_522_rst(0) <= j_d_9_d_2_d_be_mux_1_d_req0_top;
  place_524_tip(0) <= oper_tmp_d_166_bool_d_req_top;
  place_524_rst(0) <= oper_tmp_d_166_bool_d_ack_top;
  place_525_tip(0) <= else_d_0_d_entry_top;
  place_525_rst(0) <= oper_tmp_d_166_bool_d_req_top;
  place_526_tip(0) <= oper_tmp_d_171_d_id_d_1_uint_d_req_top;
  place_526_rst(0) <= oper_tmp_d_171_d_id_d_1_uint_d_ack_top;
  place_527_tip(0) <= else_d_0_d_entry_top;
  place_527_rst(0) <= oper_tmp_d_171_d_id_d_1_uint_d_req_top;
  place_528_tip(0) <= oper_tmp_d_171_d_lvl_d_1_uint_d_req_top;
  place_528_rst(0) <= oper_tmp_d_171_d_lvl_d_1_uint_d_ack_top;
  place_529_tip(0) <= oper_tmp_d_171_d_id_d_1_uint_d_ack_top;
  place_529_rst(0) <= oper_tmp_d_171_d_lvl_d_1_uint_d_req_top;
  place_530_tip(0) <= tc_tmp_d_171_d_id_d_2_d_cast_d_req_top;
  place_530_rst(0) <= tc_tmp_d_171_d_id_d_2_d_cast_d_ack_top;
  place_531_tip(0) <= else_d_0_d_entry_top;
  place_531_rst(0) <= tc_tmp_d_171_d_id_d_2_d_cast_d_req_top;
  place_532_tip(0) <= oper_tmp_d_171_d_lvl_d_2_uint_d_req_top;
  place_532_rst(0) <= oper_tmp_d_171_d_lvl_d_2_uint_d_ack_top;
  place_533_tip(0) <= oper_tmp_d_171_d_lvl_d_1_uint_d_ack_top;
  place_533_rst(0) <= oper_tmp_d_171_d_lvl_d_2_uint_d_req_top;
  place_534_tip(0) <= tc_tmp_d_171_d_id_d_2_d_cast_d_ack_top;
  place_534_rst(0) <= oper_tmp_d_171_d_lvl_d_2_uint_d_req_top;
  place_535_tip(0) <= oper_tmp_d_171_d_lvl_d_2_uint_d_ack_top;
  place_535_rst(0) <= cbr_21_oper_tmp_d_166_bool_d_req_top;
  place_536_tip(0) <= oper_tmp_d_166_bool_d_ack_top;
  place_536_rst(0) <= cbr_21_oper_tmp_d_166_bool_d_req_top;
  place_537_tip(0) <= cbr_21_oper_tmp_d_166_bool_d_req_top;
  place_537_rst(0) <= else_d_0_to_else_d_1_src_top;
  place_537_rst(1) <= else_d_0_to_then_d_2_src_top;
  place_538_tip(0) <= store_8_d_req_top;
  place_538_rst(0) <= store_8_d_ack_top;
  place_539_tip(0) <= then_d_2_d_entry_top;
  place_539_rst(0) <= store_8_d_req_top;
  place_54_tip(0) <= no_exit_d_10_to_else_d_0_src_top;
  place_54_rst(0) <= else_d_0_d_entry_top;
  place_540_tip(0) <= store_8_d_ack_top;
  place_540_rst(0) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  place_541_tip(0) <= oper_tmp_d_175_d_id_d_1_uint_d_req_top;
  place_541_rst(0) <= oper_tmp_d_175_d_id_d_1_uint_d_ack_top;
  place_542_tip(0) <= then_d_2_d_entry_top;
  place_542_rst(0) <= oper_tmp_d_175_d_id_d_1_uint_d_req_top;
  place_543_tip(0) <= oper_tmp_d_175_d_lvl_d_1_uint_d_req_top;
  place_543_rst(0) <= oper_tmp_d_175_d_lvl_d_1_uint_d_ack_top;
  place_544_tip(0) <= oper_tmp_d_175_d_id_d_1_uint_d_ack_top;
  place_544_rst(0) <= oper_tmp_d_175_d_lvl_d_1_uint_d_req_top;
  place_545_tip(0) <= tc_tmp_d_175_d_id_d_2_d_cast_d_req_top;
  place_545_rst(0) <= tc_tmp_d_175_d_id_d_2_d_cast_d_ack_top;
  place_546_tip(0) <= then_d_2_d_entry_top;
  place_546_rst(0) <= tc_tmp_d_175_d_id_d_2_d_cast_d_req_top;
  place_547_tip(0) <= oper_tmp_d_175_d_lvl_d_2_uint_d_req_top;
  place_547_rst(0) <= oper_tmp_d_175_d_lvl_d_2_uint_d_ack_top;
  place_548_tip(0) <= oper_tmp_d_175_d_lvl_d_1_uint_d_ack_top;
  place_548_rst(0) <= oper_tmp_d_175_d_lvl_d_2_uint_d_req_top;
  place_549_tip(0) <= tc_tmp_d_175_d_id_d_2_d_cast_d_ack_top;
  place_549_rst(0) <= oper_tmp_d_175_d_lvl_d_2_uint_d_req_top;
  place_550_tip(0) <= oper_tmp_d_179_d_id_d_1_uint_d_req_top;
  place_550_rst(0) <= oper_tmp_d_179_d_id_d_1_uint_d_ack_top;
  place_551_tip(0) <= then_d_2_d_entry_top;
  place_551_rst(0) <= oper_tmp_d_179_d_id_d_1_uint_d_req_top;
  place_552_tip(0) <= oper_tmp_d_179_d_lvl_d_1_uint_d_req_top;
  place_552_rst(0) <= oper_tmp_d_179_d_lvl_d_1_uint_d_ack_top;
  place_553_tip(0) <= oper_tmp_d_179_d_id_d_1_uint_d_ack_top;
  place_553_rst(0) <= oper_tmp_d_179_d_lvl_d_1_uint_d_req_top;
  place_554_tip(0) <= tc_tmp_d_179_d_id_d_2_d_cast_d_req_top;
  place_554_rst(0) <= tc_tmp_d_179_d_id_d_2_d_cast_d_ack_top;
  place_555_tip(0) <= then_d_2_d_entry_top;
  place_555_rst(0) <= tc_tmp_d_179_d_id_d_2_d_cast_d_req_top;
  place_556_tip(0) <= oper_tmp_d_179_d_lvl_d_2_uint_d_req_top;
  place_556_rst(0) <= oper_tmp_d_179_d_lvl_d_2_uint_d_ack_top;
  place_557_tip(0) <= oper_tmp_d_179_d_lvl_d_1_uint_d_ack_top;
  place_557_rst(0) <= oper_tmp_d_179_d_lvl_d_2_uint_d_req_top;
  place_558_tip(0) <= tc_tmp_d_179_d_id_d_2_d_cast_d_ack_top;
  place_558_rst(0) <= oper_tmp_d_179_d_lvl_d_2_uint_d_req_top;
  place_559_tip(0) <= load_tmp_d_180_d_req_top;
  place_559_rst(0) <= load_tmp_d_180_d_ack_top;
  place_560_tip(0) <= oper_tmp_d_179_d_lvl_d_2_uint_d_ack_top;
  place_560_rst(0) <= load_tmp_d_180_d_req_top;
  place_561_tip(0) <= store_8_d_ack_top;
  place_561_rst(0) <= load_tmp_d_180_d_req_top;
  place_562_tip(0) <= store_9_d_req_top;
  place_562_rst(0) <= store_9_d_ack_top;
  place_563_tip(0) <= oper_tmp_d_175_d_lvl_d_2_uint_d_ack_top;
  place_563_rst(0) <= store_9_d_req_top;
  place_564_tip(0) <= load_tmp_d_180_d_ack_top;
  place_564_rst(0) <= store_9_d_req_top;
  place_565_tip(0) <= load_tmp_d_180_d_ack_top;
  place_565_rst(0) <= store_9_d_req_top;
  place_566_tip(0) <= store_9_d_ack_top;
  place_566_rst(0) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  place_567_tip(0) <= oper_inc_d_976_int_d_req_top;
  place_567_rst(0) <= oper_inc_d_976_int_d_ack_top;
  place_568_tip(0) <= then_d_2_d_entry_top;
  place_568_rst(0) <= oper_inc_d_976_int_d_req_top;
  place_569_tip(0) <= oper_tmp_d_14578_bool_d_req_top;
  place_569_rst(0) <= oper_tmp_d_14578_bool_d_ack_top;
  place_570_tip(0) <= oper_inc_d_976_int_d_ack_top;
  place_570_rst(0) <= oper_tmp_d_14578_bool_d_req_top;
  place_571_tip(0) <= oper_tmp_d_14578_bool_d_ack_top;
  place_571_rst(0) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  place_572_tip(0) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  place_572_rst(0) <= then_d_2_to_loopexit_d_10_src_top;
  place_572_rst(1) <= then_d_2_to_no_exit_d_10_d_backedge_src_top;
  place_573_tip(0) <= store_9_d_ack_top;
  place_573_rst(0) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  place_574_tip(0) <= store_10_d_req_top;
  place_574_rst(0) <= store_10_d_ack_top;
  place_575_tip(0) <= else_d_1_d_entry_top;
  place_575_rst(0) <= store_10_d_req_top;
  place_576_tip(0) <= store_10_d_ack_top;
  place_576_rst(0) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  place_577_tip(0) <= oper_tmp_d_188_d_id_d_1_uint_d_req_top;
  place_577_rst(0) <= oper_tmp_d_188_d_id_d_1_uint_d_ack_top;
  place_578_tip(0) <= else_d_1_d_entry_top;
  place_578_rst(0) <= oper_tmp_d_188_d_id_d_1_uint_d_req_top;
  place_579_tip(0) <= oper_tmp_d_188_d_lvl_d_1_uint_d_req_top;
  place_579_rst(0) <= oper_tmp_d_188_d_lvl_d_1_uint_d_ack_top;
  place_580_tip(0) <= oper_tmp_d_188_d_id_d_1_uint_d_ack_top;
  place_580_rst(0) <= oper_tmp_d_188_d_lvl_d_1_uint_d_req_top;
  place_581_tip(0) <= tc_tmp_d_188_d_id_d_2_d_cast_d_req_top;
  place_581_rst(0) <= tc_tmp_d_188_d_id_d_2_d_cast_d_ack_top;
  place_582_tip(0) <= else_d_1_d_entry_top;
  place_582_rst(0) <= tc_tmp_d_188_d_id_d_2_d_cast_d_req_top;
  place_583_tip(0) <= oper_tmp_d_188_d_lvl_d_2_uint_d_req_top;
  place_583_rst(0) <= oper_tmp_d_188_d_lvl_d_2_uint_d_ack_top;
  place_584_tip(0) <= oper_tmp_d_188_d_lvl_d_1_uint_d_ack_top;
  place_584_rst(0) <= oper_tmp_d_188_d_lvl_d_2_uint_d_req_top;
  place_585_tip(0) <= tc_tmp_d_188_d_id_d_2_d_cast_d_ack_top;
  place_585_rst(0) <= oper_tmp_d_188_d_lvl_d_2_uint_d_req_top;
  place_586_tip(0) <= oper_tmp_d_192_d_id_d_1_uint_d_req_top;
  place_586_rst(0) <= oper_tmp_d_192_d_id_d_1_uint_d_ack_top;
  place_587_tip(0) <= else_d_1_d_entry_top;
  place_587_rst(0) <= oper_tmp_d_192_d_id_d_1_uint_d_req_top;
  place_588_tip(0) <= oper_tmp_d_192_d_lvl_d_1_uint_d_req_top;
  place_588_rst(0) <= oper_tmp_d_192_d_lvl_d_1_uint_d_ack_top;
  place_589_tip(0) <= oper_tmp_d_192_d_id_d_1_uint_d_ack_top;
  place_589_rst(0) <= oper_tmp_d_192_d_lvl_d_1_uint_d_req_top;
  place_59_tip(0) <= else_d_0_to_then_d_2_src_top;
  place_59_rst(0) <= then_d_2_d_entry_top;
  place_590_tip(0) <= tc_tmp_d_192_d_id_d_2_d_cast_d_req_top;
  place_590_rst(0) <= tc_tmp_d_192_d_id_d_2_d_cast_d_ack_top;
  place_591_tip(0) <= else_d_1_d_entry_top;
  place_591_rst(0) <= tc_tmp_d_192_d_id_d_2_d_cast_d_req_top;
  place_592_tip(0) <= oper_tmp_d_192_d_lvl_d_2_uint_d_req_top;
  place_592_rst(0) <= oper_tmp_d_192_d_lvl_d_2_uint_d_ack_top;
  place_593_tip(0) <= oper_tmp_d_192_d_lvl_d_1_uint_d_ack_top;
  place_593_rst(0) <= oper_tmp_d_192_d_lvl_d_2_uint_d_req_top;
  place_594_tip(0) <= tc_tmp_d_192_d_id_d_2_d_cast_d_ack_top;
  place_594_rst(0) <= oper_tmp_d_192_d_lvl_d_2_uint_d_req_top;
  place_595_tip(0) <= load_tmp_d_193_d_req_top;
  place_595_rst(0) <= load_tmp_d_193_d_ack_top;
  place_596_tip(0) <= oper_tmp_d_192_d_lvl_d_2_uint_d_ack_top;
  place_596_rst(0) <= load_tmp_d_193_d_req_top;
  place_597_tip(0) <= store_10_d_ack_top;
  place_597_rst(0) <= load_tmp_d_193_d_req_top;
  place_598_tip(0) <= store_11_d_req_top;
  place_598_rst(0) <= store_11_d_ack_top;
  place_599_tip(0) <= oper_tmp_d_188_d_lvl_d_2_uint_d_ack_top;
  place_599_rst(0) <= store_11_d_req_top;
  place_600_tip(0) <= load_tmp_d_193_d_ack_top;
  place_600_rst(0) <= store_11_d_req_top;
  place_601_tip(0) <= load_tmp_d_193_d_ack_top;
  place_601_rst(0) <= store_11_d_req_top;
  place_602_tip(0) <= store_11_d_ack_top;
  place_602_rst(0) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  place_603_tip(0) <= oper_inc_d_9_int_d_req_top;
  place_603_rst(0) <= oper_inc_d_9_int_d_ack_top;
  place_604_tip(0) <= else_d_1_d_entry_top;
  place_604_rst(0) <= oper_inc_d_9_int_d_req_top;
  place_605_tip(0) <= oper_tmp_d_14580_bool_d_req_top;
  place_605_rst(0) <= oper_tmp_d_14580_bool_d_ack_top;
  place_606_tip(0) <= oper_inc_d_9_int_d_ack_top;
  place_606_rst(0) <= oper_tmp_d_14580_bool_d_req_top;
  place_607_tip(0) <= oper_tmp_d_14580_bool_d_ack_top;
  place_607_rst(0) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  place_608_tip(0) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  place_608_rst(0) <= else_d_1_to_loopexit_d_10_src_top;
  place_608_rst(1) <= else_d_1_to_no_exit_d_10_d_backedge_src_top;
  place_609_tip(0) <= store_11_d_ack_top;
  place_609_rst(0) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  place_61_tip(0) <= else_d_0_to_else_d_1_src_top;
  place_61_rst(0) <= else_d_1_d_entry_top;
  place_610_tip(0) <= oper_indvar_d_next144_uint_d_req_top;
  place_610_rst(0) <= oper_indvar_d_next144_uint_d_ack_top;
  place_612_tip(0) <= oper_exitcond145_bool_d_req_top;
  place_612_rst(0) <= oper_exitcond145_bool_d_ack_top;
  place_613_tip(0) <= oper_indvar_d_next144_uint_d_ack_top;
  place_613_rst(0) <= oper_exitcond145_bool_d_req_top;
  place_614_tip(0) <= oper_exitcond145_bool_d_ack_top;
  place_614_rst(0) <= cbr_24_oper_exitcond145_bool_d_req_top;
  place_615_tip(0) <= cbr_24_oper_exitcond145_bool_d_req_top;
  place_615_rst(0) <= loopexit_d_10_to_loopentry_d_12_d_loopexit_src_top;
  place_615_rst(1) <= loopexit_d_10_to_no_exit_d_10_d_outer_src_top;
  place_617_tip(0) <= loopentry_d_12_d_loopexit_to_loopentry_d_12_src_top;
  place_617_rst(0) <= indvar148_mux_1_d_req1_top;
  place_618_tip(0) <= indvar148_mux_1_d_req0_top;
  place_618_tip(1) <= indvar148_mux_1_d_req1_top;
  place_618_rst(0) <= indvar148_mux_1_d_ack_top;
  place_619_tip(0) <= indvar148_mux_1_d_ack_top;
  place_619_rst(0) <= loopentry_d_12_d_pre_top;
  place_620_tip(0) <= loopexit_d_12_to_loopentry_d_12_src_top;
  place_620_rst(0) <= indvar148_mux_1_d_req0_top;
  place_621_tip(0) <= loopentry_d_12_d_loopexit_to_loopentry_d_12_src_top;
  place_621_rst(0) <= k_d_3_d_0_mux_1_d_req1_top;
  place_622_tip(0) <= k_d_3_d_0_mux_1_d_req0_top;
  place_622_tip(1) <= k_d_3_d_0_mux_1_d_req1_top;
  place_622_rst(0) <= k_d_3_d_0_mux_1_d_ack_top;
  place_623_tip(0) <= k_d_3_d_0_mux_1_d_ack_top;
  place_623_rst(0) <= loopentry_d_12_d_pre_top;
  place_624_tip(0) <= loopexit_d_12_to_loopentry_d_12_src_top;
  place_624_rst(0) <= k_d_3_d_0_mux_1_d_req0_top;
  place_625_tip(0) <= loopentry_d_12_d_entry_top;
  place_625_rst(0) <= cbr_25_oper_tmp_d_202_bool_d_req_top;
  place_626_tip(0) <= tc_i_d_4_d_0_d_req_top;
  place_626_rst(0) <= tc_i_d_4_d_0_d_ack_top;
  place_627_tip(0) <= loopentry_d_12_d_entry_top;
  place_627_rst(0) <= tc_i_d_4_d_0_d_req_top;
  place_628_tip(0) <= tc_i_d_4_d_0_d_ack_top;
  place_628_rst(0) <= cbr_25_oper_tmp_d_202_bool_d_req_top;
  place_629_tip(0) <= oper_tmp_d_202_bool_d_req_top;
  place_629_rst(0) <= oper_tmp_d_202_bool_d_ack_top;
  place_63_tip(0) <= else_d_1_to_loopexit_d_10_src_top;
  place_63_tip(1) <= then_d_1_to_loopexit_d_10_src_top;
  place_63_tip(2) <= then_d_2_to_loopexit_d_10_src_top;
  place_63_rst(0) <= oper_indvar_d_next144_uint_d_req_top;
  place_630_tip(0) <= loopentry_d_12_d_entry_top;
  place_630_rst(0) <= oper_tmp_d_202_bool_d_req_top;
  place_631_tip(0) <= oper_tmp_d_202_bool_d_ack_top;
  place_631_rst(0) <= cbr_25_oper_tmp_d_202_bool_d_req_top;
  place_632_tip(0) <= cbr_25_oper_tmp_d_202_bool_d_req_top;
  place_632_rst(0) <= loopentry_d_12_to_loopexit_d_12_src_top;
  place_632_rst(1) <= loopentry_d_12_to_no_exit_d_12_d_preheader_src_top;
  place_635_tip(0) <= indvar146_mux_1_d_req0_top;
  place_635_tip(1) <= indvar146_mux_1_d_req1_top;
  place_635_rst(0) <= indvar146_mux_1_d_ack_top;
  place_636_tip(0) <= indvar146_mux_1_d_ack_top;
  place_636_rst(0) <= no_exit_d_12_d_entry_top;
  place_637_tip(0) <= no_exit_d_12_to_no_exit_d_12_src_top;
  place_637_rst(0) <= indvar146_mux_1_d_req0_top;
  place_638_tip(0) <= tc_j_d_11_d_2_d_req_top;
  place_638_rst(0) <= tc_j_d_11_d_2_d_ack_top;
  place_639_tip(0) <= no_exit_d_12_d_entry_top;
  place_639_rst(0) <= tc_j_d_11_d_2_d_req_top;
  place_640_tip(0) <= oper_k_d_2_d_2_int_d_req_top;
  place_640_rst(0) <= oper_k_d_2_d_2_int_d_ack_top;
  place_641_tip(0) <= tc_j_d_11_d_2_d_ack_top;
  place_641_rst(0) <= oper_k_d_2_d_2_int_d_req_top;
  place_642_tip(0) <= tc_tmp_d_206_d_id_d_0_d_cast_d_req_top;
  place_642_rst(0) <= tc_tmp_d_206_d_id_d_0_d_cast_d_ack_top;
  place_643_tip(0) <= oper_k_d_2_d_2_int_d_ack_top;
  place_643_rst(0) <= tc_tmp_d_206_d_id_d_0_d_cast_d_req_top;
  place_644_tip(0) <= oper_tmp_d_206_d_lvl_d_0_uint_d_req_top;
  place_644_rst(0) <= oper_tmp_d_206_d_lvl_d_0_uint_d_ack_top;
  place_645_tip(0) <= tc_tmp_d_206_d_id_d_0_d_cast_d_ack_top;
  place_645_rst(0) <= oper_tmp_d_206_d_lvl_d_0_uint_d_req_top;
  place_646_tip(0) <= oper_tmp_d_210_d_id_d_1_uint_d_req_top;
  place_646_rst(0) <= oper_tmp_d_210_d_id_d_1_uint_d_ack_top;
  place_647_tip(0) <= no_exit_d_12_d_entry_top;
  place_647_rst(0) <= oper_tmp_d_210_d_id_d_1_uint_d_req_top;
  place_648_tip(0) <= oper_tmp_d_210_d_lvl_d_1_uint_d_req_top;
  place_648_rst(0) <= oper_tmp_d_210_d_lvl_d_1_uint_d_ack_top;
  place_649_tip(0) <= oper_tmp_d_210_d_id_d_1_uint_d_ack_top;
  place_649_rst(0) <= oper_tmp_d_210_d_lvl_d_1_uint_d_req_top;
  place_65_tip(0) <= loopexit_d_10_to_loopentry_d_12_d_loopexit_src_top;
  place_65_rst(0) <= loopentry_d_12_d_loopexit_to_loopentry_d_12_src_top;
  place_650_tip(0) <= oper_tmp_d_210_d_lvl_d_2_uint_d_req_top;
  place_650_rst(0) <= oper_tmp_d_210_d_lvl_d_2_uint_d_ack_top;
  place_651_tip(0) <= oper_tmp_d_210_d_lvl_d_1_uint_d_ack_top;
  place_651_rst(0) <= oper_tmp_d_210_d_lvl_d_2_uint_d_req_top;
  place_652_tip(0) <= load_tmp_d_211_d_req_top;
  place_652_rst(0) <= load_tmp_d_211_d_ack_top;
  place_653_tip(0) <= oper_tmp_d_210_d_lvl_d_2_uint_d_ack_top;
  place_653_rst(0) <= load_tmp_d_211_d_req_top;
  place_654_tip(0) <= store_12_d_req_top;
  place_654_rst(0) <= store_12_d_ack_top;
  place_655_tip(0) <= oper_tmp_d_206_d_lvl_d_0_uint_d_ack_top;
  place_655_rst(0) <= store_12_d_req_top;
  place_656_tip(0) <= load_tmp_d_211_d_ack_top;
  place_656_rst(0) <= store_12_d_req_top;
  place_657_tip(0) <= load_tmp_d_211_d_ack_top;
  place_657_rst(0) <= store_12_d_req_top;
  place_658_tip(0) <= store_12_d_ack_top;
  place_658_rst(0) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  place_659_tip(0) <= oper_inc_d_12_int_d_req_top;
  place_659_rst(0) <= oper_inc_d_12_int_d_ack_top;
  place_66_tip(0) <= loopentry_d_12_d_pre_top;
  place_66_rst(0) <= loopentry_d_12_d_entry_top;
  place_660_tip(0) <= tc_j_d_11_d_2_d_ack_top;
  place_660_rst(0) <= oper_inc_d_12_int_d_req_top;
  place_661_tip(0) <= oper_tmp_d_20299_bool_d_req_top;
  place_661_rst(0) <= oper_tmp_d_20299_bool_d_ack_top;
  place_662_tip(0) <= oper_inc_d_12_int_d_ack_top;
  place_662_rst(0) <= oper_tmp_d_20299_bool_d_req_top;
  place_663_tip(0) <= oper_indvar_d_next147_uint_d_req_top;
  place_663_rst(0) <= oper_indvar_d_next147_uint_d_ack_top;
  place_664_tip(0) <= no_exit_d_12_d_entry_top;
  place_664_rst(0) <= oper_indvar_d_next147_uint_d_req_top;
  place_665_tip(0) <= oper_indvar_d_next147_uint_d_ack_top;
  place_665_rst(0) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  place_666_tip(0) <= oper_tmp_d_20299_bool_d_ack_top;
  place_666_rst(0) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  place_667_tip(0) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  place_667_rst(0) <= no_exit_d_12_to_loopexit_d_12_d_loopexit_src_top;
  place_667_rst(1) <= no_exit_d_12_to_no_exit_d_12_src_top;
  place_668_tip(0) <= store_12_d_ack_top;
  place_668_rst(0) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  place_669_tip(0) <= oper_inc_d_11_int_d_req_top;
  place_669_rst(0) <= oper_inc_d_11_int_d_ack_top;
  place_671_tip(0) <= oper_inc_d_11_int_d_ack_top;
  place_671_rst(0) <= k_d_2_d_3_mux_1_d_req1_top;
  place_673_tip(0) <= k_d_2_d_3_mux_1_d_req0_top;
  place_673_tip(1) <= k_d_2_d_3_mux_1_d_req1_top;
  place_673_rst(0) <= k_d_2_d_3_mux_1_d_ack_top;
  place_674_tip(0) <= k_d_2_d_3_mux_1_d_ack_top;
  place_674_rst(0) <= loopexit_d_12_d_entry_top;
  place_675_tip(0) <= loopentry_d_12_to_loopexit_d_12_src_top;
  place_675_rst(0) <= k_d_2_d_3_mux_1_d_req0_top;
  place_676_tip(0) <= loopexit_d_12_d_entry_top;
  place_676_rst(0) <= cbr_27_oper_exitcond150_bool_d_req_top;
  place_677_tip(0) <= oper_indvar_d_next149_uint_d_req_top;
  place_677_rst(0) <= oper_indvar_d_next149_uint_d_ack_top;
  place_678_tip(0) <= loopexit_d_12_d_entry_top;
  place_678_rst(0) <= oper_indvar_d_next149_uint_d_req_top;
  place_679_tip(0) <= oper_exitcond150_bool_d_req_top;
  place_679_rst(0) <= oper_exitcond150_bool_d_ack_top;
  place_680_tip(0) <= oper_indvar_d_next149_uint_d_ack_top;
  place_680_rst(0) <= oper_exitcond150_bool_d_req_top;
  place_681_tip(0) <= oper_exitcond150_bool_d_ack_top;
  place_681_rst(0) <= cbr_27_oper_exitcond150_bool_d_req_top;
  place_682_tip(0) <= cbr_27_oper_exitcond150_bool_d_req_top;
  place_682_rst(0) <= loopexit_d_12_to_loopentry_d_12_src_top;
  place_682_rst(1) <= loopexit_d_12_to_loopentry_d_14_d_loopexit_src_top;
  place_684_tip(0) <= loopentry_d_14_d_loopexit_to_loopentry_d_14_src_top;
  place_684_rst(0) <= indvar153_mux_1_d_req1_top;
  place_685_tip(0) <= indvar153_mux_1_d_req0_top;
  place_685_tip(1) <= indvar153_mux_1_d_req1_top;
  place_685_rst(0) <= indvar153_mux_1_d_ack_top;
  place_686_tip(0) <= indvar153_mux_1_d_ack_top;
  place_686_rst(0) <= loopentry_d_14_d_pre_top;
  place_687_tip(0) <= loopexit_d_14_to_loopentry_d_14_src_top;
  place_687_rst(0) <= indvar153_mux_1_d_req0_top;
  place_688_tip(0) <= loopentry_d_14_d_loopexit_to_loopentry_d_14_src_top;
  place_688_rst(0) <= k_d_5_d_0_mux_1_d_req1_top;
  place_689_tip(0) <= k_d_5_d_0_mux_1_d_req0_top;
  place_689_tip(1) <= k_d_5_d_0_mux_1_d_req1_top;
  place_689_rst(0) <= k_d_5_d_0_mux_1_d_ack_top;
  place_69_tip(0) <= loopentry_d_12_to_no_exit_d_12_d_preheader_src_top;
  place_69_rst(0) <= indvar146_mux_1_d_req1_top;
  place_690_tip(0) <= k_d_5_d_0_mux_1_d_ack_top;
  place_690_rst(0) <= loopentry_d_14_d_pre_top;
  place_691_tip(0) <= loopexit_d_14_to_loopentry_d_14_src_top;
  place_691_rst(0) <= k_d_5_d_0_mux_1_d_req0_top;
  place_692_tip(0) <= loopentry_d_14_d_entry_top;
  place_692_rst(0) <= cbr_28_oper_tmp_d_221_bool_d_req_top;
  place_693_tip(0) <= tc_i_d_5_d_0_d_req_top;
  place_693_rst(0) <= tc_i_d_5_d_0_d_ack_top;
  place_694_tip(0) <= loopentry_d_14_d_entry_top;
  place_694_rst(0) <= tc_i_d_5_d_0_d_req_top;
  place_695_tip(0) <= oper_tmp_d_221_bool_d_req_top;
  place_695_rst(0) <= oper_tmp_d_221_bool_d_ack_top;
  place_696_tip(0) <= tc_i_d_5_d_0_d_ack_top;
  place_696_rst(0) <= oper_tmp_d_221_bool_d_req_top;
  place_697_tip(0) <= oper_tmp_d_221_bool_d_ack_top;
  place_697_rst(0) <= cbr_28_oper_tmp_d_221_bool_d_req_top;
  place_698_tip(0) <= cbr_28_oper_tmp_d_221_bool_d_req_top;
  place_698_rst(0) <= loopentry_d_14_to_loopexit_d_14_src_top;
  place_698_rst(1) <= loopentry_d_14_to_no_exit_d_14_d_preheader_src_top;
  place_7_tip(0) <= loopexit_d_1_to_loopentry_d_2_src_top;
  place_7_rst(0) <= oper_tmp_d_16_bool_d_req_top;
  place_701_tip(0) <= indvar151_mux_1_d_req0_top;
  place_701_tip(1) <= indvar151_mux_1_d_req1_top;
  place_701_rst(0) <= indvar151_mux_1_d_ack_top;
  place_702_tip(0) <= indvar151_mux_1_d_ack_top;
  place_702_rst(0) <= no_exit_d_14_d_entry_top;
  place_703_tip(0) <= no_exit_d_14_to_no_exit_d_14_src_top;
  place_703_rst(0) <= indvar151_mux_1_d_req0_top;
  place_704_tip(0) <= tc_indvar151_d_req_top;
  place_704_rst(0) <= tc_indvar151_d_ack_top;
  place_705_tip(0) <= no_exit_d_14_d_entry_top;
  place_705_rst(0) <= tc_indvar151_d_req_top;
  place_706_tip(0) <= oper_tmp_d_155_uint_d_req_top;
  place_706_rst(0) <= oper_tmp_d_155_uint_d_ack_top;
  place_707_tip(0) <= no_exit_d_14_d_entry_top;
  place_707_rst(0) <= oper_tmp_d_155_uint_d_req_top;
  place_708_tip(0) <= tc_j_d_13_d_2_d_req_top;
  place_708_rst(0) <= tc_j_d_13_d_2_d_ack_top;
  place_709_tip(0) <= oper_tmp_d_155_uint_d_ack_top;
  place_709_rst(0) <= tc_j_d_13_d_2_d_req_top;
  place_710_tip(0) <= oper_k_d_4_d_2_int_d_req_top;
  place_710_rst(0) <= oper_k_d_4_d_2_int_d_ack_top;
  place_711_tip(0) <= tc_indvar151_d_ack_top;
  place_711_rst(0) <= oper_k_d_4_d_2_int_d_req_top;
  place_712_tip(0) <= tc_tmp_d_225_d_id_d_0_d_cast_d_req_top;
  place_712_rst(0) <= tc_tmp_d_225_d_id_d_0_d_cast_d_ack_top;
  place_713_tip(0) <= oper_k_d_4_d_2_int_d_ack_top;
  place_713_rst(0) <= tc_tmp_d_225_d_id_d_0_d_cast_d_req_top;
  place_714_tip(0) <= oper_tmp_d_225_d_lvl_d_0_uint_d_req_top;
  place_714_rst(0) <= oper_tmp_d_225_d_lvl_d_0_uint_d_ack_top;
  place_715_tip(0) <= tc_tmp_d_225_d_id_d_0_d_cast_d_ack_top;
  place_715_rst(0) <= oper_tmp_d_225_d_lvl_d_0_uint_d_req_top;
  place_716_tip(0) <= oper_tmp_d_229_d_id_d_1_uint_d_req_top;
  place_716_rst(0) <= oper_tmp_d_229_d_id_d_1_uint_d_ack_top;
  place_717_tip(0) <= no_exit_d_14_d_entry_top;
  place_717_rst(0) <= oper_tmp_d_229_d_id_d_1_uint_d_req_top;
  place_718_tip(0) <= oper_tmp_d_229_d_lvl_d_1_uint_d_req_top;
  place_718_rst(0) <= oper_tmp_d_229_d_lvl_d_1_uint_d_ack_top;
  place_719_tip(0) <= oper_tmp_d_229_d_id_d_1_uint_d_ack_top;
  place_719_rst(0) <= oper_tmp_d_229_d_lvl_d_1_uint_d_req_top;
  place_72_tip(0) <= no_exit_d_12_to_loopexit_d_12_d_loopexit_src_top;
  place_72_rst(0) <= oper_inc_d_11_int_d_req_top;
  place_720_tip(0) <= oper_tmp_d_229_d_lvl_d_2_uint_d_req_top;
  place_720_rst(0) <= oper_tmp_d_229_d_lvl_d_2_uint_d_ack_top;
  place_721_tip(0) <= oper_tmp_d_229_d_lvl_d_1_uint_d_ack_top;
  place_721_rst(0) <= oper_tmp_d_229_d_lvl_d_2_uint_d_req_top;
  place_722_tip(0) <= oper_tmp_d_155_uint_d_ack_top;
  place_722_rst(0) <= oper_tmp_d_229_d_lvl_d_2_uint_d_req_top;
  place_723_tip(0) <= load_tmp_d_230_d_req_top;
  place_723_rst(0) <= load_tmp_d_230_d_ack_top;
  place_724_tip(0) <= oper_tmp_d_229_d_lvl_d_2_uint_d_ack_top;
  place_724_rst(0) <= load_tmp_d_230_d_req_top;
  place_725_tip(0) <= store_13_d_req_top;
  place_725_rst(0) <= store_13_d_ack_top;
  place_726_tip(0) <= oper_tmp_d_225_d_lvl_d_0_uint_d_ack_top;
  place_726_rst(0) <= store_13_d_req_top;
  place_727_tip(0) <= load_tmp_d_230_d_ack_top;
  place_727_rst(0) <= store_13_d_req_top;
  place_728_tip(0) <= load_tmp_d_230_d_ack_top;
  place_728_rst(0) <= store_13_d_req_top;
  place_729_tip(0) <= store_13_d_ack_top;
  place_729_rst(0) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  place_730_tip(0) <= oper_inc_d_15_int_d_req_top;
  place_730_rst(0) <= oper_inc_d_15_int_d_ack_top;
  place_731_tip(0) <= tc_j_d_13_d_2_d_ack_top;
  place_731_rst(0) <= oper_inc_d_15_int_d_req_top;
  place_732_tip(0) <= oper_tmp_d_221111_bool_d_req_top;
  place_732_rst(0) <= oper_tmp_d_221111_bool_d_ack_top;
  place_733_tip(0) <= oper_inc_d_15_int_d_ack_top;
  place_733_rst(0) <= oper_tmp_d_221111_bool_d_req_top;
  place_734_tip(0) <= oper_indvar_d_next152_uint_d_req_top;
  place_734_rst(0) <= oper_indvar_d_next152_uint_d_ack_top;
  place_735_tip(0) <= no_exit_d_14_d_entry_top;
  place_735_rst(0) <= oper_indvar_d_next152_uint_d_req_top;
  place_736_tip(0) <= oper_indvar_d_next152_uint_d_ack_top;
  place_736_rst(0) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  place_737_tip(0) <= oper_tmp_d_221111_bool_d_ack_top;
  place_737_rst(0) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  place_738_tip(0) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  place_738_rst(0) <= no_exit_d_14_to_loopexit_d_14_d_loopexit_src_top;
  place_738_rst(1) <= no_exit_d_14_to_no_exit_d_14_src_top;
  place_739_tip(0) <= store_13_d_ack_top;
  place_739_rst(0) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  place_74_tip(0) <= loopexit_d_12_to_loopentry_d_14_d_loopexit_src_top;
  place_74_rst(0) <= loopentry_d_14_d_loopexit_to_loopentry_d_14_src_top;
  place_740_tip(0) <= oper_inc_d_14_int_d_req_top;
  place_740_rst(0) <= oper_inc_d_14_int_d_ack_top;
  place_742_tip(0) <= oper_inc_d_14_int_d_ack_top;
  place_742_rst(0) <= k_d_4_d_3_mux_1_d_req1_top;
  place_744_tip(0) <= k_d_4_d_3_mux_1_d_req0_top;
  place_744_tip(1) <= k_d_4_d_3_mux_1_d_req1_top;
  place_744_rst(0) <= k_d_4_d_3_mux_1_d_ack_top;
  place_745_tip(0) <= k_d_4_d_3_mux_1_d_ack_top;
  place_745_rst(0) <= loopexit_d_14_d_entry_top;
  place_746_tip(0) <= loopentry_d_14_to_loopexit_d_14_src_top;
  place_746_rst(0) <= k_d_4_d_3_mux_1_d_req0_top;
  place_747_tip(0) <= loopexit_d_14_d_entry_top;
  place_747_rst(0) <= cbr_30_oper_exitcond158_bool_d_req_top;
  place_748_tip(0) <= oper_indvar_d_next157_uint_d_req_top;
  place_748_rst(0) <= oper_indvar_d_next157_uint_d_ack_top;
  place_749_tip(0) <= loopexit_d_14_d_entry_top;
  place_749_rst(0) <= oper_indvar_d_next157_uint_d_req_top;
  place_75_tip(0) <= loopentry_d_14_d_pre_top;
  place_75_rst(0) <= loopentry_d_14_d_entry_top;
  place_750_tip(0) <= oper_exitcond158_bool_d_req_top;
  place_750_rst(0) <= oper_exitcond158_bool_d_ack_top;
  place_751_tip(0) <= oper_indvar_d_next157_uint_d_ack_top;
  place_751_rst(0) <= oper_exitcond158_bool_d_req_top;
  place_752_tip(0) <= oper_exitcond158_bool_d_ack_top;
  place_752_rst(0) <= cbr_30_oper_exitcond158_bool_d_req_top;
  place_753_tip(0) <= cbr_30_oper_exitcond158_bool_d_req_top;
  place_753_rst(0) <= loopexit_d_14_to_loopentry_d_14_src_top;
  place_753_rst(1) <= loopexit_d_14_to_return_src_top;
  place_77_tip(0) <= loopentry_d_14_to_no_exit_d_14_d_preheader_src_top;
  place_77_rst(0) <= indvar151_mux_1_d_req1_top;
  place_81_tip(0) <= no_exit_d_14_to_loopexit_d_14_d_loopexit_src_top;
  place_81_rst(0) <= oper_inc_d_14_int_d_req_top;
  place_83_tip(0) <= loopexit_d_14_to_return_src_top;
  place_83_rst(0) <= fin_top;
  place_84_tip(0) <= fin_top;
  place_84_rst(0) <= init_top;
  place_86_tip(0) <= init_top;
  place_86_rst(0) <= load_noofelem_d_req_top;
  place_87_tip(0) <= load_noofelem_d_req_top;
  place_87_rst(0) <= load_noofelem_d_ack_top;
  place_88_tip(0) <= load_noofelem_d_ack_top;
  place_88_rst(0) <= load_A_d_req_top;
  place_89_tip(0) <= load_A_d_req_top;
  place_89_rst(0) <= load_A_d_ack_top;
  place_9_tip(0) <= loopentry_d_2_to_no_exit_d_2_d_preheader_src_top;
  place_9_rst(0) <= indvar121_mux_1_d_req1_top;
  place_90_tip(0) <= load_A_d_ack_top;
  place_90_rst(0) <= load_rcoeff_d_req_top;
  place_91_tip(0) <= load_rcoeff_d_req_top;
  place_91_rst(0) <= load_rcoeff_d_ack_top;
  place_92_tip(0) <= load_rcoeff_d_ack_top;
  place_92_rst(0) <= load_ccoeff_d_req_top;
  place_93_tip(0) <= load_ccoeff_d_req_top;
  place_93_rst(0) <= load_ccoeff_d_ack_top;
  place_94_tip(0) <= load_ccoeff_d_ack_top;
  place_94_rst(0) <= load_l_array_d_req_top;
  place_95_tip(0) <= load_l_array_d_req_top;
  place_95_rst(0) <= load_l_array_d_ack_top;
  place_96_tip(0) <= load_l_array_d_ack_top;
  place_96_rst(0) <= load_u_array_d_req_top;
  place_97_tip(0) <= load_u_array_d_req_top;
  place_97_rst(0) <= load_u_array_d_ack_top;
  place_99_tip(0) <= loopexit_d_1_to_no_exit_d_1_d_outer_src_top;
  place_99_rst(0) <= indvar118_d_ph_d_ph_mux_1_d_req1_top;

  cbr_10_oper_tmp_d_42_bool_d_req_tip(0) <= place_216_top;
  cbr_10_oper_tmp_d_42_bool_d_req_tip(1) <= place_221_top;
  cbr_11_oper_tmp_d_54_bool_d_req_tip(0) <= place_239_top;
  cbr_11_oper_tmp_d_54_bool_d_req_tip(1) <= place_244_top;
  cbr_11_oper_tmp_d_54_bool_d_req_tip(2) <= place_255_top;
  cbr_12_oper_tmp_d_4223_bool_d_req_tip(0) <= place_263_top;
  cbr_12_oper_tmp_d_4223_bool_d_req_tip(1) <= place_264_top;
  cbr_13_oper_exitcond128_bool_d_req_tip(0) <= place_299_top;
  cbr_13_oper_exitcond128_bool_d_req_tip(1) <= place_304_top;
  cbr_13_oper_exitcond128_bool_d_req_tip(2) <= place_309_top;
  cbr_13_oper_exitcond128_bool_d_req_tip(3) <= place_311_top;
  cbr_14_oper_exitcond131_bool_d_req_tip(0) <= place_314_top;
  cbr_14_oper_exitcond131_bool_d_req_tip(1) <= place_319_top;
  cbr_15_oper_tmp_d_92_bool_d_req_tip(0) <= place_360_top;
  cbr_16_oper_tmp_d_11348_bool_d_req_tip(0) <= place_389_top;
  cbr_16_oper_tmp_d_11348_bool_d_req_tip(1) <= place_390_top;
  cbr_16_oper_tmp_d_11348_bool_d_req_tip(2) <= place_392_top;
  cbr_17_oper_tmp_d_113_bool_d_req_tip(0) <= place_440_top;
  cbr_17_oper_tmp_d_113_bool_d_req_tip(1) <= place_447_top;
  cbr_17_oper_tmp_d_113_bool_d_req_tip(2) <= place_448_top;
  cbr_17_oper_tmp_d_113_bool_d_req_tip(3) <= place_450_top;
  cbr_18_oper_exitcond142_bool_d_req_tip(0) <= place_453_top;
  cbr_19_oper_tmp_d_149_bool_d_req_tip(0) <= place_469_top;
  cbr_20_oper_tmp_d_14574_bool_d_req_tip(0) <= place_495_top;
  cbr_20_oper_tmp_d_14574_bool_d_req_tip(1) <= place_508_top;
  cbr_20_oper_tmp_d_14574_bool_d_req_tip(2) <= place_513_top;
  cbr_20_oper_tmp_d_14574_bool_d_req_tip(3) <= place_515_top;
  cbr_21_oper_tmp_d_166_bool_d_req_tip(0) <= place_535_top;
  cbr_21_oper_tmp_d_166_bool_d_req_tip(1) <= place_536_top;
  cbr_22_oper_tmp_d_14578_bool_d_req_tip(0) <= place_540_top;
  cbr_22_oper_tmp_d_14578_bool_d_req_tip(1) <= place_566_top;
  cbr_22_oper_tmp_d_14578_bool_d_req_tip(2) <= place_571_top;
  cbr_22_oper_tmp_d_14578_bool_d_req_tip(3) <= place_573_top;
  cbr_23_oper_tmp_d_14580_bool_d_req_tip(0) <= place_576_top;
  cbr_23_oper_tmp_d_14580_bool_d_req_tip(1) <= place_602_top;
  cbr_23_oper_tmp_d_14580_bool_d_req_tip(2) <= place_607_top;
  cbr_23_oper_tmp_d_14580_bool_d_req_tip(3) <= place_609_top;
  cbr_24_oper_exitcond145_bool_d_req_tip(0) <= place_614_top;
  cbr_25_oper_tmp_d_202_bool_d_req_tip(0) <= place_625_top;
  cbr_25_oper_tmp_d_202_bool_d_req_tip(1) <= place_628_top;
  cbr_25_oper_tmp_d_202_bool_d_req_tip(2) <= place_631_top;
  cbr_26_oper_tmp_d_20299_bool_d_req_tip(0) <= place_658_top;
  cbr_26_oper_tmp_d_20299_bool_d_req_tip(1) <= place_665_top;
  cbr_26_oper_tmp_d_20299_bool_d_req_tip(2) <= place_666_top;
  cbr_26_oper_tmp_d_20299_bool_d_req_tip(3) <= place_668_top;
  cbr_27_oper_exitcond150_bool_d_req_tip(0) <= place_676_top;
  cbr_27_oper_exitcond150_bool_d_req_tip(1) <= place_681_top;
  cbr_28_oper_tmp_d_221_bool_d_req_tip(0) <= place_692_top;
  cbr_28_oper_tmp_d_221_bool_d_req_tip(1) <= place_697_top;
  cbr_29_oper_tmp_d_221111_bool_d_req_tip(0) <= place_729_top;
  cbr_29_oper_tmp_d_221111_bool_d_req_tip(1) <= place_736_top;
  cbr_29_oper_tmp_d_221111_bool_d_req_tip(2) <= place_737_top;
  cbr_29_oper_tmp_d_221111_bool_d_req_tip(3) <= place_739_top;
  cbr_30_oper_exitcond158_bool_d_req_tip(0) <= place_747_top;
  cbr_30_oper_exitcond158_bool_d_req_tip(1) <= place_752_top;
  cbr_6_oper_exitcond_bool_d_req_tip(0) <= place_116_top;
  cbr_6_oper_exitcond_bool_d_req_tip(1) <= place_121_top;
  cbr_6_oper_exitcond_bool_d_req_tip(2) <= place_123_top;
  cbr_7_oper_exitcond120_bool_d_req_tip(0) <= place_128_top;
  cbr_8_oper_tmp_d_16_bool_d_req_tip(0) <= place_132_top;
  cbr_9_oper_tmp_d_1614_bool_d_req_tip(0) <= place_170_top;
  cbr_9_oper_tmp_d_1614_bool_d_req_tip(1) <= place_177_top;
  cbr_9_oper_tmp_d_1614_bool_d_req_tip(2) <= place_178_top;
  cbr_9_oper_tmp_d_1614_bool_d_req_tip(3) <= place_180_top;
  else_d_0_d_entry_tip(0) <= place_54_top;
  else_d_0_to_else_d_1_src_tip(0) <= place_537_top;
  else_d_0_to_then_d_2_src_tip(0) <= place_537_top;
  else_d_1_d_entry_tip(0) <= place_61_top;
  else_d_1_to_loopexit_d_10_src_tip(0) <= place_608_top;
  else_d_1_to_no_exit_d_10_d_backedge_src_tip(0) <= place_608_top;
  fin_tip(0) <= place_83_top;
  indvar118_d_ph_d_ph_mux_1_d_ack_tip(0) <= place_100_top;
  indvar118_d_ph_d_ph_mux_1_d_req0_tip(0) <= place_1_top;
  indvar118_d_ph_d_ph_mux_1_d_req1_tip(0) <= place_99_top;
  indvar121_mux_1_d_ack_tip(0) <= place_136_top;
  indvar121_mux_1_d_req0_tip(0) <= place_138_top;
  indvar121_mux_1_d_req1_tip(0) <= place_9_top;
  indvar123_mux_1_d_ack_tip(0) <= place_232_top;
  indvar123_mux_1_d_req0_tip(0) <= place_234_top;
  indvar123_mux_1_d_req1_tip(0) <= place_231_top;
  indvar126_mux_1_d_ack_tip(0) <= place_273_top;
  indvar126_mux_1_d_req0_tip(0) <= place_275_top;
  indvar126_mux_1_d_req1_tip(0) <= place_269_top;
  indvar129_mux_1_d_ack_tip(0) <= place_184_top;
  indvar129_mux_1_d_req0_tip(0) <= place_186_top;
  indvar129_mux_1_d_req1_tip(0) <= place_183_top;
  indvar132_mux_1_d_ack_tip(0) <= place_399_top;
  indvar132_mux_1_d_req0_tip(0) <= place_401_top;
  indvar132_mux_1_d_req1_tip(0) <= place_40_top;
  indvar134_mux_1_d_ack_tip(0) <= place_323_top;
  indvar134_mux_1_d_req0_tip(0) <= place_325_top;
  indvar134_mux_1_d_req1_tip(0) <= place_322_top;
  indvar138_mux_1_d_ack_tip(0) <= place_349_top;
  indvar138_mux_1_d_req0_tip(0) <= place_351_top;
  indvar138_mux_1_d_req1_tip(0) <= place_396_top;
  indvar143_mux_1_d_ack_tip(0) <= place_457_top;
  indvar143_mux_1_d_req0_tip(0) <= place_459_top;
  indvar143_mux_1_d_req1_tip(0) <= place_48_top;
  indvar146_mux_1_d_ack_tip(0) <= place_635_top;
  indvar146_mux_1_d_req0_tip(0) <= place_637_top;
  indvar146_mux_1_d_req1_tip(0) <= place_69_top;
  indvar148_mux_1_d_ack_tip(0) <= place_618_top;
  indvar148_mux_1_d_req0_tip(0) <= place_620_top;
  indvar148_mux_1_d_req1_tip(0) <= place_617_top;
  indvar151_mux_1_d_ack_tip(0) <= place_701_top;
  indvar151_mux_1_d_req0_tip(0) <= place_703_top;
  indvar151_mux_1_d_req1_tip(0) <= place_77_top;
  indvar153_mux_1_d_ack_tip(0) <= place_685_top;
  indvar153_mux_1_d_req0_tip(0) <= place_687_top;
  indvar153_mux_1_d_req1_tip(0) <= place_684_top;
  indvar_mux_1_d_ack_tip(0) <= place_105_top;
  indvar_mux_1_d_req0_tip(0) <= place_107_top;
  indvar_mux_1_d_req1_tip(0) <= place_101_top;
  init_tip(0) <= place_84_top;
  j_d_3_d_in_d_ph_mux_1_d_ack_tip(0) <= place_188_top;
  j_d_3_d_in_d_ph_mux_1_d_req0_tip(0) <= place_190_top;
  j_d_3_d_in_d_ph_mux_1_d_req1_tip(0) <= place_187_top;
  j_d_3_d_in_mux_1_d_ack_tip(0) <= place_209_top;
  j_d_3_d_in_mux_1_d_req0_tip(0) <= place_211_top;
  j_d_3_d_in_mux_1_d_req1_tip(0) <= place_208_top;
  j_d_9_d_2_d_be_mux_1_d_ack_tip(0) <= place_520_top;
  j_d_9_d_2_d_be_mux_1_d_req0_tip(0) <= place_522_top;
  j_d_9_d_2_d_be_mux_1_d_req1_tip(0) <= place_519_top;
  j_d_9_d_2_d_be_mux_2_d_ack_tip(0) <= place_517_top;
  j_d_9_d_2_d_be_mux_2_d_req0_tip(0) <= place_521_top;
  j_d_9_d_2_d_be_mux_2_d_req1_tip(0) <= place_516_top;
  j_d_9_d_2_mux_1_d_ack_tip(0) <= place_464_top;
  j_d_9_d_2_mux_1_d_req0_tip(0) <= place_462_top;
  j_d_9_d_2_mux_1_d_req1_tip(0) <= place_518_top;
  k_d_1_d_in_d_ph_mux_1_d_ack_tip(0) <= place_327_top;
  k_d_1_d_in_d_ph_mux_1_d_req0_tip(0) <= place_329_top;
  k_d_1_d_in_d_ph_mux_1_d_req1_tip(0) <= place_326_top;
  k_d_2_d_3_mux_1_d_ack_tip(0) <= place_673_top;
  k_d_2_d_3_mux_1_d_req0_tip(0) <= place_675_top;
  k_d_2_d_3_mux_1_d_req1_tip(0) <= place_671_top;
  k_d_3_d_0_mux_1_d_ack_tip(0) <= place_622_top;
  k_d_3_d_0_mux_1_d_req0_tip(0) <= place_624_top;
  k_d_3_d_0_mux_1_d_req1_tip(0) <= place_621_top;
  k_d_4_d_3_mux_1_d_ack_tip(0) <= place_744_top;
  k_d_4_d_3_mux_1_d_req0_tip(0) <= place_746_top;
  k_d_4_d_3_mux_1_d_req1_tip(0) <= place_742_top;
  k_d_5_d_0_mux_1_d_ack_tip(0) <= place_689_top;
  k_d_5_d_0_mux_1_d_req0_tip(0) <= place_691_top;
  k_d_5_d_0_mux_1_d_req1_tip(0) <= place_688_top;
  load_A_d_ack_tip(0) <= place_89_top;
  load_A_d_req_tip(0) <= place_88_top;
  load_ccoeff_d_ack_tip(0) <= place_93_top;
  load_ccoeff_d_req_tip(0) <= place_92_top;
  load_l_array_d_ack_tip(0) <= place_95_top;
  load_l_array_d_req_tip(0) <= place_94_top;
  load_noofelem_d_ack_tip(0) <= place_87_top;
  load_noofelem_d_req_tip(0) <= place_86_top;
  load_rcoeff_d_ack_tip(0) <= place_91_top;
  load_rcoeff_d_req_tip(0) <= place_90_top;
  load_start_call_divide_0_return_d_ack_tip(0) <= place_384_top;
  load_start_call_divide_0_return_d_req_tip(0) <= place_383_top;
  load_tmp_d_103_d_ack_tip(0) <= place_370_top;
  load_tmp_d_103_d_req_tip(0) <= place_371_top;
  load_tmp_d_108_d_ack_tip(0) <= place_372_top;
  load_tmp_d_108_d_req_tip(0) <= place_373_top;
  load_tmp_d_108_d_req_tip(1) <= place_374_top;
  load_tmp_d_123_d_ack_tip(0) <= place_415_top;
  load_tmp_d_123_d_req_tip(0) <= place_416_top;
  load_tmp_d_128_d_ack_tip(0) <= place_417_top;
  load_tmp_d_128_d_req_tip(0) <= place_418_top;
  load_tmp_d_128_d_req_tip(1) <= place_419_top;
  load_tmp_d_133_d_ack_tip(0) <= place_427_top;
  load_tmp_d_133_d_req_tip(0) <= place_428_top;
  load_tmp_d_133_d_req_tip(1) <= place_429_top;
  load_tmp_d_159_d_ack_tip(0) <= place_489_top;
  load_tmp_d_159_d_req_tip(0) <= place_490_top;
  load_tmp_d_180_d_ack_tip(0) <= place_559_top;
  load_tmp_d_180_d_req_tip(0) <= place_560_top;
  load_tmp_d_180_d_req_tip(1) <= place_561_top;
  load_tmp_d_193_d_ack_tip(0) <= place_595_top;
  load_tmp_d_193_d_req_tip(0) <= place_596_top;
  load_tmp_d_193_d_req_tip(1) <= place_597_top;
  load_tmp_d_211_d_ack_tip(0) <= place_652_top;
  load_tmp_d_211_d_req_tip(0) <= place_653_top;
  load_tmp_d_21_d_ack_tip(0) <= place_143_top;
  load_tmp_d_21_d_req_tip(0) <= place_144_top;
  load_tmp_d_230_d_ack_tip(0) <= place_723_top;
  load_tmp_d_230_d_req_tip(0) <= place_724_top;
  load_tmp_d_26_d_ack_tip(0) <= place_147_top;
  load_tmp_d_26_d_req_tip(0) <= place_148_top;
  load_tmp_d_26_d_req_tip(1) <= place_149_top;
  load_tmp_d_31_d_ack_tip(0) <= place_163_top;
  load_tmp_d_31_d_req_tip(0) <= place_164_top;
  load_tmp_d_31_d_req_tip(1) <= place_165_top;
  load_tmp_d_48_d_ack_tip(0) <= place_251_top;
  load_tmp_d_48_d_req_tip(0) <= place_252_top;
  load_tmp_d_53_d_ack_tip(0) <= place_225_top;
  load_tmp_d_53_d_req_tip(0) <= place_226_top;
  load_tmp_d_66_d_ack_tip(0) <= place_282_top;
  load_tmp_d_66_d_req_tip(0) <= place_283_top;
  load_tmp_d_75_d_ack_tip(0) <= place_292_top;
  load_tmp_d_75_d_req_tip(0) <= place_293_top;
  load_tmp_d_75_d_req_tip(1) <= place_294_top;
  load_u_array_d_ack_tip(0) <= place_97_top;
  load_u_array_d_req_tip(0) <= place_96_top;
  loopentry_d_12_d_entry_tip(0) <= place_66_top;
  loopentry_d_12_d_loopexit_to_loopentry_d_12_src_tip(0) <= place_65_top;
  loopentry_d_12_d_pre_tip(0) <= place_619_top;
  loopentry_d_12_d_pre_tip(1) <= place_623_top;
  loopentry_d_12_to_loopexit_d_12_src_tip(0) <= place_632_top;
  loopentry_d_12_to_no_exit_d_12_d_preheader_src_tip(0) <= place_632_top;
  loopentry_d_14_d_entry_tip(0) <= place_75_top;
  loopentry_d_14_d_loopexit_to_loopentry_d_14_src_tip(0) <= place_74_top;
  loopentry_d_14_d_pre_tip(0) <= place_686_top;
  loopentry_d_14_d_pre_tip(1) <= place_690_top;
  loopentry_d_14_to_loopexit_d_14_src_tip(0) <= place_698_top;
  loopentry_d_14_to_no_exit_d_14_d_preheader_src_tip(0) <= place_698_top;
  loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_tip(0) <= place_133_top;
  loopentry_d_2_to_no_exit_d_2_d_preheader_src_tip(0) <= place_133_top;
  loopentry_d_4_d_entry_tip(0) <= place_17_top;
  loopentry_d_4_d_loopexit_to_loopentry_d_4_src_tip(0) <= place_25_top;
  loopentry_d_4_d_outer_d_entry_tip(0) <= place_16_top;
  loopentry_d_4_d_outer_d_pre_tip(0) <= place_185_top;
  loopentry_d_4_d_outer_d_pre_tip(1) <= place_189_top;
  loopentry_d_4_d_outer_d_pre_tip(2) <= place_194_top;
  loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_tip(0) <= place_14_top;
  loopentry_d_4_d_outer_to_loopentry_d_4_src_tip(0) <= place_191_top;
  loopentry_d_4_d_outer_to_loopentry_d_4_src_tip(1) <= place_196_top;
  loopentry_d_4_d_outer_to_loopentry_d_4_src_tip(2) <= place_199_top;
  loopentry_d_4_d_outer_to_loopentry_d_4_src_tip(3) <= place_206_top;
  loopentry_d_4_d_pre_tip(0) <= place_210_top;
  loopentry_d_4_d_pre_tip(1) <= place_214_top;
  loopentry_d_4_to_no_exit_d_4_d_preheader_src_tip(0) <= place_222_top;
  loopentry_d_4_to_no_exit_d_5_d_preheader_src_tip(0) <= place_222_top;
  loopentry_d_7_d_outer_d_entry_tip(0) <= place_33_top;
  loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_tip(0) <= place_32_top;
  loopentry_d_7_d_outer_d_pre_tip(0) <= place_324_top;
  loopentry_d_7_d_outer_d_pre_tip(1) <= place_328_top;
  loopentry_d_7_d_outer_to_loopentry_d_7_src_tip(0) <= place_330_top;
  loopentry_d_7_d_outer_to_loopentry_d_7_src_tip(1) <= place_339_top;
  loopentry_d_7_d_outer_to_loopentry_d_7_src_tip(2) <= place_344_top;
  loopentry_d_7_d_outer_to_loopentry_d_7_src_tip(3) <= place_347_top;
  loopentry_d_7_to_loopexit_d_7_src_tip(0) <= place_361_top;
  loopentry_d_7_to_no_exit_d_7_src_tip(0) <= place_361_top;
  loopexit_d_10_to_loopentry_d_12_d_loopexit_src_tip(0) <= place_615_top;
  loopexit_d_10_to_no_exit_d_10_d_outer_src_tip(0) <= place_615_top;
  loopexit_d_12_d_entry_tip(0) <= place_674_top;
  loopexit_d_12_to_loopentry_d_12_src_tip(0) <= place_682_top;
  loopexit_d_12_to_loopentry_d_14_d_loopexit_src_tip(0) <= place_682_top;
  loopexit_d_14_d_entry_tip(0) <= place_745_top;
  loopexit_d_14_to_loopentry_d_14_src_tip(0) <= place_753_top;
  loopexit_d_14_to_return_src_tip(0) <= place_753_top;
  loopexit_d_1_to_loopentry_d_2_src_tip(0) <= place_129_top;
  loopexit_d_1_to_no_exit_d_1_d_outer_src_tip(0) <= place_129_top;
  loopexit_d_5_d_entry_tip(0) <= place_30_top;
  loopexit_d_5_to_loopentry_d_4_d_outer_src_tip(0) <= place_320_top;
  loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_tip(0) <= place_320_top;
  loopexit_d_7_to_loopentry_d_7_d_outer_src_tip(0) <= place_454_top;
  loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_tip(0) <= place_454_top;
  maxcoeff_d_2_d_2_mux_1_d_ack_tip(0) <= place_236_top;
  maxcoeff_d_2_d_2_mux_1_d_req0_tip(0) <= place_238_top;
  maxcoeff_d_2_d_2_mux_1_d_req1_tip(0) <= place_235_top;
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_tip(0) <= place_268_top;
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_tip(0) <= place_270_top;
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_tip(0) <= place_27_top;
  maxcoeff_d_2_d_ph_mux_1_d_ack_tip(0) <= place_193_top;
  maxcoeff_d_2_d_ph_mux_1_d_req0_tip(0) <= place_195_top;
  maxcoeff_d_2_d_ph_mux_1_d_req1_tip(0) <= place_192_top;
  maxcoeff_d_2_mux_1_d_ack_tip(0) <= place_213_top;
  maxcoeff_d_2_mux_1_d_req0_tip(0) <= place_215_top;
  maxcoeff_d_2_mux_1_d_req1_tip(0) <= place_212_top;
  no_exit_d_10_to_else_d_0_src_tip(0) <= place_470_top;
  no_exit_d_10_to_then_d_1_src_tip(0) <= place_470_top;
  no_exit_d_12_d_entry_tip(0) <= place_636_top;
  no_exit_d_12_to_loopexit_d_12_d_loopexit_src_tip(0) <= place_667_top;
  no_exit_d_12_to_no_exit_d_12_src_tip(0) <= place_667_top;
  no_exit_d_14_d_entry_tip(0) <= place_702_top;
  no_exit_d_14_to_loopexit_d_14_d_loopexit_src_tip(0) <= place_738_top;
  no_exit_d_14_to_no_exit_d_14_src_tip(0) <= place_738_top;
  no_exit_d_1_d_entry_tip(0) <= place_106_top;
  no_exit_d_1_to_loopexit_d_1_src_tip(0) <= place_122_top;
  no_exit_d_1_to_no_exit_d_1_src_tip(0) <= place_122_top;
  no_exit_d_2_d_entry_tip(0) <= place_137_top;
  no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_tip(0) <= place_179_top;
  no_exit_d_2_to_no_exit_d_2_src_tip(0) <= place_179_top;
  no_exit_d_4_d_entry_tip(0) <= place_22_top;
  no_exit_d_4_d_pre_tip(0) <= place_233_top;
  no_exit_d_4_d_pre_tip(1) <= place_237_top;
  no_exit_d_4_d_preheader_d_entry_tip(0) <= place_20_top;
  no_exit_d_4_d_preheader_to_no_exit_d_4_src_tip(0) <= place_227_top;
  no_exit_d_4_d_preheader_to_no_exit_d_4_src_tip(1) <= place_230_top;
  no_exit_d_4_to_loopentry_d_4_d_loopexit_src_tip(0) <= place_256_top;
  no_exit_d_4_to_then_d_0_src_tip(0) <= place_256_top;
  no_exit_d_5_d_entry_tip(0) <= place_274_top;
  no_exit_d_5_to_loopexit_d_5_src_tip(0) <= place_310_top;
  no_exit_d_5_to_no_exit_d_5_src_tip(0) <= place_310_top;
  no_exit_d_7_d_entry_tip(0) <= place_36_top;
  no_exit_d_7_to_loopentry_d_7_d_backedge_src_tip(0) <= place_391_top;
  no_exit_d_7_to_no_exit_d_8_d_preheader_src_tip(0) <= place_391_top;
  no_exit_d_8_d_entry_tip(0) <= place_400_top;
  no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_tip(0) <= place_449_top;
  no_exit_d_8_to_no_exit_d_8_src_tip(0) <= place_449_top;
  oper_exitcond120_bool_d_ack_tip(0) <= place_126_top;
  oper_exitcond120_bool_d_req_tip(0) <= place_127_top;
  oper_exitcond128_bool_d_ack_tip(0) <= place_307_top;
  oper_exitcond128_bool_d_req_tip(0) <= place_308_top;
  oper_exitcond131_bool_d_ack_tip(0) <= place_317_top;
  oper_exitcond131_bool_d_req_tip(0) <= place_318_top;
  oper_exitcond142_bool_d_ack_tip(0) <= place_451_top;
  oper_exitcond142_bool_d_req_tip(0) <= place_38_top;
  oper_exitcond145_bool_d_ack_tip(0) <= place_612_top;
  oper_exitcond145_bool_d_req_tip(0) <= place_613_top;
  oper_exitcond150_bool_d_ack_tip(0) <= place_679_top;
  oper_exitcond150_bool_d_req_tip(0) <= place_680_top;
  oper_exitcond158_bool_d_ack_tip(0) <= place_750_top;
  oper_exitcond158_bool_d_req_tip(0) <= place_751_top;
  oper_exitcond_bool_d_ack_tip(0) <= place_119_top;
  oper_exitcond_bool_d_req_tip(0) <= place_120_top;
  oper_inc_d_11_int_d_ack_tip(0) <= place_669_top;
  oper_inc_d_11_int_d_req_tip(0) <= place_72_top;
  oper_inc_d_12_int_d_ack_tip(0) <= place_659_top;
  oper_inc_d_12_int_d_req_tip(0) <= place_660_top;
  oper_inc_d_14_int_d_ack_tip(0) <= place_740_top;
  oper_inc_d_14_int_d_req_tip(0) <= place_81_top;
  oper_inc_d_15_int_d_ack_tip(0) <= place_730_top;
  oper_inc_d_15_int_d_req_tip(0) <= place_731_top;
  oper_inc_d_2_int_d_ack_tip(0) <= place_171_top;
  oper_inc_d_2_int_d_req_tip(0) <= place_172_top;
  oper_inc_d_5_int_d_ack_tip(0) <= place_312_top;
  oper_inc_d_5_int_d_req_tip(0) <= place_313_top;
  oper_inc_d_960_int_d_ack_tip(0) <= place_509_top;
  oper_inc_d_960_int_d_req_tip(0) <= place_510_top;
  oper_inc_d_976_int_d_ack_tip(0) <= place_567_top;
  oper_inc_d_976_int_d_req_tip(0) <= place_568_top;
  oper_inc_d_9_int_d_ack_tip(0) <= place_603_top;
  oper_inc_d_9_int_d_req_tip(0) <= place_604_top;
  oper_indvar_d_next119_uint_d_ack_tip(0) <= place_124_top;
  oper_indvar_d_next119_uint_d_req_tip(0) <= place_5_top;
  oper_indvar_d_next122_uint_d_ack_tip(0) <= place_175_top;
  oper_indvar_d_next122_uint_d_req_tip(0) <= place_176_top;
  oper_indvar_d_next124_uint_d_ack_tip(0) <= place_261_top;
  oper_indvar_d_next124_uint_d_req_tip(0) <= place_262_top;
  oper_indvar_d_next127_uint_d_ack_tip(0) <= place_305_top;
  oper_indvar_d_next127_uint_d_req_tip(0) <= place_306_top;
  oper_indvar_d_next130_uint_d_ack_tip(0) <= place_315_top;
  oper_indvar_d_next130_uint_d_req_tip(0) <= place_316_top;
  oper_indvar_d_next133_uint_d_ack_tip(0) <= place_445_top;
  oper_indvar_d_next133_uint_d_req_tip(0) <= place_446_top;
  oper_indvar_d_next139_uint_d_ack_tip(0) <= place_394_top;
  oper_indvar_d_next139_uint_d_req_tip(0) <= place_46_top;
  oper_indvar_d_next144_uint_d_ack_tip(0) <= place_610_top;
  oper_indvar_d_next144_uint_d_req_tip(0) <= place_63_top;
  oper_indvar_d_next147_uint_d_ack_tip(0) <= place_663_top;
  oper_indvar_d_next147_uint_d_req_tip(0) <= place_664_top;
  oper_indvar_d_next149_uint_d_ack_tip(0) <= place_677_top;
  oper_indvar_d_next149_uint_d_req_tip(0) <= place_678_top;
  oper_indvar_d_next152_uint_d_ack_tip(0) <= place_734_top;
  oper_indvar_d_next152_uint_d_req_tip(0) <= place_735_top;
  oper_indvar_d_next157_uint_d_ack_tip(0) <= place_748_top;
  oper_indvar_d_next157_uint_d_req_tip(0) <= place_749_top;
  oper_indvar_d_next_uint_d_ack_tip(0) <= place_117_top;
  oper_indvar_d_next_uint_d_req_tip(0) <= place_118_top;
  oper_j_d_321_int_d_ack_tip(0) <= place_257_top;
  oper_j_d_321_int_d_req_tip(0) <= place_258_top;
  oper_j_d_3_int_d_ack_tip(0) <= place_217_top;
  oper_j_d_3_int_d_req_tip(0) <= place_218_top;
  oper_j_d_746_int_d_ack_tip(0) <= place_340_top;
  oper_j_d_746_int_d_req_tip(0) <= place_341_top;
  oper_j_d_7_int_d_ack_tip(0) <= place_441_top;
  oper_j_d_7_int_d_req_tip(0) <= place_442_top;
  oper_k_d_1_d_in_int_d_ack_tip(0) <= place_354_top;
  oper_k_d_1_d_in_int_d_req_tip(0) <= place_355_top;
  oper_k_d_1_int_d_ack_tip(0) <= place_356_top;
  oper_k_d_1_int_d_req_tip(0) <= place_357_top;
  oper_k_d_2_d_2_int_d_ack_tip(0) <= place_640_top;
  oper_k_d_2_d_2_int_d_req_tip(0) <= place_641_top;
  oper_k_d_4_d_2_int_d_ack_tip(0) <= place_710_top;
  oper_k_d_4_d_2_int_d_req_tip(0) <= place_711_top;
  oper_tmp_d_107_d_id_d_1_uint_d_ack_tip(0) <= place_333_top;
  oper_tmp_d_107_d_id_d_1_uint_d_req_tip(0) <= place_334_top;
  oper_tmp_d_107_d_lvl_d_1_uint_d_ack_tip(0) <= place_335_top;
  oper_tmp_d_107_d_lvl_d_1_uint_d_req_tip(0) <= place_336_top;
  oper_tmp_d_107_d_lvl_d_2_uint_d_ack_tip(0) <= place_337_top;
  oper_tmp_d_107_d_lvl_d_2_uint_d_req_tip(0) <= place_338_top;
  oper_tmp_d_11348_bool_d_ack_tip(0) <= place_342_top;
  oper_tmp_d_11348_bool_d_req_tip(0) <= place_343_top;
  oper_tmp_d_113_bool_d_ack_tip(0) <= place_443_top;
  oper_tmp_d_113_bool_d_req_tip(0) <= place_444_top;
  oper_tmp_d_118_d_id_d_1_uint_d_ack_tip(0) <= place_408_top;
  oper_tmp_d_118_d_id_d_1_uint_d_req_tip(0) <= place_409_top;
  oper_tmp_d_118_d_lvl_d_1_uint_d_ack_tip(0) <= place_410_top;
  oper_tmp_d_118_d_lvl_d_1_uint_d_req_tip(0) <= place_411_top;
  oper_tmp_d_118_d_lvl_d_2_uint_d_ack_tip(0) <= place_412_top;
  oper_tmp_d_118_d_lvl_d_2_uint_d_req_tip(0) <= place_413_top;
  oper_tmp_d_118_d_lvl_d_2_uint_d_req_tip(1) <= place_414_top;
  oper_tmp_d_11_d_id_d_1_uint_d_ack_tip(0) <= place_108_top;
  oper_tmp_d_11_d_id_d_1_uint_d_req_tip(0) <= place_109_top;
  oper_tmp_d_11_d_lvl_d_1_uint_d_ack_tip(0) <= place_110_top;
  oper_tmp_d_11_d_lvl_d_1_uint_d_req_tip(0) <= place_111_top;
  oper_tmp_d_11_d_lvl_d_2_uint_d_ack_tip(0) <= place_112_top;
  oper_tmp_d_11_d_lvl_d_2_uint_d_req_tip(0) <= place_113_top;
  oper_tmp_d_125_uint_d_ack_tip(0) <= place_240_top;
  oper_tmp_d_125_uint_d_req_tip(0) <= place_241_top;
  oper_tmp_d_132_d_id_d_1_uint_d_ack_tip(0) <= place_420_top;
  oper_tmp_d_132_d_id_d_1_uint_d_req_tip(0) <= place_421_top;
  oper_tmp_d_132_d_lvl_d_1_uint_d_ack_tip(0) <= place_422_top;
  oper_tmp_d_132_d_lvl_d_1_uint_d_req_tip(0) <= place_423_top;
  oper_tmp_d_132_d_lvl_d_2_uint_d_ack_tip(0) <= place_424_top;
  oper_tmp_d_132_d_lvl_d_2_uint_d_req_tip(0) <= place_425_top;
  oper_tmp_d_132_d_lvl_d_2_uint_d_req_tip(1) <= place_426_top;
  oper_tmp_d_134_float_d_ack_tip(0) <= place_430_top;
  oper_tmp_d_134_float_d_req_tip(0) <= place_431_top;
  oper_tmp_d_134_float_d_req_tip(1) <= place_432_top;
  oper_tmp_d_135_float_d_ack_tip(0) <= place_433_top;
  oper_tmp_d_135_float_d_req_tip(0) <= place_434_top;
  oper_tmp_d_135_float_d_req_tip(1) <= place_435_top;
  oper_tmp_d_136_uint_d_ack_tip(0) <= place_345_top;
  oper_tmp_d_136_uint_d_req_tip(0) <= place_346_top;
  oper_tmp_d_137_uint_d_ack_tip(0) <= place_402_top;
  oper_tmp_d_137_uint_d_req_tip(0) <= place_403_top;
  oper_tmp_d_14574_bool_d_ack_tip(0) <= place_511_top;
  oper_tmp_d_14574_bool_d_req_tip(0) <= place_512_top;
  oper_tmp_d_14578_bool_d_ack_tip(0) <= place_569_top;
  oper_tmp_d_14578_bool_d_req_tip(0) <= place_570_top;
  oper_tmp_d_14580_bool_d_ack_tip(0) <= place_605_top;
  oper_tmp_d_14580_bool_d_req_tip(0) <= place_606_top;
  oper_tmp_d_149_bool_d_ack_tip(0) <= place_467_top;
  oper_tmp_d_149_bool_d_req_tip(0) <= place_465_top;
  oper_tmp_d_154_d_id_d_1_uint_d_ack_tip(0) <= place_471_top;
  oper_tmp_d_154_d_id_d_1_uint_d_req_tip(0) <= place_472_top;
  oper_tmp_d_154_d_lvl_d_1_uint_d_ack_tip(0) <= place_473_top;
  oper_tmp_d_154_d_lvl_d_1_uint_d_req_tip(0) <= place_474_top;
  oper_tmp_d_154_d_lvl_d_2_uint_d_ack_tip(0) <= place_477_top;
  oper_tmp_d_154_d_lvl_d_2_uint_d_req_tip(0) <= place_478_top;
  oper_tmp_d_154_d_lvl_d_2_uint_d_req_tip(1) <= place_479_top;
  oper_tmp_d_155_uint_d_ack_tip(0) <= place_706_top;
  oper_tmp_d_155_uint_d_req_tip(0) <= place_707_top;
  oper_tmp_d_158_d_id_d_1_uint_d_ack_tip(0) <= place_480_top;
  oper_tmp_d_158_d_id_d_1_uint_d_req_tip(0) <= place_481_top;
  oper_tmp_d_158_d_lvl_d_1_uint_d_ack_tip(0) <= place_482_top;
  oper_tmp_d_158_d_lvl_d_1_uint_d_req_tip(0) <= place_483_top;
  oper_tmp_d_158_d_lvl_d_2_uint_d_ack_tip(0) <= place_486_top;
  oper_tmp_d_158_d_lvl_d_2_uint_d_req_tip(0) <= place_487_top;
  oper_tmp_d_158_d_lvl_d_2_uint_d_req_tip(1) <= place_488_top;
  oper_tmp_d_1614_bool_d_ack_tip(0) <= place_173_top;
  oper_tmp_d_1614_bool_d_req_tip(0) <= place_174_top;
  oper_tmp_d_163_d_id_d_1_uint_d_ack_tip(0) <= place_496_top;
  oper_tmp_d_163_d_id_d_1_uint_d_req_tip(0) <= place_497_top;
  oper_tmp_d_163_d_lvl_d_1_uint_d_ack_tip(0) <= place_498_top;
  oper_tmp_d_163_d_lvl_d_1_uint_d_req_tip(0) <= place_499_top;
  oper_tmp_d_163_d_lvl_d_2_uint_d_ack_tip(0) <= place_502_top;
  oper_tmp_d_163_d_lvl_d_2_uint_d_req_tip(0) <= place_503_top;
  oper_tmp_d_163_d_lvl_d_2_uint_d_req_tip(1) <= place_504_top;
  oper_tmp_d_166_bool_d_ack_tip(0) <= place_524_top;
  oper_tmp_d_166_bool_d_req_tip(0) <= place_525_top;
  oper_tmp_d_16_bool_d_ack_tip(0) <= place_130_top;
  oper_tmp_d_16_bool_d_req_tip(0) <= place_7_top;
  oper_tmp_d_171_d_id_d_1_uint_d_ack_tip(0) <= place_526_top;
  oper_tmp_d_171_d_id_d_1_uint_d_req_tip(0) <= place_527_top;
  oper_tmp_d_171_d_lvl_d_1_uint_d_ack_tip(0) <= place_528_top;
  oper_tmp_d_171_d_lvl_d_1_uint_d_req_tip(0) <= place_529_top;
  oper_tmp_d_171_d_lvl_d_2_uint_d_ack_tip(0) <= place_532_top;
  oper_tmp_d_171_d_lvl_d_2_uint_d_req_tip(0) <= place_533_top;
  oper_tmp_d_171_d_lvl_d_2_uint_d_req_tip(1) <= place_534_top;
  oper_tmp_d_175_d_id_d_1_uint_d_ack_tip(0) <= place_541_top;
  oper_tmp_d_175_d_id_d_1_uint_d_req_tip(0) <= place_542_top;
  oper_tmp_d_175_d_lvl_d_1_uint_d_ack_tip(0) <= place_543_top;
  oper_tmp_d_175_d_lvl_d_1_uint_d_req_tip(0) <= place_544_top;
  oper_tmp_d_175_d_lvl_d_2_uint_d_ack_tip(0) <= place_547_top;
  oper_tmp_d_175_d_lvl_d_2_uint_d_req_tip(0) <= place_548_top;
  oper_tmp_d_175_d_lvl_d_2_uint_d_req_tip(1) <= place_549_top;
  oper_tmp_d_179_d_id_d_1_uint_d_ack_tip(0) <= place_550_top;
  oper_tmp_d_179_d_id_d_1_uint_d_req_tip(0) <= place_551_top;
  oper_tmp_d_179_d_lvl_d_1_uint_d_ack_tip(0) <= place_552_top;
  oper_tmp_d_179_d_lvl_d_1_uint_d_req_tip(0) <= place_553_top;
  oper_tmp_d_179_d_lvl_d_2_uint_d_ack_tip(0) <= place_556_top;
  oper_tmp_d_179_d_lvl_d_2_uint_d_req_tip(0) <= place_557_top;
  oper_tmp_d_179_d_lvl_d_2_uint_d_req_tip(1) <= place_558_top;
  oper_tmp_d_188_d_id_d_1_uint_d_ack_tip(0) <= place_577_top;
  oper_tmp_d_188_d_id_d_1_uint_d_req_tip(0) <= place_578_top;
  oper_tmp_d_188_d_lvl_d_1_uint_d_ack_tip(0) <= place_579_top;
  oper_tmp_d_188_d_lvl_d_1_uint_d_req_tip(0) <= place_580_top;
  oper_tmp_d_188_d_lvl_d_2_uint_d_ack_tip(0) <= place_583_top;
  oper_tmp_d_188_d_lvl_d_2_uint_d_req_tip(0) <= place_584_top;
  oper_tmp_d_188_d_lvl_d_2_uint_d_req_tip(1) <= place_585_top;
  oper_tmp_d_192_d_id_d_1_uint_d_ack_tip(0) <= place_586_top;
  oper_tmp_d_192_d_id_d_1_uint_d_req_tip(0) <= place_587_top;
  oper_tmp_d_192_d_lvl_d_1_uint_d_ack_tip(0) <= place_588_top;
  oper_tmp_d_192_d_lvl_d_1_uint_d_req_tip(0) <= place_589_top;
  oper_tmp_d_192_d_lvl_d_2_uint_d_ack_tip(0) <= place_592_top;
  oper_tmp_d_192_d_lvl_d_2_uint_d_req_tip(0) <= place_593_top;
  oper_tmp_d_192_d_lvl_d_2_uint_d_req_tip(1) <= place_594_top;
  oper_tmp_d_20299_bool_d_ack_tip(0) <= place_661_top;
  oper_tmp_d_20299_bool_d_req_tip(0) <= place_662_top;
  oper_tmp_d_202_bool_d_ack_tip(0) <= place_629_top;
  oper_tmp_d_202_bool_d_req_tip(0) <= place_630_top;
  oper_tmp_d_206_d_lvl_d_0_uint_d_ack_tip(0) <= place_644_top;
  oper_tmp_d_206_d_lvl_d_0_uint_d_req_tip(0) <= place_645_top;
  oper_tmp_d_20_d_lvl_d_0_uint_d_ack_tip(0) <= place_141_top;
  oper_tmp_d_20_d_lvl_d_0_uint_d_req_tip(0) <= place_142_top;
  oper_tmp_d_210_d_id_d_1_uint_d_ack_tip(0) <= place_646_top;
  oper_tmp_d_210_d_id_d_1_uint_d_req_tip(0) <= place_647_top;
  oper_tmp_d_210_d_lvl_d_1_uint_d_ack_tip(0) <= place_648_top;
  oper_tmp_d_210_d_lvl_d_1_uint_d_req_tip(0) <= place_649_top;
  oper_tmp_d_210_d_lvl_d_2_uint_d_ack_tip(0) <= place_650_top;
  oper_tmp_d_210_d_lvl_d_2_uint_d_req_tip(0) <= place_651_top;
  oper_tmp_d_221111_bool_d_ack_tip(0) <= place_732_top;
  oper_tmp_d_221111_bool_d_req_tip(0) <= place_733_top;
  oper_tmp_d_221_bool_d_ack_tip(0) <= place_695_top;
  oper_tmp_d_221_bool_d_req_tip(0) <= place_696_top;
  oper_tmp_d_225_d_lvl_d_0_uint_d_ack_tip(0) <= place_714_top;
  oper_tmp_d_225_d_lvl_d_0_uint_d_req_tip(0) <= place_715_top;
  oper_tmp_d_229_d_id_d_1_uint_d_ack_tip(0) <= place_716_top;
  oper_tmp_d_229_d_id_d_1_uint_d_req_tip(0) <= place_717_top;
  oper_tmp_d_229_d_lvl_d_1_uint_d_ack_tip(0) <= place_718_top;
  oper_tmp_d_229_d_lvl_d_1_uint_d_req_tip(0) <= place_719_top;
  oper_tmp_d_229_d_lvl_d_2_uint_d_ack_tip(0) <= place_720_top;
  oper_tmp_d_229_d_lvl_d_2_uint_d_req_tip(0) <= place_721_top;
  oper_tmp_d_229_d_lvl_d_2_uint_d_req_tip(1) <= place_722_top;
  oper_tmp_d_25_d_lvl_d_0_uint_d_ack_tip(0) <= place_145_top;
  oper_tmp_d_25_d_lvl_d_0_uint_d_req_tip(0) <= place_146_top;
  oper_tmp_d_27_d_id_d_1_uint_d_ack_tip(0) <= place_152_top;
  oper_tmp_d_27_d_id_d_1_uint_d_req_tip(0) <= place_153_top;
  oper_tmp_d_27_d_lvl_d_1_uint_d_ack_tip(0) <= place_154_top;
  oper_tmp_d_27_d_lvl_d_1_uint_d_req_tip(0) <= place_155_top;
  oper_tmp_d_27_d_lvl_d_2_uint_d_ack_tip(0) <= place_158_top;
  oper_tmp_d_27_d_lvl_d_2_uint_d_req_tip(0) <= place_159_top;
  oper_tmp_d_27_d_lvl_d_2_uint_d_req_tip(1) <= place_160_top;
  oper_tmp_d_30_d_lvl_d_0_uint_d_ack_tip(0) <= place_161_top;
  oper_tmp_d_30_d_lvl_d_0_uint_d_req_tip(0) <= place_162_top;
  oper_tmp_d_4223_bool_d_ack_tip(0) <= place_259_top;
  oper_tmp_d_4223_bool_d_req_tip(0) <= place_260_top;
  oper_tmp_d_42_bool_d_ack_tip(0) <= place_219_top;
  oper_tmp_d_42_bool_d_req_tip(0) <= place_220_top;
  oper_tmp_d_47_d_id_d_1_uint_d_ack_tip(0) <= place_245_top;
  oper_tmp_d_47_d_id_d_1_uint_d_req_tip(0) <= place_246_top;
  oper_tmp_d_47_d_lvl_d_1_uint_d_ack_tip(0) <= place_247_top;
  oper_tmp_d_47_d_lvl_d_1_uint_d_req_tip(0) <= place_248_top;
  oper_tmp_d_47_d_lvl_d_2_uint_d_ack_tip(0) <= place_249_top;
  oper_tmp_d_47_d_lvl_d_2_uint_d_req_tip(0) <= place_250_top;
  oper_tmp_d_52_d_id_d_1_uint_d_ack_tip(0) <= place_200_top;
  oper_tmp_d_52_d_id_d_1_uint_d_req_tip(0) <= place_201_top;
  oper_tmp_d_52_d_lvl_d_1_uint_d_ack_tip(0) <= place_202_top;
  oper_tmp_d_52_d_lvl_d_1_uint_d_req_tip(0) <= place_203_top;
  oper_tmp_d_52_d_lvl_d_2_uint_d_ack_tip(0) <= place_204_top;
  oper_tmp_d_52_d_lvl_d_2_uint_d_req_tip(0) <= place_205_top;
  oper_tmp_d_54_bool_d_ack_tip(0) <= place_253_top;
  oper_tmp_d_54_bool_d_req_tip(0) <= place_254_top;
  oper_tmp_d_65_d_id_d_1_uint_d_ack_tip(0) <= place_276_top;
  oper_tmp_d_65_d_id_d_1_uint_d_req_tip(0) <= place_277_top;
  oper_tmp_d_65_d_lvl_d_1_uint_d_ack_tip(0) <= place_278_top;
  oper_tmp_d_65_d_lvl_d_1_uint_d_req_tip(0) <= place_279_top;
  oper_tmp_d_65_d_lvl_d_2_uint_d_ack_tip(0) <= place_280_top;
  oper_tmp_d_65_d_lvl_d_2_uint_d_req_tip(0) <= place_281_top;
  oper_tmp_d_74_d_id_d_1_uint_d_ack_tip(0) <= place_286_top;
  oper_tmp_d_74_d_id_d_1_uint_d_req_tip(0) <= place_287_top;
  oper_tmp_d_74_d_lvl_d_1_uint_d_ack_tip(0) <= place_288_top;
  oper_tmp_d_74_d_lvl_d_1_uint_d_req_tip(0) <= place_289_top;
  oper_tmp_d_74_d_lvl_d_2_uint_d_ack_tip(0) <= place_290_top;
  oper_tmp_d_74_d_lvl_d_2_uint_d_req_tip(0) <= place_291_top;
  oper_tmp_d_92_bool_d_ack_tip(0) <= place_358_top;
  oper_tmp_d_92_bool_d_req_tip(0) <= place_359_top;
  oper_tmp_d_97_d_id_d_1_uint_d_ack_tip(0) <= place_364_top;
  oper_tmp_d_97_d_id_d_1_uint_d_req_tip(0) <= place_365_top;
  oper_tmp_d_97_d_lvl_d_1_uint_d_ack_tip(0) <= place_366_top;
  oper_tmp_d_97_d_lvl_d_1_uint_d_req_tip(0) <= place_367_top;
  oper_tmp_d_97_d_lvl_d_2_uint_d_ack_tip(0) <= place_368_top;
  oper_tmp_d_97_d_lvl_d_2_uint_d_req_tip(0) <= place_369_top;
  oper_tmp_d_uint_d_ack_tip(0) <= place_228_top;
  oper_tmp_d_uint_d_req_tip(0) <= place_229_top;
  start_call_divide_0_actual_0_wr_d_ack_tip(0) <= place_378_top;
  start_call_divide_0_actual_0_wr_d_req_tip(0) <= place_376_top;
  start_call_divide_0_actual_0_wr_d_req_tip(1) <= place_377_top;
  start_call_divide_0_actual_1_wr_d_ack_tip(0) <= place_381_top;
  start_call_divide_0_actual_1_wr_d_req_tip(0) <= place_379_top;
  start_call_divide_0_actual_1_wr_d_req_tip(1) <= place_380_top;
  start_call_divide_0_d_ack_tip(0) <= place_375_top;
  start_call_divide_0_d_req_tip(0) <= place_382_top;
  store_0_d_ack_tip(0) <= place_114_top;
  store_0_d_req_tip(0) <= place_115_top;
  store_10_d_ack_tip(0) <= place_574_top;
  store_10_d_req_tip(0) <= place_575_top;
  store_11_d_ack_tip(0) <= place_598_top;
  store_11_d_req_tip(0) <= place_599_top;
  store_11_d_req_tip(1) <= place_600_top;
  store_11_d_req_tip(2) <= place_601_top;
  store_12_d_ack_tip(0) <= place_654_top;
  store_12_d_req_tip(0) <= place_655_top;
  store_12_d_req_tip(1) <= place_656_top;
  store_12_d_req_tip(2) <= place_657_top;
  store_13_d_ack_tip(0) <= place_725_top;
  store_13_d_req_tip(0) <= place_726_top;
  store_13_d_req_tip(1) <= place_727_top;
  store_13_d_req_tip(2) <= place_728_top;
  store_1_d_ack_tip(0) <= place_166_top;
  store_1_d_req_tip(0) <= place_167_top;
  store_1_d_req_tip(1) <= place_168_top;
  store_1_d_req_tip(2) <= place_169_top;
  store_2_d_ack_tip(0) <= place_295_top;
  store_2_d_req_tip(0) <= place_296_top;
  store_2_d_req_tip(1) <= place_297_top;
  store_2_d_req_tip(2) <= place_298_top;
  store_3_d_ack_tip(0) <= place_300_top;
  store_3_d_req_tip(0) <= place_301_top;
  store_3_d_req_tip(1) <= place_302_top;
  store_3_d_req_tip(2) <= place_303_top;
  store_4_d_ack_tip(0) <= place_385_top;
  store_4_d_req_tip(0) <= place_386_top;
  store_4_d_req_tip(1) <= place_387_top;
  store_4_d_req_tip(2) <= place_388_top;
  store_5_d_ack_tip(0) <= place_436_top;
  store_5_d_req_tip(0) <= place_437_top;
  store_5_d_req_tip(1) <= place_438_top;
  store_5_d_req_tip(2) <= place_439_top;
  store_6_d_ack_tip(0) <= place_491_top;
  store_6_d_req_tip(0) <= place_492_top;
  store_6_d_req_tip(1) <= place_493_top;
  store_6_d_req_tip(2) <= place_494_top;
  store_7_d_ack_tip(0) <= place_505_top;
  store_7_d_req_tip(0) <= place_506_top;
  store_7_d_req_tip(1) <= place_507_top;
  store_8_d_ack_tip(0) <= place_538_top;
  store_8_d_req_tip(0) <= place_539_top;
  store_9_d_ack_tip(0) <= place_562_top;
  store_9_d_req_tip(0) <= place_563_top;
  store_9_d_req_tip(1) <= place_564_top;
  store_9_d_req_tip(2) <= place_565_top;
  tc_i_d_1_d_0_d_ack_tip(0) <= place_139_top;
  tc_i_d_1_d_0_d_req_tip(0) <= place_140_top;
  tc_i_d_2_d_0_d_ph_d_ack_tip(0) <= place_197_top;
  tc_i_d_2_d_0_d_ph_d_req_tip(0) <= place_198_top;
  tc_i_d_3_d_0_d_ph_d_ack_tip(0) <= place_460_top;
  tc_i_d_3_d_0_d_ph_d_req_tip(0) <= place_458_top;
  tc_i_d_4_d_0_d_ack_tip(0) <= place_626_top;
  tc_i_d_4_d_0_d_req_tip(0) <= place_627_top;
  tc_i_d_5_d_0_d_ack_tip(0) <= place_693_top;
  tc_i_d_5_d_0_d_req_tip(0) <= place_694_top;
  tc_indvar138_d_ack_tip(0) <= place_352_top;
  tc_indvar138_d_req_tip(0) <= place_350_top;
  tc_indvar151_d_ack_tip(0) <= place_704_top;
  tc_indvar151_d_req_tip(0) <= place_705_top;
  tc_j_d_11_d_2_d_ack_tip(0) <= place_638_top;
  tc_j_d_11_d_2_d_req_tip(0) <= place_639_top;
  tc_j_d_13_d_2_d_ack_tip(0) <= place_708_top;
  tc_j_d_13_d_2_d_req_tip(0) <= place_709_top;
  tc_j_d_3_d_2_d_ack_tip(0) <= place_242_top;
  tc_j_d_3_d_2_d_req_tip(0) <= place_243_top;
  tc_j_d_3_d_in_d_ack_tip(0) <= place_223_top;
  tc_j_d_3_d_in_d_req_tip(0) <= place_224_top;
  tc_j_d_7_d_1_d_ack_tip(0) <= place_404_top;
  tc_j_d_7_d_1_d_req_tip(0) <= place_405_top;
  tc_p_d_0_d_0_d_ph_d_ack_tip(0) <= place_331_top;
  tc_p_d_0_d_0_d_ph_d_req_tip(0) <= place_332_top;
  tc_tmp_d_118_d_id_d_1_d_cast_d_ack_tip(0) <= place_406_top;
  tc_tmp_d_118_d_id_d_1_d_cast_d_req_tip(0) <= place_407_top;
  tc_tmp_d_154_d_id_d_2_d_cast_d_ack_tip(0) <= place_475_top;
  tc_tmp_d_154_d_id_d_2_d_cast_d_req_tip(0) <= place_476_top;
  tc_tmp_d_158_d_id_d_2_d_cast_d_ack_tip(0) <= place_484_top;
  tc_tmp_d_158_d_id_d_2_d_cast_d_req_tip(0) <= place_485_top;
  tc_tmp_d_163_d_id_d_2_d_cast_d_ack_tip(0) <= place_500_top;
  tc_tmp_d_163_d_id_d_2_d_cast_d_req_tip(0) <= place_501_top;
  tc_tmp_d_171_d_id_d_2_d_cast_d_ack_tip(0) <= place_530_top;
  tc_tmp_d_171_d_id_d_2_d_cast_d_req_tip(0) <= place_531_top;
  tc_tmp_d_175_d_id_d_2_d_cast_d_ack_tip(0) <= place_545_top;
  tc_tmp_d_175_d_id_d_2_d_cast_d_req_tip(0) <= place_546_top;
  tc_tmp_d_179_d_id_d_2_d_cast_d_ack_tip(0) <= place_554_top;
  tc_tmp_d_179_d_id_d_2_d_cast_d_req_tip(0) <= place_555_top;
  tc_tmp_d_188_d_id_d_2_d_cast_d_ack_tip(0) <= place_581_top;
  tc_tmp_d_188_d_id_d_2_d_cast_d_req_tip(0) <= place_582_top;
  tc_tmp_d_192_d_id_d_2_d_cast_d_ack_tip(0) <= place_590_top;
  tc_tmp_d_192_d_id_d_2_d_cast_d_req_tip(0) <= place_591_top;
  tc_tmp_d_206_d_id_d_0_d_cast_d_ack_tip(0) <= place_642_top;
  tc_tmp_d_206_d_id_d_0_d_cast_d_req_tip(0) <= place_643_top;
  tc_tmp_d_225_d_id_d_0_d_cast_d_ack_tip(0) <= place_712_top;
  tc_tmp_d_225_d_id_d_0_d_cast_d_req_tip(0) <= place_713_top;
  tc_tmp_d_27_d_id_d_1_d_cast_d_ack_tip(0) <= place_150_top;
  tc_tmp_d_27_d_id_d_1_d_cast_d_req_tip(0) <= place_151_top;
  tc_tmp_d_27_d_id_d_2_d_cast_d_ack_tip(0) <= place_156_top;
  tc_tmp_d_27_d_id_d_2_d_cast_d_req_tip(0) <= place_157_top;
  tc_tmp_d_74_d_id_d_1_d_cast_d_ack_tip(0) <= place_284_top;
  tc_tmp_d_74_d_id_d_1_d_cast_d_req_tip(0) <= place_285_top;
  tc_tmp_d_97_d_id_d_1_d_cast_d_ack_tip(0) <= place_362_top;
  tc_tmp_d_97_d_id_d_1_d_cast_d_req_tip(0) <= place_363_top;
  then_d_0_d_entry_tip(0) <= place_24_top;
  then_d_0_to_no_exit_d_4_src_tip(0) <= place_265_top;
  then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_tip(0) <= place_265_top;
  then_d_1_d_entry_tip(0) <= place_52_top;
  then_d_1_to_loopexit_d_10_src_tip(0) <= place_514_top;
  then_d_1_to_no_exit_d_10_d_backedge_src_tip(0) <= place_514_top;
  then_d_2_d_entry_tip(0) <= place_59_top;
  then_d_2_to_loopexit_d_10_src_tip(0) <= place_572_top;
  then_d_2_to_no_exit_d_10_d_backedge_src_tip(0) <= place_572_top;

  cbr_10_oper_tmp_d_42_bool_d_req_ge <= '1';
  op(59) <= cbr_10_oper_tmp_d_42_bool_d_req_top;
  cbr_11_oper_tmp_d_54_bool_d_req_ge <= '1';
  op(74) <= cbr_11_oper_tmp_d_54_bool_d_req_top;
  cbr_12_oper_tmp_d_4223_bool_d_req_ge <= '1';
  op(78) <= cbr_12_oper_tmp_d_4223_bool_d_req_top;
  cbr_13_oper_exitcond128_bool_d_req_ge <= '1';
  op(96) <= cbr_13_oper_exitcond128_bool_d_req_top;
  cbr_14_oper_exitcond131_bool_d_req_ge <= '1';
  op(100) <= cbr_14_oper_exitcond131_bool_d_req_top;
  cbr_15_oper_tmp_d_92_bool_d_req_ge <= '1';
  op(118) <= cbr_15_oper_tmp_d_92_bool_d_req_top;
  cbr_16_oper_tmp_d_11348_bool_d_req_ge <= '1';
  op(130) <= cbr_16_oper_tmp_d_11348_bool_d_req_top;
  cbr_17_oper_tmp_d_113_bool_d_req_ge <= '1';
  op(152) <= cbr_17_oper_tmp_d_113_bool_d_req_top;
  cbr_18_oper_exitcond142_bool_d_req_ge <= '1';
  op(154) <= cbr_18_oper_exitcond142_bool_d_req_top;
  cbr_19_oper_tmp_d_149_bool_d_req_ge <= '1';
  op(161) <= cbr_19_oper_tmp_d_149_bool_d_req_top;
  cbr_20_oper_tmp_d_14574_bool_d_req_ge <= '1';
  op(179) <= cbr_20_oper_tmp_d_14574_bool_d_req_top;
  cbr_21_oper_tmp_d_166_bool_d_req_ge <= '1';
  op(189) <= cbr_21_oper_tmp_d_166_bool_d_req_top;
  cbr_22_oper_tmp_d_14578_bool_d_req_ge <= '1';
  op(203) <= cbr_22_oper_tmp_d_14578_bool_d_req_top;
  cbr_23_oper_tmp_d_14580_bool_d_req_ge <= '1';
  op(217) <= cbr_23_oper_tmp_d_14580_bool_d_req_top;
  cbr_24_oper_exitcond145_bool_d_req_ge <= '1';
  op(220) <= cbr_24_oper_exitcond145_bool_d_req_top;
  cbr_25_oper_tmp_d_202_bool_d_req_ge <= '1';
  op(227) <= cbr_25_oper_tmp_d_202_bool_d_req_top;
  cbr_26_oper_tmp_d_20299_bool_d_req_ge <= '1';
  op(242) <= cbr_26_oper_tmp_d_20299_bool_d_req_top;
  cbr_27_oper_exitcond150_bool_d_req_ge <= '1';
  op(248) <= cbr_27_oper_exitcond150_bool_d_req_top;
  cbr_28_oper_tmp_d_221_bool_d_req_ge <= '1';
  op(255) <= cbr_28_oper_tmp_d_221_bool_d_req_top;
  cbr_29_oper_tmp_d_221111_bool_d_req_ge <= '1';
  op(272) <= cbr_29_oper_tmp_d_221111_bool_d_req_top;
  cbr_30_oper_exitcond158_bool_d_req_ge <= '1';
  op(278) <= cbr_30_oper_exitcond158_bool_d_req_top;
  cbr_6_oper_exitcond_bool_d_req_ge <= '1';
  op(18) <= cbr_6_oper_exitcond_bool_d_req_top;
  cbr_7_oper_exitcond120_bool_d_req_ge <= '1';
  op(21) <= cbr_7_oper_exitcond120_bool_d_req_top;
  cbr_8_oper_tmp_d_16_bool_d_req_ge <= '1';
  op(23) <= cbr_8_oper_tmp_d_16_bool_d_req_top;
  cbr_9_oper_tmp_d_1614_bool_d_req_ge <= '1';
  op(42) <= cbr_9_oper_tmp_d_1614_bool_d_req_top;
  else_d_0_d_entry_ge <= '1';
  else_d_0_to_else_d_1_src_ge <= ip(185);
  else_d_0_to_then_d_2_src_ge <= ip(184);
  else_d_1_d_entry_ge <= '1';
  else_d_1_to_loopexit_d_10_src_ge <= ip(215);
  else_d_1_to_no_exit_d_10_d_backedge_src_ge <= ip(214);
  fin_ge <= '1';
  op(1) <= fin_top;
  indvar118_d_ph_d_ph_mux_1_d_ack_ge <= ip(8);
  indvar118_d_ph_d_ph_mux_1_d_req0_ge <= '1';
  op(9) <= indvar118_d_ph_d_ph_mux_1_d_req0_top;
  indvar118_d_ph_d_ph_mux_1_d_req1_ge <= '1';
  op(8) <= indvar118_d_ph_d_ph_mux_1_d_req1_top;
  indvar121_mux_1_d_ack_ge <= ip(25);
  indvar121_mux_1_d_req0_ge <= '1';
  op(25) <= indvar121_mux_1_d_req0_top;
  indvar121_mux_1_d_req1_ge <= '1';
  op(24) <= indvar121_mux_1_d_req1_top;
  indvar123_mux_1_d_ack_ge <= ip(60);
  indvar123_mux_1_d_req0_ge <= '1';
  op(64) <= indvar123_mux_1_d_req0_top;
  indvar123_mux_1_d_req1_ge <= '1';
  op(63) <= indvar123_mux_1_d_req1_top;
  indvar126_mux_1_d_ack_ge <= ip(77);
  indvar126_mux_1_d_req0_ge <= '1';
  op(82) <= indvar126_mux_1_d_req0_top;
  indvar126_mux_1_d_req1_ge <= '1';
  op(81) <= indvar126_mux_1_d_req1_top;
  indvar129_mux_1_d_ack_ge <= ip(44);
  indvar129_mux_1_d_req0_ge <= '1';
  op(44) <= indvar129_mux_1_d_req0_top;
  indvar129_mux_1_d_req1_ge <= '1';
  op(43) <= indvar129_mux_1_d_req1_top;
  indvar132_mux_1_d_ack_ge <= ip(128);
  indvar132_mux_1_d_req0_ge <= '1';
  op(133) <= indvar132_mux_1_d_req0_top;
  indvar132_mux_1_d_req1_ge <= '1';
  op(132) <= indvar132_mux_1_d_req1_top;
  indvar134_mux_1_d_ack_ge <= ip(98);
  indvar134_mux_1_d_req0_ge <= '1';
  op(102) <= indvar134_mux_1_d_req0_top;
  indvar134_mux_1_d_req1_ge <= '1';
  op(101) <= indvar134_mux_1_d_req1_top;
  indvar138_mux_1_d_ack_ge <= ip(107);
  indvar138_mux_1_d_req0_ge <= '1';
  op(113) <= indvar138_mux_1_d_req0_top;
  indvar138_mux_1_d_req1_ge <= '1';
  op(112) <= indvar138_mux_1_d_req1_top;
  indvar143_mux_1_d_ack_ge <= ip(152);
  indvar143_mux_1_d_req0_ge <= '1';
  op(156) <= indvar143_mux_1_d_req0_top;
  indvar143_mux_1_d_req1_ge <= '1';
  op(155) <= indvar143_mux_1_d_req1_top;
  indvar146_mux_1_d_ack_ge <= ip(226);
  indvar146_mux_1_d_req0_ge <= '1';
  op(229) <= indvar146_mux_1_d_req0_top;
  indvar146_mux_1_d_req1_ge <= '1';
  op(228) <= indvar146_mux_1_d_req1_top;
  indvar148_mux_1_d_ack_ge <= ip(220);
  indvar148_mux_1_d_req0_ge <= '1';
  op(222) <= indvar148_mux_1_d_req0_top;
  indvar148_mux_1_d_req1_ge <= '1';
  op(221) <= indvar148_mux_1_d_req1_top;
  indvar151_mux_1_d_ack_ge <= ip(253);
  indvar151_mux_1_d_req0_ge <= '1';
  op(257) <= indvar151_mux_1_d_req0_top;
  indvar151_mux_1_d_req1_ge <= '1';
  op(256) <= indvar151_mux_1_d_req1_top;
  indvar153_mux_1_d_ack_ge <= ip(247);
  indvar153_mux_1_d_req0_ge <= '1';
  op(250) <= indvar153_mux_1_d_req0_top;
  indvar153_mux_1_d_req1_ge <= '1';
  op(249) <= indvar153_mux_1_d_req1_top;
  indvar_mux_1_d_ack_ge <= ip(9);
  indvar_mux_1_d_req0_ge <= '1';
  op(11) <= indvar_mux_1_d_req0_top;
  indvar_mux_1_d_req1_ge <= '1';
  op(10) <= indvar_mux_1_d_req1_top;
  init_ge <= ip(1);
  j_d_3_d_in_d_ph_mux_1_d_ack_ge <= ip(45);
  j_d_3_d_in_d_ph_mux_1_d_req0_ge <= '1';
  op(46) <= j_d_3_d_in_d_ph_mux_1_d_req0_top;
  j_d_3_d_in_d_ph_mux_1_d_req1_ge <= '1';
  op(45) <= j_d_3_d_in_d_ph_mux_1_d_req1_top;
  j_d_3_d_in_mux_1_d_ack_ge <= ip(51);
  j_d_3_d_in_mux_1_d_req0_ge <= '1';
  op(54) <= j_d_3_d_in_mux_1_d_req0_top;
  j_d_3_d_in_mux_1_d_req1_ge <= '1';
  op(53) <= j_d_3_d_in_mux_1_d_req1_top;
  j_d_9_d_2_d_be_mux_1_d_ack_ge <= ip(178);
  j_d_9_d_2_d_be_mux_1_d_req0_ge <= '1';
  op(183) <= j_d_9_d_2_d_be_mux_1_d_req0_top;
  j_d_9_d_2_d_be_mux_1_d_req1_ge <= '1';
  op(182) <= j_d_9_d_2_d_be_mux_1_d_req1_top;
  j_d_9_d_2_d_be_mux_2_d_ack_ge <= ip(177);
  j_d_9_d_2_d_be_mux_2_d_req0_ge <= '1';
  op(181) <= j_d_9_d_2_d_be_mux_2_d_req0_top;
  j_d_9_d_2_d_be_mux_2_d_req1_ge <= '1';
  op(180) <= j_d_9_d_2_d_be_mux_2_d_req1_top;
  j_d_9_d_2_mux_1_d_ack_ge <= ip(154);
  j_d_9_d_2_mux_1_d_req0_ge <= '1';
  op(159) <= j_d_9_d_2_mux_1_d_req0_top;
  j_d_9_d_2_mux_1_d_req1_ge <= '1';
  op(158) <= j_d_9_d_2_mux_1_d_req1_top;
  k_d_1_d_in_d_ph_mux_1_d_ack_ge <= ip(99);
  k_d_1_d_in_d_ph_mux_1_d_req0_ge <= '1';
  op(104) <= k_d_1_d_in_d_ph_mux_1_d_req0_top;
  k_d_1_d_in_d_ph_mux_1_d_req1_ge <= '1';
  op(103) <= k_d_1_d_in_d_ph_mux_1_d_req1_top;
  k_d_2_d_3_mux_1_d_ack_ge <= ip(242);
  k_d_2_d_3_mux_1_d_req0_ge <= '1';
  op(245) <= k_d_2_d_3_mux_1_d_req0_top;
  k_d_2_d_3_mux_1_d_req1_ge <= '1';
  op(244) <= k_d_2_d_3_mux_1_d_req1_top;
  k_d_3_d_0_mux_1_d_ack_ge <= ip(221);
  k_d_3_d_0_mux_1_d_req0_ge <= '1';
  op(224) <= k_d_3_d_0_mux_1_d_req0_top;
  k_d_3_d_0_mux_1_d_req1_ge <= '1';
  op(223) <= k_d_3_d_0_mux_1_d_req1_top;
  k_d_4_d_3_mux_1_d_ack_ge <= ip(271);
  k_d_4_d_3_mux_1_d_req0_ge <= '1';
  op(275) <= k_d_4_d_3_mux_1_d_req0_top;
  k_d_4_d_3_mux_1_d_req1_ge <= '1';
  op(274) <= k_d_4_d_3_mux_1_d_req1_top;
  k_d_5_d_0_mux_1_d_ack_ge <= ip(248);
  k_d_5_d_0_mux_1_d_req0_ge <= '1';
  op(252) <= k_d_5_d_0_mux_1_d_req0_top;
  k_d_5_d_0_mux_1_d_req1_ge <= '1';
  op(251) <= k_d_5_d_0_mux_1_d_req1_top;
  load_A_d_ack_ge <= ip(3);
  load_A_d_req_ge <= '1';
  op(3) <= load_A_d_req_top;
  load_ccoeff_d_ack_ge <= ip(5);
  load_ccoeff_d_req_ge <= '1';
  op(5) <= load_ccoeff_d_req_top;
  load_l_array_d_ack_ge <= ip(6);
  load_l_array_d_req_ge <= '1';
  op(6) <= load_l_array_d_req_top;
  load_noofelem_d_ack_ge <= ip(2);
  load_noofelem_d_req_ge <= '1';
  op(2) <= load_noofelem_d_req_top;
  load_rcoeff_d_ack_ge <= ip(4);
  load_rcoeff_d_req_ge <= '1';
  op(4) <= load_rcoeff_d_req_top;
  load_start_call_divide_0_return_d_ack_ge <= ip(123);
  load_start_call_divide_0_return_d_req_ge <= '1';
  op(128) <= load_start_call_divide_0_return_d_req_top;
  load_tmp_d_103_d_ack_ge <= ip(118);
  load_tmp_d_103_d_req_ge <= '1';
  op(123) <= load_tmp_d_103_d_req_top;
  load_tmp_d_108_d_ack_ge <= ip(119);
  load_tmp_d_108_d_req_ge <= '1';
  op(124) <= load_tmp_d_108_d_req_top;
  load_tmp_d_123_d_ack_ge <= ip(135);
  load_tmp_d_123_d_req_ge <= '1';
  op(140) <= load_tmp_d_123_d_req_top;
  load_tmp_d_128_d_ack_ge <= ip(136);
  load_tmp_d_128_d_req_ge <= '1';
  op(141) <= load_tmp_d_128_d_req_top;
  load_tmp_d_133_d_ack_ge <= ip(140);
  load_tmp_d_133_d_req_ge <= '1';
  op(145) <= load_tmp_d_133_d_req_top;
  load_tmp_d_159_d_ack_ge <= ip(166);
  load_tmp_d_159_d_req_ge <= '1';
  op(170) <= load_tmp_d_159_d_req_top;
  load_tmp_d_180_d_ack_ge <= ip(195);
  load_tmp_d_180_d_req_ge <= '1';
  op(199) <= load_tmp_d_180_d_req_top;
  load_tmp_d_193_d_ack_ge <= ip(210);
  load_tmp_d_193_d_req_ge <= '1';
  op(213) <= load_tmp_d_193_d_req_top;
  load_tmp_d_211_d_ack_ge <= ip(234);
  load_tmp_d_211_d_req_ge <= '1';
  op(237) <= load_tmp_d_211_d_req_top;
  load_tmp_d_21_d_ack_ge <= ip(28);
  load_tmp_d_21_d_req_ge <= '1';
  op(28) <= load_tmp_d_21_d_req_top;
  load_tmp_d_230_d_ack_ge <= ip(263);
  load_tmp_d_230_d_req_ge <= '1';
  op(267) <= load_tmp_d_230_d_req_top;
  load_tmp_d_26_d_ack_ge <= ip(30);
  load_tmp_d_26_d_req_ge <= '1';
  op(30) <= load_tmp_d_26_d_req_top;
  load_tmp_d_31_d_ack_ge <= ip(37);
  load_tmp_d_31_d_req_ge <= '1';
  op(37) <= load_tmp_d_31_d_req_top;
  load_tmp_d_48_d_ack_ge <= ip(67);
  load_tmp_d_48_d_req_ge <= '1';
  op(72) <= load_tmp_d_48_d_req_top;
  load_tmp_d_53_d_ack_ge <= ip(58);
  load_tmp_d_53_d_req_ge <= '1';
  op(61) <= load_tmp_d_53_d_req_top;
  load_tmp_d_66_d_ack_ge <= ip(81);
  load_tmp_d_66_d_req_ge <= '1';
  op(86) <= load_tmp_d_66_d_req_top;
  load_tmp_d_75_d_ack_ge <= ip(86);
  load_tmp_d_75_d_req_ge <= '1';
  op(91) <= load_tmp_d_75_d_req_top;
  load_u_array_d_ack_ge <= ip(7);
  load_u_array_d_req_ge <= '1';
  op(7) <= load_u_array_d_req_top;
  loopentry_d_12_d_entry_ge <= '1';
  loopentry_d_12_d_loopexit_to_loopentry_d_12_src_ge <= '1';
  loopentry_d_12_d_pre_ge <= '1';
  loopentry_d_12_to_loopexit_d_12_src_ge <= ip(224);
  loopentry_d_12_to_no_exit_d_12_d_preheader_src_ge <= ip(225);
  loopentry_d_14_d_entry_ge <= '1';
  loopentry_d_14_d_loopexit_to_loopentry_d_14_src_ge <= '1';
  loopentry_d_14_d_pre_ge <= '1';
  loopentry_d_14_to_loopexit_d_14_src_ge <= ip(252);
  loopentry_d_14_to_no_exit_d_14_d_preheader_src_ge <= ip(251);
  loopentry_d_2_to_loopentry_d_4_d_outer_d_preheader_src_ge <= ip(24);
  loopentry_d_2_to_no_exit_d_2_d_preheader_src_ge <= ip(23);
  loopentry_d_4_d_entry_ge <= '1';
  loopentry_d_4_d_loopexit_to_loopentry_d_4_src_ge <= '1';
  loopentry_d_4_d_outer_d_entry_ge <= '1';
  loopentry_d_4_d_outer_d_pre_ge <= '1';
  loopentry_d_4_d_outer_d_preheader_to_loopentry_d_4_d_outer_src_ge <= '1';
  loopentry_d_4_d_outer_to_loopentry_d_4_src_ge <= '1';
  loopentry_d_4_d_pre_ge <= '1';
  loopentry_d_4_to_no_exit_d_4_d_preheader_src_ge <= ip(55);
  loopentry_d_4_to_no_exit_d_5_d_preheader_src_ge <= ip(56);
  loopentry_d_7_d_outer_d_entry_ge <= '1';
  loopentry_d_7_d_outer_d_loopexit_to_loopentry_d_7_d_outer_src_ge <= '1';
  loopentry_d_7_d_outer_d_pre_ge <= '1';
  loopentry_d_7_d_outer_to_loopentry_d_7_src_ge <= '1';
  loopentry_d_7_to_loopexit_d_7_src_ge <= ip(113);
  loopentry_d_7_to_no_exit_d_7_src_ge <= ip(112);
  loopexit_d_10_to_loopentry_d_12_d_loopexit_src_ge <= ip(218);
  loopexit_d_10_to_no_exit_d_10_d_outer_src_ge <= ip(219);
  loopexit_d_12_d_entry_ge <= '1';
  loopexit_d_12_to_loopentry_d_12_src_ge <= ip(246);
  loopexit_d_12_to_loopentry_d_14_d_loopexit_src_ge <= ip(245);
  loopexit_d_14_d_entry_ge <= '1';
  loopexit_d_14_to_loopentry_d_14_src_ge <= ip(275);
  loopexit_d_14_to_return_src_ge <= ip(274);
  loopexit_d_1_to_loopentry_d_2_src_ge <= ip(20);
  loopexit_d_1_to_no_exit_d_1_d_outer_src_ge <= ip(21);
  loopexit_d_5_d_entry_ge <= '1';
  loopexit_d_5_to_loopentry_d_4_d_outer_src_ge <= ip(97);
  loopexit_d_5_to_loopentry_d_7_d_outer_d_loopexit_src_ge <= ip(96);
  loopexit_d_7_to_loopentry_d_7_d_outer_src_ge <= ip(151);
  loopexit_d_7_to_no_exit_d_10_d_outer_d_loopexit_src_ge <= ip(150);
  maxcoeff_d_2_d_2_mux_1_d_ack_ge <= ip(61);
  maxcoeff_d_2_d_2_mux_1_d_req0_ge <= '1';
  op(66) <= maxcoeff_d_2_d_2_mux_1_d_req0_top;
  maxcoeff_d_2_d_2_mux_1_d_req1_ge <= '1';
  op(65) <= maxcoeff_d_2_d_2_mux_1_d_req1_top;
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_ack_ge <= ip(76);
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_ge <= '1';
  op(80) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req0_top;
  maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_ge <= '1';
  op(79) <= maxcoeff_d_2_d_3_d_ph_d_ph_d_ph_mux_1_d_req1_top;
  maxcoeff_d_2_d_ph_mux_1_d_ack_ge <= ip(46);
  maxcoeff_d_2_d_ph_mux_1_d_req0_ge <= '1';
  op(48) <= maxcoeff_d_2_d_ph_mux_1_d_req0_top;
  maxcoeff_d_2_d_ph_mux_1_d_req1_ge <= '1';
  op(47) <= maxcoeff_d_2_d_ph_mux_1_d_req1_top;
  maxcoeff_d_2_mux_1_d_ack_ge <= ip(52);
  maxcoeff_d_2_mux_1_d_req0_ge <= '1';
  op(56) <= maxcoeff_d_2_mux_1_d_req0_top;
  maxcoeff_d_2_mux_1_d_req1_ge <= '1';
  op(55) <= maxcoeff_d_2_mux_1_d_req1_top;
  no_exit_d_10_to_else_d_0_src_ge <= ip(157);
  no_exit_d_10_to_then_d_1_src_ge <= ip(156);
  no_exit_d_12_d_entry_ge <= '1';
  no_exit_d_12_to_loopexit_d_12_d_loopexit_src_ge <= ip(239);
  no_exit_d_12_to_no_exit_d_12_src_ge <= ip(240);
  no_exit_d_14_d_entry_ge <= '1';
  no_exit_d_14_to_loopexit_d_14_d_loopexit_src_ge <= ip(269);
  no_exit_d_14_to_no_exit_d_14_src_ge <= ip(268);
  no_exit_d_1_d_entry_ge <= '1';
  no_exit_d_1_to_loopexit_d_1_src_ge <= ip(16);
  no_exit_d_1_to_no_exit_d_1_src_ge <= ip(17);
  no_exit_d_2_d_entry_ge <= '1';
  no_exit_d_2_to_loopentry_d_4_d_outer_d_loopexit_src_ge <= ip(43);
  no_exit_d_2_to_no_exit_d_2_src_ge <= ip(42);
  no_exit_d_4_d_entry_ge <= '1';
  no_exit_d_4_d_pre_ge <= '1';
  no_exit_d_4_d_preheader_d_entry_ge <= '1';
  no_exit_d_4_d_preheader_to_no_exit_d_4_src_ge <= '1';
  no_exit_d_4_to_loopentry_d_4_d_loopexit_src_ge <= ip(70);
  no_exit_d_4_to_then_d_0_src_ge <= ip(69);
  no_exit_d_5_d_entry_ge <= '1';
  no_exit_d_5_to_loopexit_d_5_src_ge <= ip(91);
  no_exit_d_5_to_no_exit_d_5_src_ge <= ip(92);
  no_exit_d_7_d_entry_ge <= '1';
  no_exit_d_7_to_loopentry_d_7_d_backedge_src_ge <= ip(126);
  no_exit_d_7_to_no_exit_d_8_d_preheader_src_ge <= ip(125);
  no_exit_d_8_d_entry_ge <= '1';
  no_exit_d_8_to_loopentry_d_7_d_backedge_d_loopexit_src_ge <= ip(148);
  no_exit_d_8_to_no_exit_d_8_src_ge <= ip(147);
  oper_exitcond120_bool_d_ack_ge <= ip(19);
  oper_exitcond120_bool_d_req_ge <= '1';
  op(20) <= oper_exitcond120_bool_d_req_top;
  oper_exitcond128_bool_d_ack_ge <= ip(90);
  oper_exitcond128_bool_d_req_ge <= '1';
  op(95) <= oper_exitcond128_bool_d_req_top;
  oper_exitcond131_bool_d_ack_ge <= ip(95);
  oper_exitcond131_bool_d_req_ge <= '1';
  op(99) <= oper_exitcond131_bool_d_req_top;
  oper_exitcond142_bool_d_ack_ge <= ip(149);
  oper_exitcond142_bool_d_req_ge <= '1';
  op(153) <= oper_exitcond142_bool_d_req_top;
  oper_exitcond145_bool_d_ack_ge <= ip(217);
  oper_exitcond145_bool_d_req_ge <= '1';
  op(219) <= oper_exitcond145_bool_d_req_top;
  oper_exitcond150_bool_d_ack_ge <= ip(244);
  oper_exitcond150_bool_d_req_ge <= '1';
  op(247) <= oper_exitcond150_bool_d_req_top;
  oper_exitcond158_bool_d_ack_ge <= ip(273);
  oper_exitcond158_bool_d_req_ge <= '1';
  op(277) <= oper_exitcond158_bool_d_req_top;
  oper_exitcond_bool_d_ack_ge <= ip(15);
  oper_exitcond_bool_d_req_ge <= '1';
  op(17) <= oper_exitcond_bool_d_req_top;
  oper_inc_d_11_int_d_ack_ge <= ip(241);
  oper_inc_d_11_int_d_req_ge <= '1';
  op(243) <= oper_inc_d_11_int_d_req_top;
  oper_inc_d_12_int_d_ack_ge <= ip(236);
  oper_inc_d_12_int_d_req_ge <= '1';
  op(239) <= oper_inc_d_12_int_d_req_top;
  oper_inc_d_14_int_d_ack_ge <= ip(270);
  oper_inc_d_14_int_d_req_ge <= '1';
  op(273) <= oper_inc_d_14_int_d_req_top;
  oper_inc_d_15_int_d_ack_ge <= ip(265);
  oper_inc_d_15_int_d_req_ge <= '1';
  op(269) <= oper_inc_d_15_int_d_req_top;
  oper_inc_d_2_int_d_ack_ge <= ip(39);
  oper_inc_d_2_int_d_req_ge <= '1';
  op(39) <= oper_inc_d_2_int_d_req_top;
  oper_inc_d_5_int_d_ack_ge <= ip(93);
  oper_inc_d_5_int_d_req_ge <= '1';
  op(97) <= oper_inc_d_5_int_d_req_top;
  oper_inc_d_960_int_d_ack_ge <= ip(173);
  oper_inc_d_960_int_d_req_ge <= '1';
  op(177) <= oper_inc_d_960_int_d_req_top;
  oper_inc_d_976_int_d_ack_ge <= ip(197);
  oper_inc_d_976_int_d_req_ge <= '1';
  op(201) <= oper_inc_d_976_int_d_req_top;
  oper_inc_d_9_int_d_ack_ge <= ip(212);
  oper_inc_d_9_int_d_req_ge <= '1';
  op(215) <= oper_inc_d_9_int_d_req_top;
  oper_indvar_d_next119_uint_d_ack_ge <= ip(18);
  oper_indvar_d_next119_uint_d_req_ge <= '1';
  op(19) <= oper_indvar_d_next119_uint_d_req_top;
  oper_indvar_d_next122_uint_d_ack_ge <= ip(41);
  oper_indvar_d_next122_uint_d_req_ge <= '1';
  op(41) <= oper_indvar_d_next122_uint_d_req_top;
  oper_indvar_d_next124_uint_d_ack_ge <= ip(73);
  oper_indvar_d_next124_uint_d_req_ge <= '1';
  op(77) <= oper_indvar_d_next124_uint_d_req_top;
  oper_indvar_d_next127_uint_d_ack_ge <= ip(89);
  oper_indvar_d_next127_uint_d_req_ge <= '1';
  op(94) <= oper_indvar_d_next127_uint_d_req_top;
  oper_indvar_d_next130_uint_d_ack_ge <= ip(94);
  oper_indvar_d_next130_uint_d_req_ge <= '1';
  op(98) <= oper_indvar_d_next130_uint_d_req_top;
  oper_indvar_d_next133_uint_d_ack_ge <= ip(146);
  oper_indvar_d_next133_uint_d_req_ge <= '1';
  op(151) <= oper_indvar_d_next133_uint_d_req_top;
  oper_indvar_d_next139_uint_d_ack_ge <= ip(127);
  oper_indvar_d_next139_uint_d_req_ge <= '1';
  op(131) <= oper_indvar_d_next139_uint_d_req_top;
  oper_indvar_d_next144_uint_d_ack_ge <= ip(216);
  oper_indvar_d_next144_uint_d_req_ge <= '1';
  op(218) <= oper_indvar_d_next144_uint_d_req_top;
  oper_indvar_d_next147_uint_d_ack_ge <= ip(238);
  oper_indvar_d_next147_uint_d_req_ge <= '1';
  op(241) <= oper_indvar_d_next147_uint_d_req_top;
  oper_indvar_d_next149_uint_d_ack_ge <= ip(243);
  oper_indvar_d_next149_uint_d_req_ge <= '1';
  op(246) <= oper_indvar_d_next149_uint_d_req_top;
  oper_indvar_d_next152_uint_d_ack_ge <= ip(267);
  oper_indvar_d_next152_uint_d_req_ge <= '1';
  op(271) <= oper_indvar_d_next152_uint_d_req_top;
  oper_indvar_d_next157_uint_d_ack_ge <= ip(272);
  oper_indvar_d_next157_uint_d_req_ge <= '1';
  op(276) <= oper_indvar_d_next157_uint_d_req_top;
  oper_indvar_d_next_uint_d_ack_ge <= ip(14);
  oper_indvar_d_next_uint_d_req_ge <= '1';
  op(16) <= oper_indvar_d_next_uint_d_req_top;
  oper_j_d_321_int_d_ack_ge <= ip(71);
  oper_j_d_321_int_d_req_ge <= '1';
  op(75) <= oper_j_d_321_int_d_req_top;
  oper_j_d_3_int_d_ack_ge <= ip(53);
  oper_j_d_3_int_d_req_ge <= '1';
  op(57) <= oper_j_d_3_int_d_req_top;
  oper_j_d_746_int_d_ack_ge <= ip(104);
  oper_j_d_746_int_d_req_ge <= '1';
  op(109) <= oper_j_d_746_int_d_req_top;
  oper_j_d_7_int_d_ack_ge <= ip(144);
  oper_j_d_7_int_d_req_ge <= '1';
  op(149) <= oper_j_d_7_int_d_req_top;
  oper_k_d_1_d_in_int_d_ack_ge <= ip(109);
  oper_k_d_1_d_in_int_d_req_ge <= '1';
  op(115) <= oper_k_d_1_d_in_int_d_req_top;
  oper_k_d_1_int_d_ack_ge <= ip(110);
  oper_k_d_1_int_d_req_ge <= '1';
  op(116) <= oper_k_d_1_int_d_req_top;
  oper_k_d_2_d_2_int_d_ack_ge <= ip(228);
  oper_k_d_2_d_2_int_d_req_ge <= '1';
  op(231) <= oper_k_d_2_d_2_int_d_req_top;
  oper_k_d_4_d_2_int_d_ack_ge <= ip(257);
  oper_k_d_4_d_2_int_d_req_ge <= '1';
  op(261) <= oper_k_d_4_d_2_int_d_req_top;
  oper_tmp_d_107_d_id_d_1_uint_d_ack_ge <= ip(101);
  oper_tmp_d_107_d_id_d_1_uint_d_req_ge <= '1';
  op(106) <= oper_tmp_d_107_d_id_d_1_uint_d_req_top;
  oper_tmp_d_107_d_lvl_d_1_uint_d_ack_ge <= ip(102);
  oper_tmp_d_107_d_lvl_d_1_uint_d_req_ge <= '1';
  op(107) <= oper_tmp_d_107_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_107_d_lvl_d_2_uint_d_ack_ge <= ip(103);
  oper_tmp_d_107_d_lvl_d_2_uint_d_req_ge <= '1';
  op(108) <= oper_tmp_d_107_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_11348_bool_d_ack_ge <= ip(105);
  oper_tmp_d_11348_bool_d_req_ge <= '1';
  op(110) <= oper_tmp_d_11348_bool_d_req_top;
  oper_tmp_d_113_bool_d_ack_ge <= ip(145);
  oper_tmp_d_113_bool_d_req_ge <= '1';
  op(150) <= oper_tmp_d_113_bool_d_req_top;
  oper_tmp_d_118_d_id_d_1_uint_d_ack_ge <= ip(132);
  oper_tmp_d_118_d_id_d_1_uint_d_req_ge <= '1';
  op(137) <= oper_tmp_d_118_d_id_d_1_uint_d_req_top;
  oper_tmp_d_118_d_lvl_d_1_uint_d_ack_ge <= ip(133);
  oper_tmp_d_118_d_lvl_d_1_uint_d_req_ge <= '1';
  op(138) <= oper_tmp_d_118_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_118_d_lvl_d_2_uint_d_ack_ge <= ip(134);
  oper_tmp_d_118_d_lvl_d_2_uint_d_req_ge <= '1';
  op(139) <= oper_tmp_d_118_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_11_d_id_d_1_uint_d_ack_ge <= ip(10);
  oper_tmp_d_11_d_id_d_1_uint_d_req_ge <= '1';
  op(12) <= oper_tmp_d_11_d_id_d_1_uint_d_req_top;
  oper_tmp_d_11_d_lvl_d_1_uint_d_ack_ge <= ip(11);
  oper_tmp_d_11_d_lvl_d_1_uint_d_req_ge <= '1';
  op(13) <= oper_tmp_d_11_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_11_d_lvl_d_2_uint_d_ack_ge <= ip(12);
  oper_tmp_d_11_d_lvl_d_2_uint_d_req_ge <= '1';
  op(14) <= oper_tmp_d_11_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_125_uint_d_ack_ge <= ip(62);
  oper_tmp_d_125_uint_d_req_ge <= '1';
  op(67) <= oper_tmp_d_125_uint_d_req_top;
  oper_tmp_d_132_d_id_d_1_uint_d_ack_ge <= ip(137);
  oper_tmp_d_132_d_id_d_1_uint_d_req_ge <= '1';
  op(142) <= oper_tmp_d_132_d_id_d_1_uint_d_req_top;
  oper_tmp_d_132_d_lvl_d_1_uint_d_ack_ge <= ip(138);
  oper_tmp_d_132_d_lvl_d_1_uint_d_req_ge <= '1';
  op(143) <= oper_tmp_d_132_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_132_d_lvl_d_2_uint_d_ack_ge <= ip(139);
  oper_tmp_d_132_d_lvl_d_2_uint_d_req_ge <= '1';
  op(144) <= oper_tmp_d_132_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_134_float_d_ack_ge <= ip(141);
  oper_tmp_d_134_float_d_req_ge <= '1';
  op(146) <= oper_tmp_d_134_float_d_req_top;
  oper_tmp_d_135_float_d_ack_ge <= ip(142);
  oper_tmp_d_135_float_d_req_ge <= '1';
  op(147) <= oper_tmp_d_135_float_d_req_top;
  oper_tmp_d_136_uint_d_ack_ge <= ip(106);
  oper_tmp_d_136_uint_d_req_ge <= '1';
  op(111) <= oper_tmp_d_136_uint_d_req_top;
  oper_tmp_d_137_uint_d_ack_ge <= ip(129);
  oper_tmp_d_137_uint_d_req_ge <= '1';
  op(134) <= oper_tmp_d_137_uint_d_req_top;
  oper_tmp_d_14574_bool_d_ack_ge <= ip(174);
  oper_tmp_d_14574_bool_d_req_ge <= '1';
  op(178) <= oper_tmp_d_14574_bool_d_req_top;
  oper_tmp_d_14578_bool_d_ack_ge <= ip(198);
  oper_tmp_d_14578_bool_d_req_ge <= '1';
  op(202) <= oper_tmp_d_14578_bool_d_req_top;
  oper_tmp_d_14580_bool_d_ack_ge <= ip(213);
  oper_tmp_d_14580_bool_d_req_ge <= '1';
  op(216) <= oper_tmp_d_14580_bool_d_req_top;
  oper_tmp_d_149_bool_d_ack_ge <= ip(155);
  oper_tmp_d_149_bool_d_req_ge <= '1';
  op(160) <= oper_tmp_d_149_bool_d_req_top;
  oper_tmp_d_154_d_id_d_1_uint_d_ack_ge <= ip(158);
  oper_tmp_d_154_d_id_d_1_uint_d_req_ge <= '1';
  op(162) <= oper_tmp_d_154_d_id_d_1_uint_d_req_top;
  oper_tmp_d_154_d_lvl_d_1_uint_d_ack_ge <= ip(159);
  oper_tmp_d_154_d_lvl_d_1_uint_d_req_ge <= '1';
  op(163) <= oper_tmp_d_154_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_154_d_lvl_d_2_uint_d_ack_ge <= ip(161);
  oper_tmp_d_154_d_lvl_d_2_uint_d_req_ge <= '1';
  op(165) <= oper_tmp_d_154_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_155_uint_d_ack_ge <= ip(255);
  oper_tmp_d_155_uint_d_req_ge <= '1';
  op(259) <= oper_tmp_d_155_uint_d_req_top;
  oper_tmp_d_158_d_id_d_1_uint_d_ack_ge <= ip(162);
  oper_tmp_d_158_d_id_d_1_uint_d_req_ge <= '1';
  op(166) <= oper_tmp_d_158_d_id_d_1_uint_d_req_top;
  oper_tmp_d_158_d_lvl_d_1_uint_d_ack_ge <= ip(163);
  oper_tmp_d_158_d_lvl_d_1_uint_d_req_ge <= '1';
  op(167) <= oper_tmp_d_158_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_158_d_lvl_d_2_uint_d_ack_ge <= ip(165);
  oper_tmp_d_158_d_lvl_d_2_uint_d_req_ge <= '1';
  op(169) <= oper_tmp_d_158_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_1614_bool_d_ack_ge <= ip(40);
  oper_tmp_d_1614_bool_d_req_ge <= '1';
  op(40) <= oper_tmp_d_1614_bool_d_req_top;
  oper_tmp_d_163_d_id_d_1_uint_d_ack_ge <= ip(168);
  oper_tmp_d_163_d_id_d_1_uint_d_req_ge <= '1';
  op(172) <= oper_tmp_d_163_d_id_d_1_uint_d_req_top;
  oper_tmp_d_163_d_lvl_d_1_uint_d_ack_ge <= ip(169);
  oper_tmp_d_163_d_lvl_d_1_uint_d_req_ge <= '1';
  op(173) <= oper_tmp_d_163_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_163_d_lvl_d_2_uint_d_ack_ge <= ip(171);
  oper_tmp_d_163_d_lvl_d_2_uint_d_req_ge <= '1';
  op(175) <= oper_tmp_d_163_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_166_bool_d_ack_ge <= ip(179);
  oper_tmp_d_166_bool_d_req_ge <= '1';
  op(184) <= oper_tmp_d_166_bool_d_req_top;
  oper_tmp_d_16_bool_d_ack_ge <= ip(22);
  oper_tmp_d_16_bool_d_req_ge <= '1';
  op(22) <= oper_tmp_d_16_bool_d_req_top;
  oper_tmp_d_171_d_id_d_1_uint_d_ack_ge <= ip(180);
  oper_tmp_d_171_d_id_d_1_uint_d_req_ge <= '1';
  op(185) <= oper_tmp_d_171_d_id_d_1_uint_d_req_top;
  oper_tmp_d_171_d_lvl_d_1_uint_d_ack_ge <= ip(181);
  oper_tmp_d_171_d_lvl_d_1_uint_d_req_ge <= '1';
  op(186) <= oper_tmp_d_171_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_171_d_lvl_d_2_uint_d_ack_ge <= ip(183);
  oper_tmp_d_171_d_lvl_d_2_uint_d_req_ge <= '1';
  op(188) <= oper_tmp_d_171_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_175_d_id_d_1_uint_d_ack_ge <= ip(187);
  oper_tmp_d_175_d_id_d_1_uint_d_req_ge <= '1';
  op(191) <= oper_tmp_d_175_d_id_d_1_uint_d_req_top;
  oper_tmp_d_175_d_lvl_d_1_uint_d_ack_ge <= ip(188);
  oper_tmp_d_175_d_lvl_d_1_uint_d_req_ge <= '1';
  op(192) <= oper_tmp_d_175_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_175_d_lvl_d_2_uint_d_ack_ge <= ip(190);
  oper_tmp_d_175_d_lvl_d_2_uint_d_req_ge <= '1';
  op(194) <= oper_tmp_d_175_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_179_d_id_d_1_uint_d_ack_ge <= ip(191);
  oper_tmp_d_179_d_id_d_1_uint_d_req_ge <= '1';
  op(195) <= oper_tmp_d_179_d_id_d_1_uint_d_req_top;
  oper_tmp_d_179_d_lvl_d_1_uint_d_ack_ge <= ip(192);
  oper_tmp_d_179_d_lvl_d_1_uint_d_req_ge <= '1';
  op(196) <= oper_tmp_d_179_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_179_d_lvl_d_2_uint_d_ack_ge <= ip(194);
  oper_tmp_d_179_d_lvl_d_2_uint_d_req_ge <= '1';
  op(198) <= oper_tmp_d_179_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_188_d_id_d_1_uint_d_ack_ge <= ip(202);
  oper_tmp_d_188_d_id_d_1_uint_d_req_ge <= '1';
  op(205) <= oper_tmp_d_188_d_id_d_1_uint_d_req_top;
  oper_tmp_d_188_d_lvl_d_1_uint_d_ack_ge <= ip(203);
  oper_tmp_d_188_d_lvl_d_1_uint_d_req_ge <= '1';
  op(206) <= oper_tmp_d_188_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_188_d_lvl_d_2_uint_d_ack_ge <= ip(205);
  oper_tmp_d_188_d_lvl_d_2_uint_d_req_ge <= '1';
  op(208) <= oper_tmp_d_188_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_192_d_id_d_1_uint_d_ack_ge <= ip(206);
  oper_tmp_d_192_d_id_d_1_uint_d_req_ge <= '1';
  op(209) <= oper_tmp_d_192_d_id_d_1_uint_d_req_top;
  oper_tmp_d_192_d_lvl_d_1_uint_d_ack_ge <= ip(207);
  oper_tmp_d_192_d_lvl_d_1_uint_d_req_ge <= '1';
  op(210) <= oper_tmp_d_192_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_192_d_lvl_d_2_uint_d_ack_ge <= ip(209);
  oper_tmp_d_192_d_lvl_d_2_uint_d_req_ge <= '1';
  op(212) <= oper_tmp_d_192_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_20299_bool_d_ack_ge <= ip(237);
  oper_tmp_d_20299_bool_d_req_ge <= '1';
  op(240) <= oper_tmp_d_20299_bool_d_req_top;
  oper_tmp_d_202_bool_d_ack_ge <= ip(223);
  oper_tmp_d_202_bool_d_req_ge <= '1';
  op(226) <= oper_tmp_d_202_bool_d_req_top;
  oper_tmp_d_206_d_lvl_d_0_uint_d_ack_ge <= ip(230);
  oper_tmp_d_206_d_lvl_d_0_uint_d_req_ge <= '1';
  op(233) <= oper_tmp_d_206_d_lvl_d_0_uint_d_req_top;
  oper_tmp_d_20_d_lvl_d_0_uint_d_ack_ge <= ip(27);
  oper_tmp_d_20_d_lvl_d_0_uint_d_req_ge <= '1';
  op(27) <= oper_tmp_d_20_d_lvl_d_0_uint_d_req_top;
  oper_tmp_d_210_d_id_d_1_uint_d_ack_ge <= ip(231);
  oper_tmp_d_210_d_id_d_1_uint_d_req_ge <= '1';
  op(234) <= oper_tmp_d_210_d_id_d_1_uint_d_req_top;
  oper_tmp_d_210_d_lvl_d_1_uint_d_ack_ge <= ip(232);
  oper_tmp_d_210_d_lvl_d_1_uint_d_req_ge <= '1';
  op(235) <= oper_tmp_d_210_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_210_d_lvl_d_2_uint_d_ack_ge <= ip(233);
  oper_tmp_d_210_d_lvl_d_2_uint_d_req_ge <= '1';
  op(236) <= oper_tmp_d_210_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_221111_bool_d_ack_ge <= ip(266);
  oper_tmp_d_221111_bool_d_req_ge <= '1';
  op(270) <= oper_tmp_d_221111_bool_d_req_top;
  oper_tmp_d_221_bool_d_ack_ge <= ip(250);
  oper_tmp_d_221_bool_d_req_ge <= '1';
  op(254) <= oper_tmp_d_221_bool_d_req_top;
  oper_tmp_d_225_d_lvl_d_0_uint_d_ack_ge <= ip(259);
  oper_tmp_d_225_d_lvl_d_0_uint_d_req_ge <= '1';
  op(263) <= oper_tmp_d_225_d_lvl_d_0_uint_d_req_top;
  oper_tmp_d_229_d_id_d_1_uint_d_ack_ge <= ip(260);
  oper_tmp_d_229_d_id_d_1_uint_d_req_ge <= '1';
  op(264) <= oper_tmp_d_229_d_id_d_1_uint_d_req_top;
  oper_tmp_d_229_d_lvl_d_1_uint_d_ack_ge <= ip(261);
  oper_tmp_d_229_d_lvl_d_1_uint_d_req_ge <= '1';
  op(265) <= oper_tmp_d_229_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_229_d_lvl_d_2_uint_d_ack_ge <= ip(262);
  oper_tmp_d_229_d_lvl_d_2_uint_d_req_ge <= '1';
  op(266) <= oper_tmp_d_229_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_25_d_lvl_d_0_uint_d_ack_ge <= ip(29);
  oper_tmp_d_25_d_lvl_d_0_uint_d_req_ge <= '1';
  op(29) <= oper_tmp_d_25_d_lvl_d_0_uint_d_req_top;
  oper_tmp_d_27_d_id_d_1_uint_d_ack_ge <= ip(32);
  oper_tmp_d_27_d_id_d_1_uint_d_req_ge <= '1';
  op(32) <= oper_tmp_d_27_d_id_d_1_uint_d_req_top;
  oper_tmp_d_27_d_lvl_d_1_uint_d_ack_ge <= ip(33);
  oper_tmp_d_27_d_lvl_d_1_uint_d_req_ge <= '1';
  op(33) <= oper_tmp_d_27_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_27_d_lvl_d_2_uint_d_ack_ge <= ip(35);
  oper_tmp_d_27_d_lvl_d_2_uint_d_req_ge <= '1';
  op(35) <= oper_tmp_d_27_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_30_d_lvl_d_0_uint_d_ack_ge <= ip(36);
  oper_tmp_d_30_d_lvl_d_0_uint_d_req_ge <= '1';
  op(36) <= oper_tmp_d_30_d_lvl_d_0_uint_d_req_top;
  oper_tmp_d_4223_bool_d_ack_ge <= ip(72);
  oper_tmp_d_4223_bool_d_req_ge <= '1';
  op(76) <= oper_tmp_d_4223_bool_d_req_top;
  oper_tmp_d_42_bool_d_ack_ge <= ip(54);
  oper_tmp_d_42_bool_d_req_ge <= '1';
  op(58) <= oper_tmp_d_42_bool_d_req_top;
  oper_tmp_d_47_d_id_d_1_uint_d_ack_ge <= ip(64);
  oper_tmp_d_47_d_id_d_1_uint_d_req_ge <= '1';
  op(69) <= oper_tmp_d_47_d_id_d_1_uint_d_req_top;
  oper_tmp_d_47_d_lvl_d_1_uint_d_ack_ge <= ip(65);
  oper_tmp_d_47_d_lvl_d_1_uint_d_req_ge <= '1';
  op(70) <= oper_tmp_d_47_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_47_d_lvl_d_2_uint_d_ack_ge <= ip(66);
  oper_tmp_d_47_d_lvl_d_2_uint_d_req_ge <= '1';
  op(71) <= oper_tmp_d_47_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_52_d_id_d_1_uint_d_ack_ge <= ip(48);
  oper_tmp_d_52_d_id_d_1_uint_d_req_ge <= '1';
  op(50) <= oper_tmp_d_52_d_id_d_1_uint_d_req_top;
  oper_tmp_d_52_d_lvl_d_1_uint_d_ack_ge <= ip(49);
  oper_tmp_d_52_d_lvl_d_1_uint_d_req_ge <= '1';
  op(51) <= oper_tmp_d_52_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_52_d_lvl_d_2_uint_d_ack_ge <= ip(50);
  oper_tmp_d_52_d_lvl_d_2_uint_d_req_ge <= '1';
  op(52) <= oper_tmp_d_52_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_54_bool_d_ack_ge <= ip(68);
  oper_tmp_d_54_bool_d_req_ge <= '1';
  op(73) <= oper_tmp_d_54_bool_d_req_top;
  oper_tmp_d_65_d_id_d_1_uint_d_ack_ge <= ip(78);
  oper_tmp_d_65_d_id_d_1_uint_d_req_ge <= '1';
  op(83) <= oper_tmp_d_65_d_id_d_1_uint_d_req_top;
  oper_tmp_d_65_d_lvl_d_1_uint_d_ack_ge <= ip(79);
  oper_tmp_d_65_d_lvl_d_1_uint_d_req_ge <= '1';
  op(84) <= oper_tmp_d_65_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_65_d_lvl_d_2_uint_d_ack_ge <= ip(80);
  oper_tmp_d_65_d_lvl_d_2_uint_d_req_ge <= '1';
  op(85) <= oper_tmp_d_65_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_74_d_id_d_1_uint_d_ack_ge <= ip(83);
  oper_tmp_d_74_d_id_d_1_uint_d_req_ge <= '1';
  op(88) <= oper_tmp_d_74_d_id_d_1_uint_d_req_top;
  oper_tmp_d_74_d_lvl_d_1_uint_d_ack_ge <= ip(84);
  oper_tmp_d_74_d_lvl_d_1_uint_d_req_ge <= '1';
  op(89) <= oper_tmp_d_74_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_74_d_lvl_d_2_uint_d_ack_ge <= ip(85);
  oper_tmp_d_74_d_lvl_d_2_uint_d_req_ge <= '1';
  op(90) <= oper_tmp_d_74_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_92_bool_d_ack_ge <= ip(111);
  oper_tmp_d_92_bool_d_req_ge <= '1';
  op(117) <= oper_tmp_d_92_bool_d_req_top;
  oper_tmp_d_97_d_id_d_1_uint_d_ack_ge <= ip(115);
  oper_tmp_d_97_d_id_d_1_uint_d_req_ge <= '1';
  op(120) <= oper_tmp_d_97_d_id_d_1_uint_d_req_top;
  oper_tmp_d_97_d_lvl_d_1_uint_d_ack_ge <= ip(116);
  oper_tmp_d_97_d_lvl_d_1_uint_d_req_ge <= '1';
  op(121) <= oper_tmp_d_97_d_lvl_d_1_uint_d_req_top;
  oper_tmp_d_97_d_lvl_d_2_uint_d_ack_ge <= ip(117);
  oper_tmp_d_97_d_lvl_d_2_uint_d_req_ge <= '1';
  op(122) <= oper_tmp_d_97_d_lvl_d_2_uint_d_req_top;
  oper_tmp_d_uint_d_ack_ge <= ip(59);
  oper_tmp_d_uint_d_req_ge <= '1';
  op(62) <= oper_tmp_d_uint_d_req_top;
  start_call_divide_0_actual_0_wr_d_ack_ge <= ip(121);
  start_call_divide_0_actual_0_wr_d_req_ge <= '1';
  op(126) <= start_call_divide_0_actual_0_wr_d_req_top;
  start_call_divide_0_actual_1_wr_d_ack_ge <= ip(122);
  start_call_divide_0_actual_1_wr_d_req_ge <= '1';
  op(127) <= start_call_divide_0_actual_1_wr_d_req_top;
  start_call_divide_0_d_ack_ge <= ip(120);
  start_call_divide_0_d_req_ge <= '1';
  op(125) <= start_call_divide_0_d_req_top;
  store_0_d_ack_ge <= ip(13);
  store_0_d_req_ge <= '1';
  op(15) <= store_0_d_req_top;
  store_10_d_ack_ge <= ip(201);
  store_10_d_req_ge <= '1';
  op(204) <= store_10_d_req_top;
  store_11_d_ack_ge <= ip(211);
  store_11_d_req_ge <= '1';
  op(214) <= store_11_d_req_top;
  store_12_d_ack_ge <= ip(235);
  store_12_d_req_ge <= '1';
  op(238) <= store_12_d_req_top;
  store_13_d_ack_ge <= ip(264);
  store_13_d_req_ge <= '1';
  op(268) <= store_13_d_req_top;
  store_1_d_ack_ge <= ip(38);
  store_1_d_req_ge <= '1';
  op(38) <= store_1_d_req_top;
  store_2_d_ack_ge <= ip(87);
  store_2_d_req_ge <= '1';
  op(92) <= store_2_d_req_top;
  store_3_d_ack_ge <= ip(88);
  store_3_d_req_ge <= '1';
  op(93) <= store_3_d_req_top;
  store_4_d_ack_ge <= ip(124);
  store_4_d_req_ge <= '1';
  op(129) <= store_4_d_req_top;
  store_5_d_ack_ge <= ip(143);
  store_5_d_req_ge <= '1';
  op(148) <= store_5_d_req_top;
  store_6_d_ack_ge <= ip(167);
  store_6_d_req_ge <= '1';
  op(171) <= store_6_d_req_top;
  store_7_d_ack_ge <= ip(172);
  store_7_d_req_ge <= '1';
  op(176) <= store_7_d_req_top;
  store_8_d_ack_ge <= ip(186);
  store_8_d_req_ge <= '1';
  op(190) <= store_8_d_req_top;
  store_9_d_ack_ge <= ip(196);
  store_9_d_req_ge <= '1';
  op(200) <= store_9_d_req_top;
  tc_i_d_1_d_0_d_ack_ge <= ip(26);
  tc_i_d_1_d_0_d_req_ge <= '1';
  op(26) <= tc_i_d_1_d_0_d_req_top;
  tc_i_d_2_d_0_d_ph_d_ack_ge <= ip(47);
  tc_i_d_2_d_0_d_ph_d_req_ge <= '1';
  op(49) <= tc_i_d_2_d_0_d_ph_d_req_top;
  tc_i_d_3_d_0_d_ph_d_ack_ge <= ip(153);
  tc_i_d_3_d_0_d_ph_d_req_ge <= '1';
  op(157) <= tc_i_d_3_d_0_d_ph_d_req_top;
  tc_i_d_4_d_0_d_ack_ge <= ip(222);
  tc_i_d_4_d_0_d_req_ge <= '1';
  op(225) <= tc_i_d_4_d_0_d_req_top;
  tc_i_d_5_d_0_d_ack_ge <= ip(249);
  tc_i_d_5_d_0_d_req_ge <= '1';
  op(253) <= tc_i_d_5_d_0_d_req_top;
  tc_indvar138_d_ack_ge <= ip(108);
  tc_indvar138_d_req_ge <= '1';
  op(114) <= tc_indvar138_d_req_top;
  tc_indvar151_d_ack_ge <= ip(254);
  tc_indvar151_d_req_ge <= '1';
  op(258) <= tc_indvar151_d_req_top;
  tc_j_d_11_d_2_d_ack_ge <= ip(227);
  tc_j_d_11_d_2_d_req_ge <= '1';
  op(230) <= tc_j_d_11_d_2_d_req_top;
  tc_j_d_13_d_2_d_ack_ge <= ip(256);
  tc_j_d_13_d_2_d_req_ge <= '1';
  op(260) <= tc_j_d_13_d_2_d_req_top;
  tc_j_d_3_d_2_d_ack_ge <= ip(63);
  tc_j_d_3_d_2_d_req_ge <= '1';
  op(68) <= tc_j_d_3_d_2_d_req_top;
  tc_j_d_3_d_in_d_ack_ge <= ip(57);
  tc_j_d_3_d_in_d_req_ge <= '1';
  op(60) <= tc_j_d_3_d_in_d_req_top;
  tc_j_d_7_d_1_d_ack_ge <= ip(130);
  tc_j_d_7_d_1_d_req_ge <= '1';
  op(135) <= tc_j_d_7_d_1_d_req_top;
  tc_p_d_0_d_0_d_ph_d_ack_ge <= ip(100);
  tc_p_d_0_d_0_d_ph_d_req_ge <= '1';
  op(105) <= tc_p_d_0_d_0_d_ph_d_req_top;
  tc_tmp_d_118_d_id_d_1_d_cast_d_ack_ge <= ip(131);
  tc_tmp_d_118_d_id_d_1_d_cast_d_req_ge <= '1';
  op(136) <= tc_tmp_d_118_d_id_d_1_d_cast_d_req_top;
  tc_tmp_d_154_d_id_d_2_d_cast_d_ack_ge <= ip(160);
  tc_tmp_d_154_d_id_d_2_d_cast_d_req_ge <= '1';
  op(164) <= tc_tmp_d_154_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_158_d_id_d_2_d_cast_d_ack_ge <= ip(164);
  tc_tmp_d_158_d_id_d_2_d_cast_d_req_ge <= '1';
  op(168) <= tc_tmp_d_158_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_163_d_id_d_2_d_cast_d_ack_ge <= ip(170);
  tc_tmp_d_163_d_id_d_2_d_cast_d_req_ge <= '1';
  op(174) <= tc_tmp_d_163_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_171_d_id_d_2_d_cast_d_ack_ge <= ip(182);
  tc_tmp_d_171_d_id_d_2_d_cast_d_req_ge <= '1';
  op(187) <= tc_tmp_d_171_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_175_d_id_d_2_d_cast_d_ack_ge <= ip(189);
  tc_tmp_d_175_d_id_d_2_d_cast_d_req_ge <= '1';
  op(193) <= tc_tmp_d_175_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_179_d_id_d_2_d_cast_d_ack_ge <= ip(193);
  tc_tmp_d_179_d_id_d_2_d_cast_d_req_ge <= '1';
  op(197) <= tc_tmp_d_179_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_188_d_id_d_2_d_cast_d_ack_ge <= ip(204);
  tc_tmp_d_188_d_id_d_2_d_cast_d_req_ge <= '1';
  op(207) <= tc_tmp_d_188_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_192_d_id_d_2_d_cast_d_ack_ge <= ip(208);
  tc_tmp_d_192_d_id_d_2_d_cast_d_req_ge <= '1';
  op(211) <= tc_tmp_d_192_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_206_d_id_d_0_d_cast_d_ack_ge <= ip(229);
  tc_tmp_d_206_d_id_d_0_d_cast_d_req_ge <= '1';
  op(232) <= tc_tmp_d_206_d_id_d_0_d_cast_d_req_top;
  tc_tmp_d_225_d_id_d_0_d_cast_d_ack_ge <= ip(258);
  tc_tmp_d_225_d_id_d_0_d_cast_d_req_ge <= '1';
  op(262) <= tc_tmp_d_225_d_id_d_0_d_cast_d_req_top;
  tc_tmp_d_27_d_id_d_1_d_cast_d_ack_ge <= ip(31);
  tc_tmp_d_27_d_id_d_1_d_cast_d_req_ge <= '1';
  op(31) <= tc_tmp_d_27_d_id_d_1_d_cast_d_req_top;
  tc_tmp_d_27_d_id_d_2_d_cast_d_ack_ge <= ip(34);
  tc_tmp_d_27_d_id_d_2_d_cast_d_req_ge <= '1';
  op(34) <= tc_tmp_d_27_d_id_d_2_d_cast_d_req_top;
  tc_tmp_d_74_d_id_d_1_d_cast_d_ack_ge <= ip(82);
  tc_tmp_d_74_d_id_d_1_d_cast_d_req_ge <= '1';
  op(87) <= tc_tmp_d_74_d_id_d_1_d_cast_d_req_top;
  tc_tmp_d_97_d_id_d_1_d_cast_d_ack_ge <= ip(114);
  tc_tmp_d_97_d_id_d_1_d_cast_d_req_ge <= '1';
  op(119) <= tc_tmp_d_97_d_id_d_1_d_cast_d_req_top;
  then_d_0_d_entry_ge <= '1';
  then_d_0_to_no_exit_d_4_src_ge <= ip(74);
  then_d_0_to_no_exit_d_5_d_preheader_d_loopexit_src_ge <= ip(75);
  then_d_1_d_entry_ge <= '1';
  then_d_1_to_loopexit_d_10_src_ge <= ip(176);
  then_d_1_to_no_exit_d_10_d_backedge_src_ge <= ip(175);
  then_d_2_d_entry_ge <= '1';
  then_d_2_to_loopexit_d_10_src_ge <= ip(200);
  then_d_2_to_no_exit_d_10_d_backedge_src_ge <= ip(199);

end behavioral;
