
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;

entity test_floats_ln is
  port(
    clk : in std_logic;
    reset : in std_logic;
    test_floats_cp_LambdaIn : out BooleanArray(323 downto 1);
    test_floats_cp_LambdaOut : in BooleanArray(323 downto 1);
    test_floats_dp_SigmaIn : out BooleanArray(323 downto 1);
    test_floats_dp_SigmaOut : in BooleanArray(323 downto 1));
end test_floats_ln;

architecture default_arch of test_floats_ln is
begin
  test_floats_cp_LambdaIn(1) <= test_floats_dp_SigmaOut(1);
  test_floats_cp_LambdaIn(2) <= test_floats_dp_SigmaOut(2);
  test_floats_cp_LambdaIn(3) <= test_floats_dp_SigmaOut(3);
  test_floats_cp_LambdaIn(4) <= test_floats_dp_SigmaOut(4);
  test_floats_cp_LambdaIn(5) <= test_floats_dp_SigmaOut(5);
  test_floats_cp_LambdaIn(6) <= test_floats_dp_SigmaOut(6);
  test_floats_cp_LambdaIn(7) <= test_floats_dp_SigmaOut(7);
  test_floats_cp_LambdaIn(8) <= test_floats_dp_SigmaOut(8);
  test_floats_cp_LambdaIn(9) <= test_floats_dp_SigmaOut(9);
  test_floats_cp_LambdaIn(10) <= test_floats_dp_SigmaOut(10);
  test_floats_cp_LambdaIn(11) <= test_floats_dp_SigmaOut(11);
  test_floats_cp_LambdaIn(12) <= test_floats_dp_SigmaOut(12);
  test_floats_cp_LambdaIn(13) <= test_floats_dp_SigmaOut(13);
  test_floats_cp_LambdaIn(14) <= test_floats_dp_SigmaOut(14);
  test_floats_cp_LambdaIn(15) <= test_floats_dp_SigmaOut(15);
  test_floats_cp_LambdaIn(16) <= test_floats_dp_SigmaOut(16);
  test_floats_cp_LambdaIn(17) <= test_floats_dp_SigmaOut(17);
  test_floats_cp_LambdaIn(18) <= test_floats_dp_SigmaOut(18);
  test_floats_cp_LambdaIn(19) <= test_floats_dp_SigmaOut(19);
  test_floats_cp_LambdaIn(20) <= test_floats_dp_SigmaOut(20);
  test_floats_cp_LambdaIn(21) <= test_floats_dp_SigmaOut(21);
  test_floats_cp_LambdaIn(22) <= test_floats_dp_SigmaOut(22);
  test_floats_cp_LambdaIn(23) <= test_floats_dp_SigmaOut(23);
  test_floats_cp_LambdaIn(24) <= test_floats_dp_SigmaOut(24);
  test_floats_cp_LambdaIn(25) <= test_floats_dp_SigmaOut(25);
  test_floats_cp_LambdaIn(26) <= test_floats_dp_SigmaOut(26);
  test_floats_cp_LambdaIn(27) <= test_floats_dp_SigmaOut(27);
  test_floats_cp_LambdaIn(28) <= test_floats_dp_SigmaOut(28);
  test_floats_cp_LambdaIn(29) <= test_floats_dp_SigmaOut(29);
  test_floats_cp_LambdaIn(30) <= test_floats_dp_SigmaOut(30);
  test_floats_cp_LambdaIn(31) <= test_floats_dp_SigmaOut(31);
  test_floats_cp_LambdaIn(32) <= test_floats_dp_SigmaOut(32);
  test_floats_cp_LambdaIn(33) <= test_floats_dp_SigmaOut(33);
  test_floats_cp_LambdaIn(34) <= test_floats_dp_SigmaOut(34);
  test_floats_cp_LambdaIn(35) <= test_floats_dp_SigmaOut(35);
  test_floats_cp_LambdaIn(36) <= test_floats_dp_SigmaOut(36);
  test_floats_cp_LambdaIn(37) <= test_floats_dp_SigmaOut(37);
  test_floats_cp_LambdaIn(38) <= test_floats_dp_SigmaOut(38);
  test_floats_cp_LambdaIn(39) <= test_floats_dp_SigmaOut(39);
  test_floats_cp_LambdaIn(40) <= test_floats_dp_SigmaOut(40);
  test_floats_cp_LambdaIn(41) <= test_floats_dp_SigmaOut(41);
  test_floats_cp_LambdaIn(42) <= test_floats_dp_SigmaOut(42);
  test_floats_cp_LambdaIn(43) <= test_floats_dp_SigmaOut(43);
  test_floats_cp_LambdaIn(44) <= test_floats_dp_SigmaOut(44);
  test_floats_cp_LambdaIn(45) <= test_floats_dp_SigmaOut(45);
  test_floats_cp_LambdaIn(46) <= test_floats_dp_SigmaOut(46);
  test_floats_cp_LambdaIn(47) <= test_floats_dp_SigmaOut(47);
  test_floats_cp_LambdaIn(48) <= test_floats_dp_SigmaOut(48);
  test_floats_cp_LambdaIn(49) <= test_floats_dp_SigmaOut(49);
  test_floats_cp_LambdaIn(50) <= test_floats_dp_SigmaOut(50);
  test_floats_cp_LambdaIn(51) <= test_floats_dp_SigmaOut(51);
  test_floats_cp_LambdaIn(52) <= test_floats_dp_SigmaOut(52);
  test_floats_cp_LambdaIn(53) <= test_floats_dp_SigmaOut(53);
  test_floats_cp_LambdaIn(54) <= test_floats_dp_SigmaOut(54);
  test_floats_cp_LambdaIn(55) <= test_floats_dp_SigmaOut(55);
  test_floats_cp_LambdaIn(56) <= test_floats_dp_SigmaOut(56);
  test_floats_cp_LambdaIn(57) <= test_floats_dp_SigmaOut(57);
  test_floats_cp_LambdaIn(58) <= test_floats_dp_SigmaOut(58);
  test_floats_cp_LambdaIn(59) <= test_floats_dp_SigmaOut(59);
  test_floats_cp_LambdaIn(60) <= test_floats_dp_SigmaOut(60);
  test_floats_cp_LambdaIn(61) <= test_floats_dp_SigmaOut(61);
  test_floats_cp_LambdaIn(62) <= test_floats_dp_SigmaOut(62);
  test_floats_cp_LambdaIn(63) <= test_floats_dp_SigmaOut(63);
  test_floats_cp_LambdaIn(64) <= test_floats_dp_SigmaOut(64);
  test_floats_cp_LambdaIn(65) <= test_floats_dp_SigmaOut(65);
  test_floats_cp_LambdaIn(66) <= test_floats_dp_SigmaOut(66);
  test_floats_cp_LambdaIn(67) <= test_floats_dp_SigmaOut(67);
  test_floats_cp_LambdaIn(68) <= test_floats_dp_SigmaOut(68);
  test_floats_cp_LambdaIn(69) <= test_floats_dp_SigmaOut(69);
  test_floats_cp_LambdaIn(70) <= test_floats_dp_SigmaOut(70);
  test_floats_cp_LambdaIn(71) <= test_floats_dp_SigmaOut(71);
  test_floats_cp_LambdaIn(72) <= test_floats_dp_SigmaOut(72);
  test_floats_cp_LambdaIn(73) <= test_floats_dp_SigmaOut(73);
  test_floats_cp_LambdaIn(74) <= test_floats_dp_SigmaOut(74);
  test_floats_cp_LambdaIn(75) <= test_floats_dp_SigmaOut(75);
  test_floats_cp_LambdaIn(76) <= test_floats_dp_SigmaOut(76);
  test_floats_cp_LambdaIn(77) <= test_floats_dp_SigmaOut(77);
  test_floats_cp_LambdaIn(78) <= test_floats_dp_SigmaOut(78);
  test_floats_cp_LambdaIn(79) <= test_floats_dp_SigmaOut(79);
  test_floats_cp_LambdaIn(80) <= test_floats_dp_SigmaOut(80);
  test_floats_cp_LambdaIn(81) <= test_floats_dp_SigmaOut(81);
  test_floats_cp_LambdaIn(82) <= test_floats_dp_SigmaOut(82);
  test_floats_cp_LambdaIn(83) <= test_floats_dp_SigmaOut(83);
  test_floats_cp_LambdaIn(84) <= test_floats_dp_SigmaOut(84);
  test_floats_cp_LambdaIn(85) <= test_floats_dp_SigmaOut(85);
  test_floats_cp_LambdaIn(86) <= test_floats_dp_SigmaOut(86);
  test_floats_cp_LambdaIn(87) <= test_floats_dp_SigmaOut(87);
  test_floats_cp_LambdaIn(88) <= test_floats_dp_SigmaOut(88);
  test_floats_cp_LambdaIn(89) <= test_floats_dp_SigmaOut(89);
  test_floats_cp_LambdaIn(90) <= test_floats_dp_SigmaOut(90);
  test_floats_cp_LambdaIn(91) <= test_floats_dp_SigmaOut(91);
  test_floats_cp_LambdaIn(92) <= test_floats_dp_SigmaOut(92);
  test_floats_cp_LambdaIn(93) <= test_floats_dp_SigmaOut(93);
  test_floats_cp_LambdaIn(94) <= test_floats_dp_SigmaOut(94);
  test_floats_cp_LambdaIn(95) <= test_floats_dp_SigmaOut(95);
  test_floats_cp_LambdaIn(96) <= test_floats_dp_SigmaOut(96);
  test_floats_cp_LambdaIn(97) <= test_floats_dp_SigmaOut(97);
  test_floats_cp_LambdaIn(98) <= test_floats_dp_SigmaOut(98);
  test_floats_cp_LambdaIn(99) <= test_floats_dp_SigmaOut(99);
  test_floats_cp_LambdaIn(100) <= test_floats_dp_SigmaOut(100);
  test_floats_cp_LambdaIn(101) <= test_floats_dp_SigmaOut(101);
  test_floats_cp_LambdaIn(102) <= test_floats_dp_SigmaOut(102);
  test_floats_cp_LambdaIn(103) <= test_floats_dp_SigmaOut(103);
  test_floats_cp_LambdaIn(104) <= test_floats_dp_SigmaOut(104);
  test_floats_cp_LambdaIn(105) <= test_floats_dp_SigmaOut(105);
  test_floats_cp_LambdaIn(106) <= test_floats_dp_SigmaOut(106);
  test_floats_cp_LambdaIn(107) <= test_floats_dp_SigmaOut(107);
  test_floats_cp_LambdaIn(108) <= test_floats_dp_SigmaOut(108);
  test_floats_cp_LambdaIn(109) <= test_floats_dp_SigmaOut(109);
  test_floats_cp_LambdaIn(110) <= test_floats_dp_SigmaOut(110);
  test_floats_cp_LambdaIn(111) <= test_floats_dp_SigmaOut(111);
  test_floats_cp_LambdaIn(112) <= test_floats_dp_SigmaOut(112);
  test_floats_cp_LambdaIn(113) <= test_floats_dp_SigmaOut(113);
  test_floats_cp_LambdaIn(114) <= test_floats_dp_SigmaOut(114);
  test_floats_cp_LambdaIn(115) <= test_floats_dp_SigmaOut(115);
  test_floats_cp_LambdaIn(116) <= test_floats_dp_SigmaOut(116);
  test_floats_cp_LambdaIn(117) <= test_floats_dp_SigmaOut(117);
  test_floats_cp_LambdaIn(118) <= test_floats_dp_SigmaOut(118);
  test_floats_cp_LambdaIn(119) <= test_floats_dp_SigmaOut(119);
  test_floats_cp_LambdaIn(120) <= test_floats_dp_SigmaOut(120);
  test_floats_cp_LambdaIn(121) <= test_floats_dp_SigmaOut(121);
  test_floats_cp_LambdaIn(122) <= test_floats_dp_SigmaOut(122);
  test_floats_cp_LambdaIn(123) <= test_floats_dp_SigmaOut(123);
  test_floats_cp_LambdaIn(124) <= test_floats_dp_SigmaOut(124);
  test_floats_cp_LambdaIn(125) <= test_floats_dp_SigmaOut(125);
  test_floats_cp_LambdaIn(126) <= test_floats_dp_SigmaOut(126);
  test_floats_cp_LambdaIn(127) <= test_floats_dp_SigmaOut(127);
  test_floats_cp_LambdaIn(128) <= test_floats_dp_SigmaOut(128);
  test_floats_cp_LambdaIn(129) <= test_floats_dp_SigmaOut(129);
  test_floats_cp_LambdaIn(130) <= test_floats_dp_SigmaOut(130);
  test_floats_cp_LambdaIn(131) <= test_floats_dp_SigmaOut(131);
  test_floats_cp_LambdaIn(132) <= test_floats_dp_SigmaOut(132);
  test_floats_cp_LambdaIn(133) <= test_floats_dp_SigmaOut(133);
  test_floats_cp_LambdaIn(134) <= test_floats_dp_SigmaOut(134);
  test_floats_cp_LambdaIn(135) <= test_floats_dp_SigmaOut(135);
  test_floats_cp_LambdaIn(136) <= test_floats_dp_SigmaOut(136);
  test_floats_cp_LambdaIn(137) <= test_floats_dp_SigmaOut(137);
  test_floats_cp_LambdaIn(138) <= test_floats_dp_SigmaOut(138);
  test_floats_cp_LambdaIn(139) <= test_floats_dp_SigmaOut(139);
  test_floats_cp_LambdaIn(140) <= test_floats_dp_SigmaOut(140);
  test_floats_cp_LambdaIn(141) <= test_floats_dp_SigmaOut(141);
  test_floats_cp_LambdaIn(142) <= test_floats_dp_SigmaOut(142);
  test_floats_cp_LambdaIn(143) <= test_floats_dp_SigmaOut(143);
  test_floats_cp_LambdaIn(144) <= test_floats_dp_SigmaOut(144);
  test_floats_cp_LambdaIn(145) <= test_floats_dp_SigmaOut(145);
  test_floats_cp_LambdaIn(146) <= test_floats_dp_SigmaOut(146);
  test_floats_cp_LambdaIn(147) <= test_floats_dp_SigmaOut(147);
  test_floats_cp_LambdaIn(148) <= test_floats_dp_SigmaOut(148);
  test_floats_cp_LambdaIn(149) <= test_floats_dp_SigmaOut(149);
  test_floats_cp_LambdaIn(150) <= test_floats_dp_SigmaOut(150);
  test_floats_cp_LambdaIn(151) <= test_floats_dp_SigmaOut(151);
  test_floats_cp_LambdaIn(152) <= test_floats_dp_SigmaOut(152);
  test_floats_cp_LambdaIn(153) <= test_floats_dp_SigmaOut(153);
  test_floats_cp_LambdaIn(154) <= test_floats_dp_SigmaOut(154);
  test_floats_cp_LambdaIn(155) <= test_floats_dp_SigmaOut(155);
  test_floats_cp_LambdaIn(156) <= test_floats_dp_SigmaOut(156);
  test_floats_cp_LambdaIn(157) <= test_floats_dp_SigmaOut(157);
  test_floats_cp_LambdaIn(158) <= test_floats_dp_SigmaOut(158);
  test_floats_cp_LambdaIn(159) <= test_floats_dp_SigmaOut(159);
  test_floats_cp_LambdaIn(160) <= test_floats_dp_SigmaOut(160);
  test_floats_cp_LambdaIn(161) <= test_floats_dp_SigmaOut(161);
  test_floats_cp_LambdaIn(162) <= test_floats_dp_SigmaOut(162);
  test_floats_cp_LambdaIn(163) <= test_floats_dp_SigmaOut(163);
  test_floats_cp_LambdaIn(164) <= test_floats_dp_SigmaOut(164);
  test_floats_cp_LambdaIn(165) <= test_floats_dp_SigmaOut(165);
  test_floats_cp_LambdaIn(166) <= test_floats_dp_SigmaOut(166);
  test_floats_cp_LambdaIn(167) <= test_floats_dp_SigmaOut(167);
  test_floats_cp_LambdaIn(168) <= test_floats_dp_SigmaOut(168);
  test_floats_cp_LambdaIn(169) <= test_floats_dp_SigmaOut(169);
  test_floats_cp_LambdaIn(170) <= test_floats_dp_SigmaOut(170);
  test_floats_cp_LambdaIn(171) <= test_floats_dp_SigmaOut(171);
  test_floats_cp_LambdaIn(172) <= test_floats_dp_SigmaOut(172);
  test_floats_cp_LambdaIn(173) <= test_floats_dp_SigmaOut(173);
  test_floats_cp_LambdaIn(174) <= test_floats_dp_SigmaOut(174);
  test_floats_cp_LambdaIn(175) <= test_floats_dp_SigmaOut(175);
  test_floats_cp_LambdaIn(176) <= test_floats_dp_SigmaOut(176);
  test_floats_cp_LambdaIn(177) <= test_floats_dp_SigmaOut(177);
  test_floats_cp_LambdaIn(178) <= test_floats_dp_SigmaOut(178);
  test_floats_cp_LambdaIn(179) <= test_floats_dp_SigmaOut(179);
  test_floats_cp_LambdaIn(180) <= test_floats_dp_SigmaOut(180);
  test_floats_cp_LambdaIn(181) <= test_floats_dp_SigmaOut(181);
  test_floats_cp_LambdaIn(182) <= test_floats_dp_SigmaOut(182);
  test_floats_cp_LambdaIn(183) <= test_floats_dp_SigmaOut(183);
  test_floats_cp_LambdaIn(184) <= test_floats_dp_SigmaOut(184);
  test_floats_cp_LambdaIn(185) <= test_floats_dp_SigmaOut(185);
  test_floats_cp_LambdaIn(186) <= test_floats_dp_SigmaOut(186);
  test_floats_cp_LambdaIn(187) <= test_floats_dp_SigmaOut(187);
  test_floats_cp_LambdaIn(188) <= test_floats_dp_SigmaOut(188);
  test_floats_cp_LambdaIn(189) <= test_floats_dp_SigmaOut(189);
  test_floats_cp_LambdaIn(190) <= test_floats_dp_SigmaOut(190);
  test_floats_cp_LambdaIn(191) <= test_floats_dp_SigmaOut(191);
  test_floats_cp_LambdaIn(192) <= test_floats_dp_SigmaOut(192);
  test_floats_cp_LambdaIn(193) <= test_floats_dp_SigmaOut(193);
  test_floats_cp_LambdaIn(194) <= test_floats_dp_SigmaOut(194);
  test_floats_cp_LambdaIn(195) <= test_floats_dp_SigmaOut(195);
  test_floats_cp_LambdaIn(196) <= test_floats_dp_SigmaOut(196);
  test_floats_cp_LambdaIn(197) <= test_floats_dp_SigmaOut(197);
  test_floats_cp_LambdaIn(198) <= test_floats_dp_SigmaOut(198);
  test_floats_cp_LambdaIn(199) <= test_floats_dp_SigmaOut(199);
  test_floats_cp_LambdaIn(200) <= test_floats_dp_SigmaOut(200);
  test_floats_cp_LambdaIn(201) <= test_floats_dp_SigmaOut(201);
  test_floats_cp_LambdaIn(202) <= test_floats_dp_SigmaOut(202);
  test_floats_cp_LambdaIn(203) <= test_floats_dp_SigmaOut(203);
  test_floats_cp_LambdaIn(204) <= test_floats_dp_SigmaOut(204);
  test_floats_cp_LambdaIn(205) <= test_floats_dp_SigmaOut(205);
  test_floats_cp_LambdaIn(206) <= test_floats_dp_SigmaOut(206);
  test_floats_cp_LambdaIn(207) <= test_floats_dp_SigmaOut(207);
  test_floats_cp_LambdaIn(208) <= test_floats_dp_SigmaOut(208);
  test_floats_cp_LambdaIn(209) <= test_floats_dp_SigmaOut(209);
  test_floats_cp_LambdaIn(210) <= test_floats_dp_SigmaOut(210);
  test_floats_cp_LambdaIn(211) <= test_floats_dp_SigmaOut(211);
  test_floats_cp_LambdaIn(212) <= test_floats_dp_SigmaOut(212);
  test_floats_cp_LambdaIn(213) <= test_floats_dp_SigmaOut(213);
  test_floats_cp_LambdaIn(214) <= test_floats_dp_SigmaOut(214);
  test_floats_cp_LambdaIn(215) <= test_floats_dp_SigmaOut(215);
  test_floats_cp_LambdaIn(216) <= test_floats_dp_SigmaOut(216);
  test_floats_cp_LambdaIn(217) <= test_floats_dp_SigmaOut(217);
  test_floats_cp_LambdaIn(218) <= test_floats_dp_SigmaOut(218);
  test_floats_cp_LambdaIn(219) <= test_floats_dp_SigmaOut(219);
  test_floats_cp_LambdaIn(220) <= test_floats_dp_SigmaOut(220);
  test_floats_cp_LambdaIn(221) <= test_floats_dp_SigmaOut(221);
  test_floats_cp_LambdaIn(222) <= test_floats_dp_SigmaOut(222);
  test_floats_cp_LambdaIn(223) <= test_floats_dp_SigmaOut(223);
  test_floats_cp_LambdaIn(224) <= test_floats_dp_SigmaOut(224);
  test_floats_cp_LambdaIn(225) <= test_floats_dp_SigmaOut(225);
  test_floats_cp_LambdaIn(226) <= test_floats_dp_SigmaOut(226);
  test_floats_cp_LambdaIn(227) <= test_floats_dp_SigmaOut(227);
  test_floats_cp_LambdaIn(228) <= test_floats_dp_SigmaOut(228);
  test_floats_cp_LambdaIn(229) <= test_floats_dp_SigmaOut(229);
  test_floats_cp_LambdaIn(230) <= test_floats_dp_SigmaOut(230);
  test_floats_cp_LambdaIn(231) <= test_floats_dp_SigmaOut(231);
  test_floats_cp_LambdaIn(232) <= test_floats_dp_SigmaOut(232);
  test_floats_cp_LambdaIn(233) <= test_floats_dp_SigmaOut(233);
  test_floats_cp_LambdaIn(234) <= test_floats_dp_SigmaOut(234);
  test_floats_cp_LambdaIn(235) <= test_floats_dp_SigmaOut(235);
  test_floats_cp_LambdaIn(236) <= test_floats_dp_SigmaOut(236);
  test_floats_cp_LambdaIn(237) <= test_floats_dp_SigmaOut(237);
  test_floats_cp_LambdaIn(238) <= test_floats_dp_SigmaOut(238);
  test_floats_cp_LambdaIn(239) <= test_floats_dp_SigmaOut(239);
  test_floats_cp_LambdaIn(240) <= test_floats_dp_SigmaOut(240);
  test_floats_cp_LambdaIn(241) <= test_floats_dp_SigmaOut(241);
  test_floats_cp_LambdaIn(242) <= test_floats_dp_SigmaOut(242);
  test_floats_cp_LambdaIn(243) <= test_floats_dp_SigmaOut(243);
  test_floats_cp_LambdaIn(244) <= test_floats_dp_SigmaOut(244);
  test_floats_cp_LambdaIn(245) <= test_floats_dp_SigmaOut(245);
  test_floats_cp_LambdaIn(246) <= test_floats_dp_SigmaOut(246);
  test_floats_cp_LambdaIn(247) <= test_floats_dp_SigmaOut(247);
  test_floats_cp_LambdaIn(248) <= test_floats_dp_SigmaOut(248);
  test_floats_cp_LambdaIn(249) <= test_floats_dp_SigmaOut(249);
  test_floats_cp_LambdaIn(250) <= test_floats_dp_SigmaOut(250);
  test_floats_cp_LambdaIn(251) <= test_floats_dp_SigmaOut(251);
  test_floats_cp_LambdaIn(252) <= test_floats_dp_SigmaOut(252);
  test_floats_cp_LambdaIn(253) <= test_floats_dp_SigmaOut(253);
  test_floats_cp_LambdaIn(254) <= test_floats_dp_SigmaOut(254);
  test_floats_cp_LambdaIn(255) <= test_floats_dp_SigmaOut(255);
  test_floats_cp_LambdaIn(256) <= test_floats_dp_SigmaOut(256);
  test_floats_cp_LambdaIn(257) <= test_floats_dp_SigmaOut(257);
  test_floats_cp_LambdaIn(258) <= test_floats_dp_SigmaOut(258);
  test_floats_cp_LambdaIn(259) <= test_floats_dp_SigmaOut(259);
  test_floats_cp_LambdaIn(260) <= test_floats_dp_SigmaOut(260);
  test_floats_cp_LambdaIn(261) <= test_floats_dp_SigmaOut(261);
  test_floats_cp_LambdaIn(262) <= test_floats_dp_SigmaOut(262);
  test_floats_cp_LambdaIn(263) <= test_floats_dp_SigmaOut(263);
  test_floats_cp_LambdaIn(264) <= test_floats_dp_SigmaOut(264);
  test_floats_cp_LambdaIn(265) <= test_floats_dp_SigmaOut(265);
  test_floats_cp_LambdaIn(266) <= test_floats_dp_SigmaOut(266);
  test_floats_cp_LambdaIn(267) <= test_floats_dp_SigmaOut(267);
  test_floats_cp_LambdaIn(268) <= test_floats_dp_SigmaOut(268);
  test_floats_cp_LambdaIn(269) <= test_floats_dp_SigmaOut(269);
  test_floats_cp_LambdaIn(270) <= test_floats_dp_SigmaOut(270);
  test_floats_cp_LambdaIn(271) <= test_floats_dp_SigmaOut(271);
  test_floats_cp_LambdaIn(272) <= test_floats_dp_SigmaOut(272);
  test_floats_cp_LambdaIn(273) <= test_floats_dp_SigmaOut(273);
  test_floats_cp_LambdaIn(274) <= test_floats_dp_SigmaOut(274);
  test_floats_cp_LambdaIn(275) <= test_floats_dp_SigmaOut(275);
  test_floats_cp_LambdaIn(276) <= test_floats_dp_SigmaOut(276);
  test_floats_cp_LambdaIn(277) <= test_floats_dp_SigmaOut(277);
  test_floats_cp_LambdaIn(278) <= test_floats_dp_SigmaOut(278);
  test_floats_cp_LambdaIn(279) <= test_floats_dp_SigmaOut(279);
  test_floats_cp_LambdaIn(280) <= test_floats_dp_SigmaOut(280);
  test_floats_cp_LambdaIn(281) <= test_floats_dp_SigmaOut(281);
  test_floats_cp_LambdaIn(282) <= test_floats_dp_SigmaOut(282);
  test_floats_cp_LambdaIn(283) <= test_floats_dp_SigmaOut(283);
  test_floats_cp_LambdaIn(284) <= test_floats_dp_SigmaOut(284);
  test_floats_cp_LambdaIn(285) <= test_floats_dp_SigmaOut(285);
  test_floats_cp_LambdaIn(286) <= test_floats_dp_SigmaOut(286);
  test_floats_cp_LambdaIn(287) <= test_floats_dp_SigmaOut(287);
  test_floats_cp_LambdaIn(288) <= test_floats_dp_SigmaOut(288);
  test_floats_cp_LambdaIn(289) <= test_floats_dp_SigmaOut(289);
  test_floats_cp_LambdaIn(290) <= test_floats_dp_SigmaOut(290);
  test_floats_cp_LambdaIn(291) <= test_floats_dp_SigmaOut(291);
  test_floats_cp_LambdaIn(292) <= test_floats_dp_SigmaOut(292);
  test_floats_cp_LambdaIn(293) <= test_floats_dp_SigmaOut(293);
  test_floats_cp_LambdaIn(294) <= test_floats_dp_SigmaOut(294);
  test_floats_cp_LambdaIn(295) <= test_floats_dp_SigmaOut(295);
  test_floats_cp_LambdaIn(296) <= test_floats_dp_SigmaOut(296);
  test_floats_cp_LambdaIn(297) <= test_floats_dp_SigmaOut(297);
  test_floats_cp_LambdaIn(298) <= test_floats_dp_SigmaOut(298);
  test_floats_cp_LambdaIn(299) <= test_floats_dp_SigmaOut(299);
  test_floats_cp_LambdaIn(300) <= test_floats_dp_SigmaOut(300);
  test_floats_cp_LambdaIn(301) <= test_floats_dp_SigmaOut(301);
  test_floats_cp_LambdaIn(302) <= test_floats_dp_SigmaOut(302);
  test_floats_cp_LambdaIn(303) <= test_floats_dp_SigmaOut(303);
  test_floats_cp_LambdaIn(304) <= test_floats_dp_SigmaOut(304);
  test_floats_cp_LambdaIn(305) <= test_floats_dp_SigmaOut(305);
  test_floats_cp_LambdaIn(306) <= test_floats_dp_SigmaOut(306);
  test_floats_cp_LambdaIn(307) <= test_floats_dp_SigmaOut(307);
  test_floats_cp_LambdaIn(308) <= test_floats_dp_SigmaOut(308);
  test_floats_cp_LambdaIn(309) <= test_floats_dp_SigmaOut(309);
  test_floats_cp_LambdaIn(310) <= test_floats_dp_SigmaOut(310);
  test_floats_cp_LambdaIn(311) <= test_floats_dp_SigmaOut(311);
  test_floats_cp_LambdaIn(312) <= test_floats_dp_SigmaOut(312);
  test_floats_cp_LambdaIn(313) <= test_floats_dp_SigmaOut(313);
  test_floats_cp_LambdaIn(314) <= test_floats_dp_SigmaOut(314);
  test_floats_cp_LambdaIn(315) <= test_floats_dp_SigmaOut(315);
  test_floats_cp_LambdaIn(316) <= test_floats_dp_SigmaOut(316);
  test_floats_cp_LambdaIn(317) <= test_floats_dp_SigmaOut(317);
  test_floats_cp_LambdaIn(318) <= test_floats_dp_SigmaOut(318);
  test_floats_cp_LambdaIn(319) <= test_floats_dp_SigmaOut(319);
  test_floats_cp_LambdaIn(320) <= test_floats_dp_SigmaOut(320);
  test_floats_cp_LambdaIn(321) <= test_floats_dp_SigmaOut(321);
  test_floats_cp_LambdaIn(322) <= test_floats_dp_SigmaOut(322);
  test_floats_cp_LambdaIn(323) <= test_floats_dp_SigmaOut(323);

  test_floats_dp_SigmaIn(1) <= test_floats_cp_LambdaOut(1);
  test_floats_dp_SigmaIn(2) <= test_floats_cp_LambdaOut(2);
  test_floats_dp_SigmaIn(3) <= test_floats_cp_LambdaOut(3);
  test_floats_dp_SigmaIn(4) <= test_floats_cp_LambdaOut(4);
  test_floats_dp_SigmaIn(5) <= test_floats_cp_LambdaOut(5);
  test_floats_dp_SigmaIn(6) <= test_floats_cp_LambdaOut(6);
  test_floats_dp_SigmaIn(7) <= test_floats_cp_LambdaOut(7);
  test_floats_dp_SigmaIn(8) <= test_floats_cp_LambdaOut(8);
  test_floats_dp_SigmaIn(9) <= test_floats_cp_LambdaOut(9);
  test_floats_dp_SigmaIn(10) <= test_floats_cp_LambdaOut(10);
  test_floats_dp_SigmaIn(11) <= test_floats_cp_LambdaOut(11);
  test_floats_dp_SigmaIn(12) <= test_floats_cp_LambdaOut(12);
  test_floats_dp_SigmaIn(13) <= test_floats_cp_LambdaOut(13);
  test_floats_dp_SigmaIn(14) <= test_floats_cp_LambdaOut(14);
  test_floats_dp_SigmaIn(15) <= test_floats_cp_LambdaOut(15);
  test_floats_dp_SigmaIn(16) <= test_floats_cp_LambdaOut(16);
  test_floats_dp_SigmaIn(17) <= test_floats_cp_LambdaOut(17);
  test_floats_dp_SigmaIn(18) <= test_floats_cp_LambdaOut(18);
  test_floats_dp_SigmaIn(19) <= test_floats_cp_LambdaOut(19);
  test_floats_dp_SigmaIn(20) <= test_floats_cp_LambdaOut(20);
  test_floats_dp_SigmaIn(21) <= test_floats_cp_LambdaOut(21);
  test_floats_dp_SigmaIn(22) <= test_floats_cp_LambdaOut(22);
  test_floats_dp_SigmaIn(23) <= test_floats_cp_LambdaOut(23);
  test_floats_dp_SigmaIn(24) <= test_floats_cp_LambdaOut(24);
  test_floats_dp_SigmaIn(25) <= test_floats_cp_LambdaOut(25);
  test_floats_dp_SigmaIn(26) <= test_floats_cp_LambdaOut(26);
  test_floats_dp_SigmaIn(27) <= test_floats_cp_LambdaOut(27);
  test_floats_dp_SigmaIn(28) <= test_floats_cp_LambdaOut(28);
  test_floats_dp_SigmaIn(29) <= test_floats_cp_LambdaOut(29);
  test_floats_dp_SigmaIn(30) <= test_floats_cp_LambdaOut(30);
  test_floats_dp_SigmaIn(31) <= test_floats_cp_LambdaOut(31);
  test_floats_dp_SigmaIn(32) <= test_floats_cp_LambdaOut(32);
  test_floats_dp_SigmaIn(33) <= test_floats_cp_LambdaOut(33);
  test_floats_dp_SigmaIn(34) <= test_floats_cp_LambdaOut(34);
  test_floats_dp_SigmaIn(35) <= test_floats_cp_LambdaOut(35);
  test_floats_dp_SigmaIn(36) <= test_floats_cp_LambdaOut(36);
  test_floats_dp_SigmaIn(37) <= test_floats_cp_LambdaOut(37);
  test_floats_dp_SigmaIn(38) <= test_floats_cp_LambdaOut(38);
  test_floats_dp_SigmaIn(39) <= test_floats_cp_LambdaOut(39);
  test_floats_dp_SigmaIn(40) <= test_floats_cp_LambdaOut(40);
  test_floats_dp_SigmaIn(41) <= test_floats_cp_LambdaOut(41);
  test_floats_dp_SigmaIn(42) <= test_floats_cp_LambdaOut(42);
  test_floats_dp_SigmaIn(43) <= test_floats_cp_LambdaOut(43);
  test_floats_dp_SigmaIn(44) <= test_floats_cp_LambdaOut(44);
  test_floats_dp_SigmaIn(45) <= test_floats_cp_LambdaOut(45);
  test_floats_dp_SigmaIn(46) <= test_floats_cp_LambdaOut(46);
  test_floats_dp_SigmaIn(47) <= test_floats_cp_LambdaOut(47);
  test_floats_dp_SigmaIn(48) <= test_floats_cp_LambdaOut(48);
  test_floats_dp_SigmaIn(49) <= test_floats_cp_LambdaOut(49);
  test_floats_dp_SigmaIn(50) <= test_floats_cp_LambdaOut(50);
  test_floats_dp_SigmaIn(51) <= test_floats_cp_LambdaOut(51);
  test_floats_dp_SigmaIn(52) <= test_floats_cp_LambdaOut(52);
  test_floats_dp_SigmaIn(53) <= test_floats_cp_LambdaOut(53);
  test_floats_dp_SigmaIn(54) <= test_floats_cp_LambdaOut(54);
  test_floats_dp_SigmaIn(55) <= test_floats_cp_LambdaOut(55);
  test_floats_dp_SigmaIn(56) <= test_floats_cp_LambdaOut(56);
  test_floats_dp_SigmaIn(57) <= test_floats_cp_LambdaOut(57);
  test_floats_dp_SigmaIn(58) <= test_floats_cp_LambdaOut(58);
  test_floats_dp_SigmaIn(59) <= test_floats_cp_LambdaOut(59);
  test_floats_dp_SigmaIn(60) <= test_floats_cp_LambdaOut(60);
  test_floats_dp_SigmaIn(61) <= test_floats_cp_LambdaOut(61);
  test_floats_dp_SigmaIn(62) <= test_floats_cp_LambdaOut(62);
  test_floats_dp_SigmaIn(63) <= test_floats_cp_LambdaOut(63);
  test_floats_dp_SigmaIn(64) <= test_floats_cp_LambdaOut(64);
  test_floats_dp_SigmaIn(65) <= test_floats_cp_LambdaOut(65);
  test_floats_dp_SigmaIn(66) <= test_floats_cp_LambdaOut(66);
  test_floats_dp_SigmaIn(67) <= test_floats_cp_LambdaOut(67);
  test_floats_dp_SigmaIn(68) <= test_floats_cp_LambdaOut(68);
  test_floats_dp_SigmaIn(69) <= test_floats_cp_LambdaOut(69);
  test_floats_dp_SigmaIn(70) <= test_floats_cp_LambdaOut(70);
  test_floats_dp_SigmaIn(71) <= test_floats_cp_LambdaOut(71);
  test_floats_dp_SigmaIn(72) <= test_floats_cp_LambdaOut(72);
  test_floats_dp_SigmaIn(73) <= test_floats_cp_LambdaOut(73);
  test_floats_dp_SigmaIn(74) <= test_floats_cp_LambdaOut(74);
  test_floats_dp_SigmaIn(75) <= test_floats_cp_LambdaOut(75);
  test_floats_dp_SigmaIn(76) <= test_floats_cp_LambdaOut(76);
  test_floats_dp_SigmaIn(77) <= test_floats_cp_LambdaOut(77);
  test_floats_dp_SigmaIn(78) <= test_floats_cp_LambdaOut(78);
  test_floats_dp_SigmaIn(79) <= test_floats_cp_LambdaOut(79);
  test_floats_dp_SigmaIn(80) <= test_floats_cp_LambdaOut(80);
  test_floats_dp_SigmaIn(81) <= test_floats_cp_LambdaOut(81);
  test_floats_dp_SigmaIn(82) <= test_floats_cp_LambdaOut(82);
  test_floats_dp_SigmaIn(83) <= test_floats_cp_LambdaOut(83);
  test_floats_dp_SigmaIn(84) <= test_floats_cp_LambdaOut(84);
  test_floats_dp_SigmaIn(85) <= test_floats_cp_LambdaOut(85);
  test_floats_dp_SigmaIn(86) <= test_floats_cp_LambdaOut(86);
  test_floats_dp_SigmaIn(87) <= test_floats_cp_LambdaOut(87);
  test_floats_dp_SigmaIn(88) <= test_floats_cp_LambdaOut(88);
  test_floats_dp_SigmaIn(89) <= test_floats_cp_LambdaOut(89);
  test_floats_dp_SigmaIn(90) <= test_floats_cp_LambdaOut(90);
  test_floats_dp_SigmaIn(91) <= test_floats_cp_LambdaOut(91);
  test_floats_dp_SigmaIn(92) <= test_floats_cp_LambdaOut(92);
  test_floats_dp_SigmaIn(93) <= test_floats_cp_LambdaOut(93);
  test_floats_dp_SigmaIn(94) <= test_floats_cp_LambdaOut(94);
  test_floats_dp_SigmaIn(95) <= test_floats_cp_LambdaOut(95);
  test_floats_dp_SigmaIn(96) <= test_floats_cp_LambdaOut(96);
  test_floats_dp_SigmaIn(97) <= test_floats_cp_LambdaOut(97);
  test_floats_dp_SigmaIn(98) <= test_floats_cp_LambdaOut(98);
  test_floats_dp_SigmaIn(99) <= test_floats_cp_LambdaOut(99);
  test_floats_dp_SigmaIn(100) <= test_floats_cp_LambdaOut(100);
  test_floats_dp_SigmaIn(101) <= test_floats_cp_LambdaOut(101);
  test_floats_dp_SigmaIn(102) <= test_floats_cp_LambdaOut(102);
  test_floats_dp_SigmaIn(103) <= test_floats_cp_LambdaOut(103);
  test_floats_dp_SigmaIn(104) <= test_floats_cp_LambdaOut(104);
  test_floats_dp_SigmaIn(105) <= test_floats_cp_LambdaOut(105);
  test_floats_dp_SigmaIn(106) <= test_floats_cp_LambdaOut(106);
  test_floats_dp_SigmaIn(107) <= test_floats_cp_LambdaOut(107);
  test_floats_dp_SigmaIn(108) <= test_floats_cp_LambdaOut(108);
  test_floats_dp_SigmaIn(109) <= test_floats_cp_LambdaOut(109);
  test_floats_dp_SigmaIn(110) <= test_floats_cp_LambdaOut(110);
  test_floats_dp_SigmaIn(111) <= test_floats_cp_LambdaOut(111);
  test_floats_dp_SigmaIn(112) <= test_floats_cp_LambdaOut(112);
  test_floats_dp_SigmaIn(113) <= test_floats_cp_LambdaOut(113);
  test_floats_dp_SigmaIn(114) <= test_floats_cp_LambdaOut(114);
  test_floats_dp_SigmaIn(115) <= test_floats_cp_LambdaOut(115);
  test_floats_dp_SigmaIn(116) <= test_floats_cp_LambdaOut(116);
  test_floats_dp_SigmaIn(117) <= test_floats_cp_LambdaOut(117);
  test_floats_dp_SigmaIn(118) <= test_floats_cp_LambdaOut(118);
  test_floats_dp_SigmaIn(119) <= test_floats_cp_LambdaOut(119);
  test_floats_dp_SigmaIn(120) <= test_floats_cp_LambdaOut(120);
  test_floats_dp_SigmaIn(121) <= test_floats_cp_LambdaOut(121);
  test_floats_dp_SigmaIn(122) <= test_floats_cp_LambdaOut(122);
  test_floats_dp_SigmaIn(123) <= test_floats_cp_LambdaOut(123);
  test_floats_dp_SigmaIn(124) <= test_floats_cp_LambdaOut(124);
  test_floats_dp_SigmaIn(125) <= test_floats_cp_LambdaOut(125);
  test_floats_dp_SigmaIn(126) <= test_floats_cp_LambdaOut(126);
  test_floats_dp_SigmaIn(127) <= test_floats_cp_LambdaOut(127);
  test_floats_dp_SigmaIn(128) <= test_floats_cp_LambdaOut(128);
  test_floats_dp_SigmaIn(129) <= test_floats_cp_LambdaOut(129);
  test_floats_dp_SigmaIn(130) <= test_floats_cp_LambdaOut(130);
  test_floats_dp_SigmaIn(131) <= test_floats_cp_LambdaOut(131);
  test_floats_dp_SigmaIn(132) <= test_floats_cp_LambdaOut(132);
  test_floats_dp_SigmaIn(133) <= test_floats_cp_LambdaOut(133);
  test_floats_dp_SigmaIn(134) <= test_floats_cp_LambdaOut(134);
  test_floats_dp_SigmaIn(135) <= test_floats_cp_LambdaOut(135);
  test_floats_dp_SigmaIn(136) <= test_floats_cp_LambdaOut(136);
  test_floats_dp_SigmaIn(137) <= test_floats_cp_LambdaOut(137);
  test_floats_dp_SigmaIn(138) <= test_floats_cp_LambdaOut(138);
  test_floats_dp_SigmaIn(139) <= test_floats_cp_LambdaOut(139);
  test_floats_dp_SigmaIn(140) <= test_floats_cp_LambdaOut(140);
  test_floats_dp_SigmaIn(141) <= test_floats_cp_LambdaOut(141);
  test_floats_dp_SigmaIn(142) <= test_floats_cp_LambdaOut(142);
  test_floats_dp_SigmaIn(143) <= test_floats_cp_LambdaOut(143);
  test_floats_dp_SigmaIn(144) <= test_floats_cp_LambdaOut(144);
  test_floats_dp_SigmaIn(145) <= test_floats_cp_LambdaOut(145);
  test_floats_dp_SigmaIn(146) <= test_floats_cp_LambdaOut(146);
  test_floats_dp_SigmaIn(147) <= test_floats_cp_LambdaOut(147);
  test_floats_dp_SigmaIn(148) <= test_floats_cp_LambdaOut(148);
  test_floats_dp_SigmaIn(149) <= test_floats_cp_LambdaOut(149);
  test_floats_dp_SigmaIn(150) <= test_floats_cp_LambdaOut(150);
  test_floats_dp_SigmaIn(151) <= test_floats_cp_LambdaOut(151);
  test_floats_dp_SigmaIn(152) <= test_floats_cp_LambdaOut(152);
  test_floats_dp_SigmaIn(153) <= test_floats_cp_LambdaOut(153);
  test_floats_dp_SigmaIn(154) <= test_floats_cp_LambdaOut(154);
  test_floats_dp_SigmaIn(155) <= test_floats_cp_LambdaOut(155);
  test_floats_dp_SigmaIn(156) <= test_floats_cp_LambdaOut(156);
  test_floats_dp_SigmaIn(157) <= test_floats_cp_LambdaOut(157);
  test_floats_dp_SigmaIn(158) <= test_floats_cp_LambdaOut(158);
  test_floats_dp_SigmaIn(159) <= test_floats_cp_LambdaOut(159);
  test_floats_dp_SigmaIn(160) <= test_floats_cp_LambdaOut(160);
  test_floats_dp_SigmaIn(161) <= test_floats_cp_LambdaOut(161);
  test_floats_dp_SigmaIn(162) <= test_floats_cp_LambdaOut(162);
  test_floats_dp_SigmaIn(163) <= test_floats_cp_LambdaOut(163);
  test_floats_dp_SigmaIn(164) <= test_floats_cp_LambdaOut(164);
  test_floats_dp_SigmaIn(165) <= test_floats_cp_LambdaOut(165);
  test_floats_dp_SigmaIn(166) <= test_floats_cp_LambdaOut(166);
  test_floats_dp_SigmaIn(167) <= test_floats_cp_LambdaOut(167);
  test_floats_dp_SigmaIn(168) <= test_floats_cp_LambdaOut(168);
  test_floats_dp_SigmaIn(169) <= test_floats_cp_LambdaOut(169);
  test_floats_dp_SigmaIn(170) <= test_floats_cp_LambdaOut(170);
  test_floats_dp_SigmaIn(171) <= test_floats_cp_LambdaOut(171);
  test_floats_dp_SigmaIn(172) <= test_floats_cp_LambdaOut(172);
  test_floats_dp_SigmaIn(173) <= test_floats_cp_LambdaOut(173);
  test_floats_dp_SigmaIn(174) <= test_floats_cp_LambdaOut(174);
  test_floats_dp_SigmaIn(175) <= test_floats_cp_LambdaOut(175);
  test_floats_dp_SigmaIn(176) <= test_floats_cp_LambdaOut(176);
  test_floats_dp_SigmaIn(177) <= test_floats_cp_LambdaOut(177);
  test_floats_dp_SigmaIn(178) <= test_floats_cp_LambdaOut(178);
  test_floats_dp_SigmaIn(179) <= test_floats_cp_LambdaOut(179);
  test_floats_dp_SigmaIn(180) <= test_floats_cp_LambdaOut(180);
  test_floats_dp_SigmaIn(181) <= test_floats_cp_LambdaOut(181);
  test_floats_dp_SigmaIn(182) <= test_floats_cp_LambdaOut(182);
  test_floats_dp_SigmaIn(183) <= test_floats_cp_LambdaOut(183);
  test_floats_dp_SigmaIn(184) <= test_floats_cp_LambdaOut(184);
  test_floats_dp_SigmaIn(185) <= test_floats_cp_LambdaOut(185);
  test_floats_dp_SigmaIn(186) <= test_floats_cp_LambdaOut(186);
  test_floats_dp_SigmaIn(187) <= test_floats_cp_LambdaOut(187);
  test_floats_dp_SigmaIn(188) <= test_floats_cp_LambdaOut(188);
  test_floats_dp_SigmaIn(189) <= test_floats_cp_LambdaOut(189);
  test_floats_dp_SigmaIn(190) <= test_floats_cp_LambdaOut(190);
  test_floats_dp_SigmaIn(191) <= test_floats_cp_LambdaOut(191);
  test_floats_dp_SigmaIn(192) <= test_floats_cp_LambdaOut(192);
  test_floats_dp_SigmaIn(193) <= test_floats_cp_LambdaOut(193);
  test_floats_dp_SigmaIn(194) <= test_floats_cp_LambdaOut(194);
  test_floats_dp_SigmaIn(195) <= test_floats_cp_LambdaOut(195);
  test_floats_dp_SigmaIn(196) <= test_floats_cp_LambdaOut(196);
  test_floats_dp_SigmaIn(197) <= test_floats_cp_LambdaOut(197);
  test_floats_dp_SigmaIn(198) <= test_floats_cp_LambdaOut(198);
  test_floats_dp_SigmaIn(199) <= test_floats_cp_LambdaOut(199);
  test_floats_dp_SigmaIn(200) <= test_floats_cp_LambdaOut(200);
  test_floats_dp_SigmaIn(201) <= test_floats_cp_LambdaOut(201);
  test_floats_dp_SigmaIn(202) <= test_floats_cp_LambdaOut(202);
  test_floats_dp_SigmaIn(203) <= test_floats_cp_LambdaOut(203);
  test_floats_dp_SigmaIn(204) <= test_floats_cp_LambdaOut(204);
  test_floats_dp_SigmaIn(205) <= test_floats_cp_LambdaOut(205);
  test_floats_dp_SigmaIn(206) <= test_floats_cp_LambdaOut(206);
  test_floats_dp_SigmaIn(207) <= test_floats_cp_LambdaOut(207);
  test_floats_dp_SigmaIn(208) <= test_floats_cp_LambdaOut(208);
  test_floats_dp_SigmaIn(209) <= test_floats_cp_LambdaOut(209);
  test_floats_dp_SigmaIn(210) <= test_floats_cp_LambdaOut(210);
  test_floats_dp_SigmaIn(211) <= test_floats_cp_LambdaOut(211);
  test_floats_dp_SigmaIn(212) <= test_floats_cp_LambdaOut(212);
  test_floats_dp_SigmaIn(213) <= test_floats_cp_LambdaOut(213);
  test_floats_dp_SigmaIn(214) <= test_floats_cp_LambdaOut(214);
  test_floats_dp_SigmaIn(215) <= test_floats_cp_LambdaOut(215);
  test_floats_dp_SigmaIn(216) <= test_floats_cp_LambdaOut(216);
  test_floats_dp_SigmaIn(217) <= test_floats_cp_LambdaOut(217);
  test_floats_dp_SigmaIn(218) <= test_floats_cp_LambdaOut(218);
  test_floats_dp_SigmaIn(219) <= test_floats_cp_LambdaOut(219);
  test_floats_dp_SigmaIn(220) <= test_floats_cp_LambdaOut(220);
  test_floats_dp_SigmaIn(221) <= test_floats_cp_LambdaOut(221);
  test_floats_dp_SigmaIn(222) <= test_floats_cp_LambdaOut(222);
  test_floats_dp_SigmaIn(223) <= test_floats_cp_LambdaOut(223);
  test_floats_dp_SigmaIn(224) <= test_floats_cp_LambdaOut(224);
  test_floats_dp_SigmaIn(225) <= test_floats_cp_LambdaOut(225);
  test_floats_dp_SigmaIn(226) <= test_floats_cp_LambdaOut(226);
  test_floats_dp_SigmaIn(227) <= test_floats_cp_LambdaOut(227);
  test_floats_dp_SigmaIn(228) <= test_floats_cp_LambdaOut(228);
  test_floats_dp_SigmaIn(229) <= test_floats_cp_LambdaOut(229);
  test_floats_dp_SigmaIn(230) <= test_floats_cp_LambdaOut(230);
  test_floats_dp_SigmaIn(231) <= test_floats_cp_LambdaOut(231);
  test_floats_dp_SigmaIn(232) <= test_floats_cp_LambdaOut(232);
  test_floats_dp_SigmaIn(233) <= test_floats_cp_LambdaOut(233);
  test_floats_dp_SigmaIn(234) <= test_floats_cp_LambdaOut(234);
  test_floats_dp_SigmaIn(235) <= test_floats_cp_LambdaOut(235);
  test_floats_dp_SigmaIn(236) <= test_floats_cp_LambdaOut(236);
  test_floats_dp_SigmaIn(237) <= test_floats_cp_LambdaOut(237);
  test_floats_dp_SigmaIn(238) <= test_floats_cp_LambdaOut(238);
  test_floats_dp_SigmaIn(239) <= test_floats_cp_LambdaOut(239);
  test_floats_dp_SigmaIn(240) <= test_floats_cp_LambdaOut(240);
  test_floats_dp_SigmaIn(241) <= test_floats_cp_LambdaOut(241);
  test_floats_dp_SigmaIn(242) <= test_floats_cp_LambdaOut(242);
  test_floats_dp_SigmaIn(243) <= test_floats_cp_LambdaOut(243);
  test_floats_dp_SigmaIn(244) <= test_floats_cp_LambdaOut(244);
  test_floats_dp_SigmaIn(245) <= test_floats_cp_LambdaOut(245);
  test_floats_dp_SigmaIn(246) <= test_floats_cp_LambdaOut(246);
  test_floats_dp_SigmaIn(247) <= test_floats_cp_LambdaOut(247);
  test_floats_dp_SigmaIn(248) <= test_floats_cp_LambdaOut(248);
  test_floats_dp_SigmaIn(249) <= test_floats_cp_LambdaOut(249);
  test_floats_dp_SigmaIn(250) <= test_floats_cp_LambdaOut(250);
  test_floats_dp_SigmaIn(251) <= test_floats_cp_LambdaOut(251);
  test_floats_dp_SigmaIn(252) <= test_floats_cp_LambdaOut(252);
  test_floats_dp_SigmaIn(253) <= test_floats_cp_LambdaOut(253);
  test_floats_dp_SigmaIn(254) <= test_floats_cp_LambdaOut(254);
  test_floats_dp_SigmaIn(255) <= test_floats_cp_LambdaOut(255);
  test_floats_dp_SigmaIn(256) <= test_floats_cp_LambdaOut(256);
  test_floats_dp_SigmaIn(257) <= test_floats_cp_LambdaOut(257);
  test_floats_dp_SigmaIn(258) <= test_floats_cp_LambdaOut(258);
  test_floats_dp_SigmaIn(259) <= test_floats_cp_LambdaOut(259);
  test_floats_dp_SigmaIn(260) <= test_floats_cp_LambdaOut(260);
  test_floats_dp_SigmaIn(261) <= test_floats_cp_LambdaOut(261);
  test_floats_dp_SigmaIn(262) <= test_floats_cp_LambdaOut(262);
  test_floats_dp_SigmaIn(263) <= test_floats_cp_LambdaOut(263);
  test_floats_dp_SigmaIn(264) <= test_floats_cp_LambdaOut(264);
  test_floats_dp_SigmaIn(265) <= test_floats_cp_LambdaOut(265);
  test_floats_dp_SigmaIn(266) <= test_floats_cp_LambdaOut(266);
  test_floats_dp_SigmaIn(267) <= test_floats_cp_LambdaOut(267);
  test_floats_dp_SigmaIn(268) <= test_floats_cp_LambdaOut(268);
  test_floats_dp_SigmaIn(269) <= test_floats_cp_LambdaOut(269);
  test_floats_dp_SigmaIn(270) <= test_floats_cp_LambdaOut(270);
  test_floats_dp_SigmaIn(271) <= test_floats_cp_LambdaOut(271);
  test_floats_dp_SigmaIn(272) <= test_floats_cp_LambdaOut(272);
  test_floats_dp_SigmaIn(273) <= test_floats_cp_LambdaOut(273);
  test_floats_dp_SigmaIn(274) <= test_floats_cp_LambdaOut(274);
  test_floats_dp_SigmaIn(275) <= test_floats_cp_LambdaOut(275);
  test_floats_dp_SigmaIn(276) <= test_floats_cp_LambdaOut(276);
  test_floats_dp_SigmaIn(277) <= test_floats_cp_LambdaOut(277);
  test_floats_dp_SigmaIn(278) <= test_floats_cp_LambdaOut(278);
  test_floats_dp_SigmaIn(279) <= test_floats_cp_LambdaOut(279);
  test_floats_dp_SigmaIn(280) <= test_floats_cp_LambdaOut(280);
  test_floats_dp_SigmaIn(281) <= test_floats_cp_LambdaOut(281);
  test_floats_dp_SigmaIn(282) <= test_floats_cp_LambdaOut(282);
  test_floats_dp_SigmaIn(283) <= test_floats_cp_LambdaOut(283);
  test_floats_dp_SigmaIn(284) <= test_floats_cp_LambdaOut(284);
  test_floats_dp_SigmaIn(285) <= test_floats_cp_LambdaOut(285);
  test_floats_dp_SigmaIn(286) <= test_floats_cp_LambdaOut(286);
  test_floats_dp_SigmaIn(287) <= test_floats_cp_LambdaOut(287);
  test_floats_dp_SigmaIn(288) <= test_floats_cp_LambdaOut(288);
  test_floats_dp_SigmaIn(289) <= test_floats_cp_LambdaOut(289);
  test_floats_dp_SigmaIn(290) <= test_floats_cp_LambdaOut(290);
  test_floats_dp_SigmaIn(291) <= test_floats_cp_LambdaOut(291);
  test_floats_dp_SigmaIn(292) <= test_floats_cp_LambdaOut(292);
  test_floats_dp_SigmaIn(293) <= test_floats_cp_LambdaOut(293);
  test_floats_dp_SigmaIn(294) <= test_floats_cp_LambdaOut(294);
  test_floats_dp_SigmaIn(295) <= test_floats_cp_LambdaOut(295);
  test_floats_dp_SigmaIn(296) <= test_floats_cp_LambdaOut(296);
  test_floats_dp_SigmaIn(297) <= test_floats_cp_LambdaOut(297);
  test_floats_dp_SigmaIn(298) <= test_floats_cp_LambdaOut(298);
  test_floats_dp_SigmaIn(299) <= test_floats_cp_LambdaOut(299);
  test_floats_dp_SigmaIn(300) <= test_floats_cp_LambdaOut(300);
  test_floats_dp_SigmaIn(301) <= test_floats_cp_LambdaOut(301);
  test_floats_dp_SigmaIn(302) <= test_floats_cp_LambdaOut(302);
  test_floats_dp_SigmaIn(303) <= test_floats_cp_LambdaOut(303);
  test_floats_dp_SigmaIn(304) <= test_floats_cp_LambdaOut(304);
  test_floats_dp_SigmaIn(305) <= test_floats_cp_LambdaOut(305);
  test_floats_dp_SigmaIn(306) <= test_floats_cp_LambdaOut(306);
  test_floats_dp_SigmaIn(307) <= test_floats_cp_LambdaOut(307);
  test_floats_dp_SigmaIn(308) <= test_floats_cp_LambdaOut(308);
  test_floats_dp_SigmaIn(309) <= test_floats_cp_LambdaOut(309);
  test_floats_dp_SigmaIn(310) <= test_floats_cp_LambdaOut(310);
  test_floats_dp_SigmaIn(311) <= test_floats_cp_LambdaOut(311);
  test_floats_dp_SigmaIn(312) <= test_floats_cp_LambdaOut(312);
  test_floats_dp_SigmaIn(313) <= test_floats_cp_LambdaOut(313);
  test_floats_dp_SigmaIn(314) <= test_floats_cp_LambdaOut(314);
  test_floats_dp_SigmaIn(315) <= test_floats_cp_LambdaOut(315);
  test_floats_dp_SigmaIn(316) <= test_floats_cp_LambdaOut(316);
  test_floats_dp_SigmaIn(317) <= test_floats_cp_LambdaOut(317);
  test_floats_dp_SigmaIn(318) <= test_floats_cp_LambdaOut(318);
  test_floats_dp_SigmaIn(319) <= test_floats_cp_LambdaOut(319);
  test_floats_dp_SigmaIn(320) <= test_floats_cp_LambdaOut(320);
  test_floats_dp_SigmaIn(321) <= test_floats_cp_LambdaOut(321);
  test_floats_dp_SigmaIn(322) <= test_floats_cp_LambdaOut(322);
  test_floats_dp_SigmaIn(323) <= test_floats_cp_LambdaOut(323);
end default_arch;