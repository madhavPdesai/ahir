-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package vc_system_package is -- 
  constant GV_15_base_address : std_logic_vector(8 downto 0) := "000000000";
  constant GV_16_base_address : std_logic_vector(4 downto 0) := "00000";
  constant ahir_heap_base_address : std_logic_vector(13 downto 0) := "00000000000000";
  constant click_bc_iNtErNal_x_ZZN14LinearIPLookup4pushEiP6PacketE10complained_base_address : std_logic_vector(0 downto 0) := "0";
  constant free_queue_ram_base_address : std_logic_vector(15 downto 0) := "0000000000000000";
  constant mempool_base_address : std_logic_vector(0 downto 0) := "0";
  -- 
end package vc_system_package;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity GV_15_initializer_in_click_bc is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity GV_15_initializer_in_click_bc;
architecture Default of GV_15_initializer_in_click_bc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal GV_15_initializer_in_click_bc_CP_0_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_176_gather_scatter_req_0 : boolean;
  signal array_obj_ref_176_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_241_store_0_ack_0 : boolean;
  signal array_obj_ref_241_store_0_req_1 : boolean;
  signal array_obj_ref_241_store_0_ack_1 : boolean;
  signal array_obj_ref_176_store_0_req_0 : boolean;
  signal array_obj_ref_176_store_0_ack_0 : boolean;
  signal array_obj_ref_176_store_0_req_1 : boolean;
  signal array_obj_ref_176_store_0_ack_1 : boolean;
  signal array_obj_ref_185_gather_scatter_req_0 : boolean;
  signal array_obj_ref_185_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_185_store_0_req_0 : boolean;
  signal array_obj_ref_185_store_0_ack_0 : boolean;
  signal array_obj_ref_185_store_0_req_1 : boolean;
  signal array_obj_ref_185_store_0_ack_1 : boolean;
  signal array_obj_ref_192_gather_scatter_req_0 : boolean;
  signal array_obj_ref_192_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_192_store_0_req_0 : boolean;
  signal array_obj_ref_192_store_0_ack_0 : boolean;
  signal array_obj_ref_192_store_0_req_1 : boolean;
  signal array_obj_ref_192_store_0_ack_1 : boolean;
  signal array_obj_ref_199_gather_scatter_req_0 : boolean;
  signal array_obj_ref_199_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_199_store_0_req_0 : boolean;
  signal array_obj_ref_199_store_0_ack_0 : boolean;
  signal array_obj_ref_199_store_0_req_1 : boolean;
  signal array_obj_ref_199_store_0_ack_1 : boolean;
  signal array_obj_ref_206_gather_scatter_req_0 : boolean;
  signal array_obj_ref_206_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_0 : boolean;
  signal array_obj_ref_206_store_0_ack_0 : boolean;
  signal array_obj_ref_206_store_0_req_1 : boolean;
  signal array_obj_ref_206_store_0_ack_1 : boolean;
  signal array_obj_ref_213_gather_scatter_req_0 : boolean;
  signal array_obj_ref_213_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_213_store_0_req_0 : boolean;
  signal array_obj_ref_213_store_0_ack_0 : boolean;
  signal array_obj_ref_213_store_0_req_1 : boolean;
  signal array_obj_ref_213_store_0_ack_1 : boolean;
  signal array_obj_ref_220_gather_scatter_req_0 : boolean;
  signal array_obj_ref_220_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_220_store_0_req_0 : boolean;
  signal array_obj_ref_220_store_0_ack_0 : boolean;
  signal array_obj_ref_220_store_0_req_1 : boolean;
  signal array_obj_ref_220_store_0_ack_1 : boolean;
  signal array_obj_ref_227_gather_scatter_req_0 : boolean;
  signal array_obj_ref_227_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_227_store_0_req_0 : boolean;
  signal array_obj_ref_227_store_0_ack_0 : boolean;
  signal array_obj_ref_227_store_0_req_1 : boolean;
  signal array_obj_ref_227_store_0_ack_1 : boolean;
  signal array_obj_ref_234_gather_scatter_req_0 : boolean;
  signal array_obj_ref_234_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_0 : boolean;
  signal array_obj_ref_234_store_0_ack_0 : boolean;
  signal array_obj_ref_234_store_0_req_1 : boolean;
  signal array_obj_ref_234_store_0_ack_1 : boolean;
  signal array_obj_ref_241_gather_scatter_req_0 : boolean;
  signal array_obj_ref_241_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_241_store_0_req_0 : boolean;
  signal array_obj_ref_248_gather_scatter_req_0 : boolean;
  signal array_obj_ref_248_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_248_store_0_req_0 : boolean;
  signal array_obj_ref_248_store_0_ack_0 : boolean;
  signal array_obj_ref_248_store_0_req_1 : boolean;
  signal array_obj_ref_248_store_0_ack_1 : boolean;
  signal array_obj_ref_255_gather_scatter_req_0 : boolean;
  signal array_obj_ref_255_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_255_store_0_req_0 : boolean;
  signal array_obj_ref_255_store_0_ack_0 : boolean;
  signal array_obj_ref_255_store_0_req_1 : boolean;
  signal array_obj_ref_255_store_0_ack_1 : boolean;
  signal array_obj_ref_262_gather_scatter_req_0 : boolean;
  signal array_obj_ref_262_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_0 : boolean;
  signal array_obj_ref_262_store_0_ack_0 : boolean;
  signal array_obj_ref_262_store_0_req_1 : boolean;
  signal array_obj_ref_262_store_0_ack_1 : boolean;
  signal array_obj_ref_269_gather_scatter_req_0 : boolean;
  signal array_obj_ref_269_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_269_store_0_req_0 : boolean;
  signal array_obj_ref_269_store_0_ack_0 : boolean;
  signal array_obj_ref_269_store_0_req_1 : boolean;
  signal array_obj_ref_269_store_0_ack_1 : boolean;
  signal array_obj_ref_276_gather_scatter_req_0 : boolean;
  signal array_obj_ref_276_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_0 : boolean;
  signal array_obj_ref_276_store_0_ack_0 : boolean;
  signal array_obj_ref_276_store_0_req_1 : boolean;
  signal array_obj_ref_276_store_0_ack_1 : boolean;
  signal array_obj_ref_283_gather_scatter_req_0 : boolean;
  signal array_obj_ref_283_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_283_store_0_req_0 : boolean;
  signal array_obj_ref_283_store_0_ack_0 : boolean;
  signal array_obj_ref_283_store_0_req_1 : boolean;
  signal array_obj_ref_283_store_0_ack_1 : boolean;
  signal array_obj_ref_290_gather_scatter_req_0 : boolean;
  signal array_obj_ref_290_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_290_store_0_req_0 : boolean;
  signal array_obj_ref_290_store_0_ack_0 : boolean;
  signal array_obj_ref_290_store_0_req_1 : boolean;
  signal array_obj_ref_290_store_0_ack_1 : boolean;
  signal array_obj_ref_297_gather_scatter_req_0 : boolean;
  signal array_obj_ref_297_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_297_store_0_req_0 : boolean;
  signal array_obj_ref_297_store_0_ack_0 : boolean;
  signal array_obj_ref_297_store_0_req_1 : boolean;
  signal array_obj_ref_297_store_0_ack_1 : boolean;
  signal array_obj_ref_304_gather_scatter_req_0 : boolean;
  signal array_obj_ref_304_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_0 : boolean;
  signal array_obj_ref_304_store_0_ack_0 : boolean;
  signal array_obj_ref_304_store_0_req_1 : boolean;
  signal array_obj_ref_304_store_0_ack_1 : boolean;
  signal array_obj_ref_311_gather_scatter_req_0 : boolean;
  signal array_obj_ref_311_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_311_store_0_req_0 : boolean;
  signal array_obj_ref_311_store_0_ack_0 : boolean;
  signal array_obj_ref_311_store_0_req_1 : boolean;
  signal array_obj_ref_311_store_0_ack_1 : boolean;
  signal array_obj_ref_318_gather_scatter_req_0 : boolean;
  signal array_obj_ref_318_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_0 : boolean;
  signal array_obj_ref_318_store_0_ack_0 : boolean;
  signal array_obj_ref_318_store_0_req_1 : boolean;
  signal array_obj_ref_318_store_0_ack_1 : boolean;
  signal array_obj_ref_325_gather_scatter_req_0 : boolean;
  signal array_obj_ref_325_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_325_store_0_req_0 : boolean;
  signal array_obj_ref_325_store_0_ack_0 : boolean;
  signal array_obj_ref_325_store_0_req_1 : boolean;
  signal array_obj_ref_325_store_0_ack_1 : boolean;
  signal array_obj_ref_332_gather_scatter_req_0 : boolean;
  signal array_obj_ref_332_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_332_store_0_req_0 : boolean;
  signal array_obj_ref_332_store_0_ack_0 : boolean;
  signal array_obj_ref_332_store_0_req_1 : boolean;
  signal array_obj_ref_332_store_0_ack_1 : boolean;
  signal array_obj_ref_339_gather_scatter_req_0 : boolean;
  signal array_obj_ref_339_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_339_store_0_req_0 : boolean;
  signal array_obj_ref_339_store_0_ack_0 : boolean;
  signal array_obj_ref_339_store_0_req_1 : boolean;
  signal array_obj_ref_339_store_0_ack_1 : boolean;
  signal array_obj_ref_346_gather_scatter_req_0 : boolean;
  signal array_obj_ref_346_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_0 : boolean;
  signal array_obj_ref_346_store_0_ack_0 : boolean;
  signal array_obj_ref_346_store_0_req_1 : boolean;
  signal array_obj_ref_346_store_0_ack_1 : boolean;
  signal array_obj_ref_353_gather_scatter_req_0 : boolean;
  signal array_obj_ref_353_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_353_store_0_req_0 : boolean;
  signal array_obj_ref_353_store_0_ack_0 : boolean;
  signal array_obj_ref_353_store_0_req_1 : boolean;
  signal array_obj_ref_353_store_0_ack_1 : boolean;
  signal array_obj_ref_360_gather_scatter_req_0 : boolean;
  signal array_obj_ref_360_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_360_store_0_req_0 : boolean;
  signal array_obj_ref_360_store_0_ack_0 : boolean;
  signal array_obj_ref_360_store_0_req_1 : boolean;
  signal array_obj_ref_360_store_0_ack_1 : boolean;
  signal array_obj_ref_367_gather_scatter_req_0 : boolean;
  signal array_obj_ref_367_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_367_store_0_req_0 : boolean;
  signal array_obj_ref_367_store_0_ack_0 : boolean;
  signal array_obj_ref_367_store_0_req_1 : boolean;
  signal array_obj_ref_367_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  GV_15_initializer_in_click_bc_CP_0: Block -- control-path 
    signal cp_elements: BooleanArray(84 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(84);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(84), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    split_req_12_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => array_obj_ref_176_gather_scatter_req_0); -- 
    split_ack_13_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_gather_scatter_ack_0, ack => cp_elements(1)); -- 
    rr_20_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => array_obj_ref_176_store_0_req_0); -- 
    ra_21_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_store_0_ack_0, ack => cp_elements(2)); -- 
    cr_22_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => array_obj_ref_176_store_0_req_1); -- 
    ca_23_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_176_store_0_ack_1, ack => cp_elements(3)); -- 
    split_req_33_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => array_obj_ref_185_gather_scatter_req_0); -- 
    split_ack_34_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_gather_scatter_ack_0, ack => cp_elements(4)); -- 
    rr_41_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => array_obj_ref_185_store_0_req_0); -- 
    ra_42_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_store_0_ack_0, ack => cp_elements(5)); -- 
    cr_43_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => array_obj_ref_185_store_0_req_1); -- 
    ca_44_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_185_store_0_ack_1, ack => cp_elements(6)); -- 
    split_req_54_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => array_obj_ref_192_gather_scatter_req_0); -- 
    split_ack_55_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_gather_scatter_ack_0, ack => cp_elements(7)); -- 
    rr_62_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => array_obj_ref_192_store_0_req_0); -- 
    ra_63_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_store_0_ack_0, ack => cp_elements(8)); -- 
    cr_64_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => array_obj_ref_192_store_0_req_1); -- 
    ca_65_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_192_store_0_ack_1, ack => cp_elements(9)); -- 
    split_req_75_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => array_obj_ref_199_gather_scatter_req_0); -- 
    split_ack_76_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_83_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => array_obj_ref_199_store_0_req_0); -- 
    ra_84_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_85_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => array_obj_ref_199_store_0_req_1); -- 
    ca_86_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_199_store_0_ack_1, ack => cp_elements(12)); -- 
    split_req_96_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => array_obj_ref_206_gather_scatter_req_0); -- 
    split_ack_97_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => array_obj_ref_206_store_0_req_0); -- 
    ra_105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_store_0_ack_0, ack => cp_elements(14)); -- 
    cr_106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => array_obj_ref_206_store_0_req_1); -- 
    ca_107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_206_store_0_ack_1, ack => cp_elements(15)); -- 
    split_req_117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => array_obj_ref_213_gather_scatter_req_0); -- 
    split_ack_118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_213_store_0_req_0); -- 
    ra_126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_0, ack => cp_elements(17)); -- 
    cr_127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_213_store_0_req_1); -- 
    ca_128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_213_store_0_ack_1, ack => cp_elements(18)); -- 
    split_req_138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_220_gather_scatter_req_0); -- 
    split_ack_139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_gather_scatter_ack_0, ack => cp_elements(19)); -- 
    rr_146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => array_obj_ref_220_store_0_req_0); -- 
    ra_147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_store_0_ack_0, ack => cp_elements(20)); -- 
    cr_148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => array_obj_ref_220_store_0_req_1); -- 
    ca_149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_220_store_0_ack_1, ack => cp_elements(21)); -- 
    split_req_159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_227_gather_scatter_req_0); -- 
    split_ack_160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    rr_167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_227_store_0_req_0); -- 
    ra_168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_store_0_ack_0, ack => cp_elements(23)); -- 
    cr_169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_227_store_0_req_1); -- 
    ca_170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_227_store_0_ack_1, ack => cp_elements(24)); -- 
    split_req_180_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => array_obj_ref_234_gather_scatter_req_0); -- 
    split_ack_181_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    rr_188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => array_obj_ref_234_store_0_req_0); -- 
    ra_189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_store_0_ack_0, ack => cp_elements(26)); -- 
    cr_190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => array_obj_ref_234_store_0_req_1); -- 
    ca_191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_234_store_0_ack_1, ack => cp_elements(27)); -- 
    split_req_201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_241_gather_scatter_req_0); -- 
    split_ack_202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    rr_209_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => array_obj_ref_241_store_0_req_0); -- 
    ra_210_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_store_0_ack_0, ack => cp_elements(29)); -- 
    cr_211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_241_store_0_req_1); -- 
    ca_212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_241_store_0_ack_1, ack => cp_elements(30)); -- 
    split_req_222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_248_gather_scatter_req_0); -- 
    split_ack_223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_gather_scatter_ack_0, ack => cp_elements(31)); -- 
    rr_230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_248_store_0_req_0); -- 
    ra_231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_store_0_ack_0, ack => cp_elements(32)); -- 
    cr_232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_248_store_0_req_1); -- 
    ca_233_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_248_store_0_ack_1, ack => cp_elements(33)); -- 
    split_req_243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_255_gather_scatter_req_0); -- 
    split_ack_244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_gather_scatter_ack_0, ack => cp_elements(34)); -- 
    rr_251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_255_store_0_req_0); -- 
    ra_252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_store_0_ack_0, ack => cp_elements(35)); -- 
    cr_253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_255_store_0_req_1); -- 
    ca_254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_255_store_0_ack_1, ack => cp_elements(36)); -- 
    split_req_264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_262_gather_scatter_req_0); -- 
    split_ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_gather_scatter_ack_0, ack => cp_elements(37)); -- 
    rr_272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_262_store_0_req_0); -- 
    ra_273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_store_0_ack_0, ack => cp_elements(38)); -- 
    cr_274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_262_store_0_req_1); -- 
    ca_275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_262_store_0_ack_1, ack => cp_elements(39)); -- 
    split_req_285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => array_obj_ref_269_gather_scatter_req_0); -- 
    split_ack_286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_gather_scatter_ack_0, ack => cp_elements(40)); -- 
    rr_293_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => array_obj_ref_269_store_0_req_0); -- 
    ra_294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_store_0_ack_0, ack => cp_elements(41)); -- 
    cr_295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => array_obj_ref_269_store_0_req_1); -- 
    ca_296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_269_store_0_ack_1, ack => cp_elements(42)); -- 
    split_req_306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => array_obj_ref_276_gather_scatter_req_0); -- 
    split_ack_307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_gather_scatter_ack_0, ack => cp_elements(43)); -- 
    rr_314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => array_obj_ref_276_store_0_req_0); -- 
    ra_315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_store_0_ack_0, ack => cp_elements(44)); -- 
    cr_316_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => array_obj_ref_276_store_0_req_1); -- 
    ca_317_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_276_store_0_ack_1, ack => cp_elements(45)); -- 
    split_req_327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => array_obj_ref_283_gather_scatter_req_0); -- 
    split_ack_328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_gather_scatter_ack_0, ack => cp_elements(46)); -- 
    rr_335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => array_obj_ref_283_store_0_req_0); -- 
    ra_336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_store_0_ack_0, ack => cp_elements(47)); -- 
    cr_337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => array_obj_ref_283_store_0_req_1); -- 
    ca_338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_283_store_0_ack_1, ack => cp_elements(48)); -- 
    split_req_348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => array_obj_ref_290_gather_scatter_req_0); -- 
    split_ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_gather_scatter_ack_0, ack => cp_elements(49)); -- 
    rr_356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => array_obj_ref_290_store_0_req_0); -- 
    ra_357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_store_0_ack_0, ack => cp_elements(50)); -- 
    cr_358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => array_obj_ref_290_store_0_req_1); -- 
    ca_359_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_290_store_0_ack_1, ack => cp_elements(51)); -- 
    split_req_369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_297_gather_scatter_req_0); -- 
    split_ack_370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_gather_scatter_ack_0, ack => cp_elements(52)); -- 
    rr_377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_297_store_0_req_0); -- 
    ra_378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_store_0_ack_0, ack => cp_elements(53)); -- 
    cr_379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_297_store_0_req_1); -- 
    ca_380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_store_0_ack_1, ack => cp_elements(54)); -- 
    split_req_390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_304_gather_scatter_req_0); -- 
    split_ack_391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_gather_scatter_ack_0, ack => cp_elements(55)); -- 
    rr_398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => array_obj_ref_304_store_0_req_0); -- 
    ra_399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_0, ack => cp_elements(56)); -- 
    cr_400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => array_obj_ref_304_store_0_req_1); -- 
    ca_401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_304_store_0_ack_1, ack => cp_elements(57)); -- 
    split_req_411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => array_obj_ref_311_gather_scatter_req_0); -- 
    split_ack_412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_gather_scatter_ack_0, ack => cp_elements(58)); -- 
    rr_419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => array_obj_ref_311_store_0_req_0); -- 
    ra_420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_store_0_ack_0, ack => cp_elements(59)); -- 
    cr_421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => array_obj_ref_311_store_0_req_1); -- 
    ca_422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_311_store_0_ack_1, ack => cp_elements(60)); -- 
    split_req_432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => array_obj_ref_318_gather_scatter_req_0); -- 
    split_ack_433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_gather_scatter_ack_0, ack => cp_elements(61)); -- 
    rr_440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => array_obj_ref_318_store_0_req_0); -- 
    ra_441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_store_0_ack_0, ack => cp_elements(62)); -- 
    cr_442_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => array_obj_ref_318_store_0_req_1); -- 
    ca_443_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_318_store_0_ack_1, ack => cp_elements(63)); -- 
    split_req_453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => array_obj_ref_325_gather_scatter_req_0); -- 
    split_ack_454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_gather_scatter_ack_0, ack => cp_elements(64)); -- 
    rr_461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => array_obj_ref_325_store_0_req_0); -- 
    ra_462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_store_0_ack_0, ack => cp_elements(65)); -- 
    cr_463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => array_obj_ref_325_store_0_req_1); -- 
    ca_464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_325_store_0_ack_1, ack => cp_elements(66)); -- 
    split_req_474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => array_obj_ref_332_gather_scatter_req_0); -- 
    split_ack_475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_gather_scatter_ack_0, ack => cp_elements(67)); -- 
    rr_482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => array_obj_ref_332_store_0_req_0); -- 
    ra_483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_store_0_ack_0, ack => cp_elements(68)); -- 
    cr_484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => array_obj_ref_332_store_0_req_1); -- 
    ca_485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_332_store_0_ack_1, ack => cp_elements(69)); -- 
    split_req_495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_339_gather_scatter_req_0); -- 
    split_ack_496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_gather_scatter_ack_0, ack => cp_elements(70)); -- 
    rr_503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_339_store_0_req_0); -- 
    ra_504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_store_0_ack_0, ack => cp_elements(71)); -- 
    cr_505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_339_store_0_req_1); -- 
    ca_506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_339_store_0_ack_1, ack => cp_elements(72)); -- 
    split_req_516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_346_gather_scatter_req_0); -- 
    split_ack_517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_gather_scatter_ack_0, ack => cp_elements(73)); -- 
    rr_524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_346_store_0_req_0); -- 
    ra_525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_store_0_ack_0, ack => cp_elements(74)); -- 
    cr_526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_346_store_0_req_1); -- 
    ca_527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_346_store_0_ack_1, ack => cp_elements(75)); -- 
    split_req_537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_353_gather_scatter_req_0); -- 
    split_ack_538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_gather_scatter_ack_0, ack => cp_elements(76)); -- 
    rr_545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => array_obj_ref_353_store_0_req_0); -- 
    ra_546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_store_0_ack_0, ack => cp_elements(77)); -- 
    cr_547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => array_obj_ref_353_store_0_req_1); -- 
    ca_548_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_353_store_0_ack_1, ack => cp_elements(78)); -- 
    split_req_558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => array_obj_ref_360_gather_scatter_req_0); -- 
    split_ack_559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_gather_scatter_ack_0, ack => cp_elements(79)); -- 
    rr_566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => array_obj_ref_360_store_0_req_0); -- 
    ra_567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_store_0_ack_0, ack => cp_elements(80)); -- 
    cr_568_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => array_obj_ref_360_store_0_req_1); -- 
    ca_569_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_360_store_0_ack_1, ack => cp_elements(81)); -- 
    split_req_579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_367_gather_scatter_req_0); -- 
    split_ack_580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_gather_scatter_ack_0, ack => cp_elements(82)); -- 
    rr_587_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_367_store_0_req_0); -- 
    ra_588_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_store_0_ack_0, ack => cp_elements(83)); -- 
    cr_589_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => array_obj_ref_367_store_0_req_1); -- 
    ca_590_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_367_store_0_ack_1, ack => cp_elements(84)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_176_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_176_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_185_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_185_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_192_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_192_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_199_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_199_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_206_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_206_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_213_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_213_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_220_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_220_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_227_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_227_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_234_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_234_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_241_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_241_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_248_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_248_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_255_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_255_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_262_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_262_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_269_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_269_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_276_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_276_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_283_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_283_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_290_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_290_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_297_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_297_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_304_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_304_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_311_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_311_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_318_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_318_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_325_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_325_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_332_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_332_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_339_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_339_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_346_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_346_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_353_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_353_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_360_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_360_word_address_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_367_data_0 : std_logic_vector(7 downto 0);
    signal array_obj_ref_367_word_address_0 : std_logic_vector(8 downto 0);
    signal expr_177_wire_constant : std_logic_vector(7 downto 0);
    signal expr_186_wire_constant : std_logic_vector(7 downto 0);
    signal expr_193_wire_constant : std_logic_vector(7 downto 0);
    signal expr_200_wire_constant : std_logic_vector(7 downto 0);
    signal expr_207_wire_constant : std_logic_vector(7 downto 0);
    signal expr_214_wire_constant : std_logic_vector(7 downto 0);
    signal expr_221_wire_constant : std_logic_vector(7 downto 0);
    signal expr_228_wire_constant : std_logic_vector(7 downto 0);
    signal expr_235_wire_constant : std_logic_vector(7 downto 0);
    signal expr_242_wire_constant : std_logic_vector(7 downto 0);
    signal expr_249_wire_constant : std_logic_vector(7 downto 0);
    signal expr_256_wire_constant : std_logic_vector(7 downto 0);
    signal expr_263_wire_constant : std_logic_vector(7 downto 0);
    signal expr_270_wire_constant : std_logic_vector(7 downto 0);
    signal expr_277_wire_constant : std_logic_vector(7 downto 0);
    signal expr_284_wire_constant : std_logic_vector(7 downto 0);
    signal expr_291_wire_constant : std_logic_vector(7 downto 0);
    signal expr_298_wire_constant : std_logic_vector(7 downto 0);
    signal expr_305_wire_constant : std_logic_vector(7 downto 0);
    signal expr_312_wire_constant : std_logic_vector(7 downto 0);
    signal expr_319_wire_constant : std_logic_vector(7 downto 0);
    signal expr_326_wire_constant : std_logic_vector(7 downto 0);
    signal expr_333_wire_constant : std_logic_vector(7 downto 0);
    signal expr_340_wire_constant : std_logic_vector(7 downto 0);
    signal expr_347_wire_constant : std_logic_vector(7 downto 0);
    signal expr_354_wire_constant : std_logic_vector(7 downto 0);
    signal expr_361_wire_constant : std_logic_vector(7 downto 0);
    signal expr_368_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_176_word_address_0 <= "000000000";
    array_obj_ref_185_word_address_0 <= "000000001";
    array_obj_ref_192_word_address_0 <= "000000010";
    array_obj_ref_199_word_address_0 <= "000000011";
    array_obj_ref_206_word_address_0 <= "000000100";
    array_obj_ref_213_word_address_0 <= "000000101";
    array_obj_ref_220_word_address_0 <= "000000110";
    array_obj_ref_227_word_address_0 <= "001001000";
    array_obj_ref_234_word_address_0 <= "001001001";
    array_obj_ref_241_word_address_0 <= "001001010";
    array_obj_ref_248_word_address_0 <= "001001011";
    array_obj_ref_255_word_address_0 <= "001001100";
    array_obj_ref_262_word_address_0 <= "001001101";
    array_obj_ref_269_word_address_0 <= "001001110";
    array_obj_ref_276_word_address_0 <= "010010000";
    array_obj_ref_283_word_address_0 <= "010010001";
    array_obj_ref_290_word_address_0 <= "010010010";
    array_obj_ref_297_word_address_0 <= "010010011";
    array_obj_ref_304_word_address_0 <= "010010100";
    array_obj_ref_311_word_address_0 <= "010010101";
    array_obj_ref_318_word_address_0 <= "010010110";
    array_obj_ref_325_word_address_0 <= "011011000";
    array_obj_ref_332_word_address_0 <= "011011001";
    array_obj_ref_339_word_address_0 <= "011011010";
    array_obj_ref_346_word_address_0 <= "011011011";
    array_obj_ref_353_word_address_0 <= "011011100";
    array_obj_ref_360_word_address_0 <= "011011101";
    array_obj_ref_367_word_address_0 <= "011011110";
    expr_177_wire_constant <= "01110100";
    expr_186_wire_constant <= "01101111";
    expr_193_wire_constant <= "00110000";
    expr_200_wire_constant <= "01011111";
    expr_207_wire_constant <= "01101001";
    expr_214_wire_constant <= "01101110";
    expr_221_wire_constant <= "00110000";
    expr_228_wire_constant <= "01110100";
    expr_235_wire_constant <= "01101111";
    expr_242_wire_constant <= "00110001";
    expr_249_wire_constant <= "01011111";
    expr_256_wire_constant <= "01101001";
    expr_263_wire_constant <= "01101110";
    expr_270_wire_constant <= "00110000";
    expr_277_wire_constant <= "01110100";
    expr_284_wire_constant <= "01101111";
    expr_291_wire_constant <= "00110010";
    expr_298_wire_constant <= "01011111";
    expr_305_wire_constant <= "01101001";
    expr_312_wire_constant <= "01101110";
    expr_319_wire_constant <= "00110000";
    expr_326_wire_constant <= "01110100";
    expr_333_wire_constant <= "01101111";
    expr_340_wire_constant <= "00110011";
    expr_347_wire_constant <= "01011111";
    expr_354_wire_constant <= "01101001";
    expr_361_wire_constant <= "01101110";
    expr_368_wire_constant <= "00110000";
    array_obj_ref_176_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_176_gather_scatter_ack_0 <= array_obj_ref_176_gather_scatter_req_0;
      aggregated_sig <= expr_177_wire_constant;
      array_obj_ref_176_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_185_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_185_gather_scatter_ack_0 <= array_obj_ref_185_gather_scatter_req_0;
      aggregated_sig <= expr_186_wire_constant;
      array_obj_ref_185_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_192_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_192_gather_scatter_ack_0 <= array_obj_ref_192_gather_scatter_req_0;
      aggregated_sig <= expr_193_wire_constant;
      array_obj_ref_192_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_199_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_199_gather_scatter_ack_0 <= array_obj_ref_199_gather_scatter_req_0;
      aggregated_sig <= expr_200_wire_constant;
      array_obj_ref_199_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_206_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_206_gather_scatter_ack_0 <= array_obj_ref_206_gather_scatter_req_0;
      aggregated_sig <= expr_207_wire_constant;
      array_obj_ref_206_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_213_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_213_gather_scatter_ack_0 <= array_obj_ref_213_gather_scatter_req_0;
      aggregated_sig <= expr_214_wire_constant;
      array_obj_ref_213_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_220_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_220_gather_scatter_ack_0 <= array_obj_ref_220_gather_scatter_req_0;
      aggregated_sig <= expr_221_wire_constant;
      array_obj_ref_220_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_227_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_227_gather_scatter_ack_0 <= array_obj_ref_227_gather_scatter_req_0;
      aggregated_sig <= expr_228_wire_constant;
      array_obj_ref_227_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_234_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_234_gather_scatter_ack_0 <= array_obj_ref_234_gather_scatter_req_0;
      aggregated_sig <= expr_235_wire_constant;
      array_obj_ref_234_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_241_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_241_gather_scatter_ack_0 <= array_obj_ref_241_gather_scatter_req_0;
      aggregated_sig <= expr_242_wire_constant;
      array_obj_ref_241_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_248_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_248_gather_scatter_ack_0 <= array_obj_ref_248_gather_scatter_req_0;
      aggregated_sig <= expr_249_wire_constant;
      array_obj_ref_248_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_255_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_255_gather_scatter_ack_0 <= array_obj_ref_255_gather_scatter_req_0;
      aggregated_sig <= expr_256_wire_constant;
      array_obj_ref_255_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_262_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_262_gather_scatter_ack_0 <= array_obj_ref_262_gather_scatter_req_0;
      aggregated_sig <= expr_263_wire_constant;
      array_obj_ref_262_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_269_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_269_gather_scatter_ack_0 <= array_obj_ref_269_gather_scatter_req_0;
      aggregated_sig <= expr_270_wire_constant;
      array_obj_ref_269_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_276_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_276_gather_scatter_ack_0 <= array_obj_ref_276_gather_scatter_req_0;
      aggregated_sig <= expr_277_wire_constant;
      array_obj_ref_276_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_283_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_283_gather_scatter_ack_0 <= array_obj_ref_283_gather_scatter_req_0;
      aggregated_sig <= expr_284_wire_constant;
      array_obj_ref_283_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_290_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_290_gather_scatter_ack_0 <= array_obj_ref_290_gather_scatter_req_0;
      aggregated_sig <= expr_291_wire_constant;
      array_obj_ref_290_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_297_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_297_gather_scatter_ack_0 <= array_obj_ref_297_gather_scatter_req_0;
      aggregated_sig <= expr_298_wire_constant;
      array_obj_ref_297_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_304_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_304_gather_scatter_ack_0 <= array_obj_ref_304_gather_scatter_req_0;
      aggregated_sig <= expr_305_wire_constant;
      array_obj_ref_304_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_311_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_311_gather_scatter_ack_0 <= array_obj_ref_311_gather_scatter_req_0;
      aggregated_sig <= expr_312_wire_constant;
      array_obj_ref_311_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_318_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_318_gather_scatter_ack_0 <= array_obj_ref_318_gather_scatter_req_0;
      aggregated_sig <= expr_319_wire_constant;
      array_obj_ref_318_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_325_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_325_gather_scatter_ack_0 <= array_obj_ref_325_gather_scatter_req_0;
      aggregated_sig <= expr_326_wire_constant;
      array_obj_ref_325_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_332_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_332_gather_scatter_ack_0 <= array_obj_ref_332_gather_scatter_req_0;
      aggregated_sig <= expr_333_wire_constant;
      array_obj_ref_332_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_339_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_339_gather_scatter_ack_0 <= array_obj_ref_339_gather_scatter_req_0;
      aggregated_sig <= expr_340_wire_constant;
      array_obj_ref_339_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_346_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_346_gather_scatter_ack_0 <= array_obj_ref_346_gather_scatter_req_0;
      aggregated_sig <= expr_347_wire_constant;
      array_obj_ref_346_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_353_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_353_gather_scatter_ack_0 <= array_obj_ref_353_gather_scatter_req_0;
      aggregated_sig <= expr_354_wire_constant;
      array_obj_ref_353_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_360_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_360_gather_scatter_ack_0 <= array_obj_ref_360_gather_scatter_req_0;
      aggregated_sig <= expr_361_wire_constant;
      array_obj_ref_360_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    array_obj_ref_367_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      array_obj_ref_367_gather_scatter_ack_0 <= array_obj_ref_367_gather_scatter_req_0;
      aggregated_sig <= expr_368_wire_constant;
      array_obj_ref_367_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if array_obj_ref_176_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_176_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_176_word_address_0) &  " data array_obj_ref_176_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_176_data_0) severity note; --
        end if;
        if array_obj_ref_185_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_185_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_185_word_address_0) &  " data array_obj_ref_185_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_185_data_0) severity note; --
        end if;
        if array_obj_ref_192_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_192_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_192_word_address_0) &  " data array_obj_ref_192_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_192_data_0) severity note; --
        end if;
        if array_obj_ref_199_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_199_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_199_word_address_0) &  " data array_obj_ref_199_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_199_data_0) severity note; --
        end if;
        if array_obj_ref_206_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_206_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_206_word_address_0) &  " data array_obj_ref_206_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_206_data_0) severity note; --
        end if;
        if array_obj_ref_213_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_213_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_213_word_address_0) &  " data array_obj_ref_213_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_213_data_0) severity note; --
        end if;
        if array_obj_ref_220_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_220_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_220_word_address_0) &  " data array_obj_ref_220_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_220_data_0) severity note; --
        end if;
        if array_obj_ref_227_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_227_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_227_word_address_0) &  " data array_obj_ref_227_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_227_data_0) severity note; --
        end if;
        if array_obj_ref_234_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_234_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_234_word_address_0) &  " data array_obj_ref_234_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_234_data_0) severity note; --
        end if;
        if array_obj_ref_241_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_241_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_241_word_address_0) &  " data array_obj_ref_241_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_241_data_0) severity note; --
        end if;
        if array_obj_ref_248_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_248_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_248_word_address_0) &  " data array_obj_ref_248_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_248_data_0) severity note; --
        end if;
        if array_obj_ref_255_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_255_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_255_word_address_0) &  " data array_obj_ref_255_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_255_data_0) severity note; --
        end if;
        if array_obj_ref_262_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_262_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_262_word_address_0) &  " data array_obj_ref_262_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_262_data_0) severity note; --
        end if;
        if array_obj_ref_269_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_269_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_269_word_address_0) &  " data array_obj_ref_269_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_269_data_0) severity note; --
        end if;
        if array_obj_ref_276_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_276_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_276_word_address_0) &  " data array_obj_ref_276_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_276_data_0) severity note; --
        end if;
        if array_obj_ref_283_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_283_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_283_word_address_0) &  " data array_obj_ref_283_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_283_data_0) severity note; --
        end if;
        if array_obj_ref_290_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_290_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_290_word_address_0) &  " data array_obj_ref_290_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_290_data_0) severity note; --
        end if;
        if array_obj_ref_297_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_297_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_297_word_address_0) &  " data array_obj_ref_297_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_297_data_0) severity note; --
        end if;
        if array_obj_ref_304_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_304_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_304_word_address_0) &  " data array_obj_ref_304_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_304_data_0) severity note; --
        end if;
        if array_obj_ref_311_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_311_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_311_word_address_0) &  " data array_obj_ref_311_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_311_data_0) severity note; --
        end if;
        if array_obj_ref_318_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_318_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_318_word_address_0) &  " data array_obj_ref_318_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_318_data_0) severity note; --
        end if;
        if array_obj_ref_325_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_325_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_325_word_address_0) &  " data array_obj_ref_325_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_325_data_0) severity note; --
        end if;
        if array_obj_ref_332_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_332_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_332_word_address_0) &  " data array_obj_ref_332_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_332_data_0) severity note; --
        end if;
        if array_obj_ref_339_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_339_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_339_word_address_0) &  " data array_obj_ref_339_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_339_data_0) severity note; --
        end if;
        if array_obj_ref_346_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_346_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_346_word_address_0) &  " data array_obj_ref_346_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_346_data_0) severity note; --
        end if;
        if array_obj_ref_353_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_353_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_353_word_address_0) &  " data array_obj_ref_353_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_353_data_0) severity note; --
        end if;
        if array_obj_ref_360_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_360_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_360_word_address_0) &  " data array_obj_ref_360_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_360_data_0) severity note; --
        end if;
        if array_obj_ref_367_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_1 address array_obj_ref_367_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_367_word_address_0) &  " data array_obj_ref_367_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_367_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : array_obj_ref_176_store_0 array_obj_ref_185_store_0 array_obj_ref_192_store_0 array_obj_ref_199_store_0 array_obj_ref_206_store_0 array_obj_ref_213_store_0 array_obj_ref_220_store_0 array_obj_ref_227_store_0 array_obj_ref_234_store_0 array_obj_ref_241_store_0 array_obj_ref_248_store_0 array_obj_ref_255_store_0 array_obj_ref_262_store_0 array_obj_ref_269_store_0 array_obj_ref_276_store_0 array_obj_ref_283_store_0 array_obj_ref_290_store_0 array_obj_ref_297_store_0 array_obj_ref_304_store_0 array_obj_ref_311_store_0 array_obj_ref_318_store_0 array_obj_ref_325_store_0 array_obj_ref_332_store_0 array_obj_ref_339_store_0 array_obj_ref_346_store_0 array_obj_ref_353_store_0 array_obj_ref_360_store_0 array_obj_ref_367_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(251 downto 0);
      signal data_in: std_logic_vector(223 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 27 downto 0);
      -- 
    begin -- 
      reqL(27) <= array_obj_ref_176_store_0_req_0;
      reqL(26) <= array_obj_ref_185_store_0_req_0;
      reqL(25) <= array_obj_ref_192_store_0_req_0;
      reqL(24) <= array_obj_ref_199_store_0_req_0;
      reqL(23) <= array_obj_ref_206_store_0_req_0;
      reqL(22) <= array_obj_ref_213_store_0_req_0;
      reqL(21) <= array_obj_ref_220_store_0_req_0;
      reqL(20) <= array_obj_ref_227_store_0_req_0;
      reqL(19) <= array_obj_ref_234_store_0_req_0;
      reqL(18) <= array_obj_ref_241_store_0_req_0;
      reqL(17) <= array_obj_ref_248_store_0_req_0;
      reqL(16) <= array_obj_ref_255_store_0_req_0;
      reqL(15) <= array_obj_ref_262_store_0_req_0;
      reqL(14) <= array_obj_ref_269_store_0_req_0;
      reqL(13) <= array_obj_ref_276_store_0_req_0;
      reqL(12) <= array_obj_ref_283_store_0_req_0;
      reqL(11) <= array_obj_ref_290_store_0_req_0;
      reqL(10) <= array_obj_ref_297_store_0_req_0;
      reqL(9) <= array_obj_ref_304_store_0_req_0;
      reqL(8) <= array_obj_ref_311_store_0_req_0;
      reqL(7) <= array_obj_ref_318_store_0_req_0;
      reqL(6) <= array_obj_ref_325_store_0_req_0;
      reqL(5) <= array_obj_ref_332_store_0_req_0;
      reqL(4) <= array_obj_ref_339_store_0_req_0;
      reqL(3) <= array_obj_ref_346_store_0_req_0;
      reqL(2) <= array_obj_ref_353_store_0_req_0;
      reqL(1) <= array_obj_ref_360_store_0_req_0;
      reqL(0) <= array_obj_ref_367_store_0_req_0;
      array_obj_ref_176_store_0_ack_0 <= ackL(27);
      array_obj_ref_185_store_0_ack_0 <= ackL(26);
      array_obj_ref_192_store_0_ack_0 <= ackL(25);
      array_obj_ref_199_store_0_ack_0 <= ackL(24);
      array_obj_ref_206_store_0_ack_0 <= ackL(23);
      array_obj_ref_213_store_0_ack_0 <= ackL(22);
      array_obj_ref_220_store_0_ack_0 <= ackL(21);
      array_obj_ref_227_store_0_ack_0 <= ackL(20);
      array_obj_ref_234_store_0_ack_0 <= ackL(19);
      array_obj_ref_241_store_0_ack_0 <= ackL(18);
      array_obj_ref_248_store_0_ack_0 <= ackL(17);
      array_obj_ref_255_store_0_ack_0 <= ackL(16);
      array_obj_ref_262_store_0_ack_0 <= ackL(15);
      array_obj_ref_269_store_0_ack_0 <= ackL(14);
      array_obj_ref_276_store_0_ack_0 <= ackL(13);
      array_obj_ref_283_store_0_ack_0 <= ackL(12);
      array_obj_ref_290_store_0_ack_0 <= ackL(11);
      array_obj_ref_297_store_0_ack_0 <= ackL(10);
      array_obj_ref_304_store_0_ack_0 <= ackL(9);
      array_obj_ref_311_store_0_ack_0 <= ackL(8);
      array_obj_ref_318_store_0_ack_0 <= ackL(7);
      array_obj_ref_325_store_0_ack_0 <= ackL(6);
      array_obj_ref_332_store_0_ack_0 <= ackL(5);
      array_obj_ref_339_store_0_ack_0 <= ackL(4);
      array_obj_ref_346_store_0_ack_0 <= ackL(3);
      array_obj_ref_353_store_0_ack_0 <= ackL(2);
      array_obj_ref_360_store_0_ack_0 <= ackL(1);
      array_obj_ref_367_store_0_ack_0 <= ackL(0);
      reqR(27) <= array_obj_ref_176_store_0_req_1;
      reqR(26) <= array_obj_ref_185_store_0_req_1;
      reqR(25) <= array_obj_ref_192_store_0_req_1;
      reqR(24) <= array_obj_ref_199_store_0_req_1;
      reqR(23) <= array_obj_ref_206_store_0_req_1;
      reqR(22) <= array_obj_ref_213_store_0_req_1;
      reqR(21) <= array_obj_ref_220_store_0_req_1;
      reqR(20) <= array_obj_ref_227_store_0_req_1;
      reqR(19) <= array_obj_ref_234_store_0_req_1;
      reqR(18) <= array_obj_ref_241_store_0_req_1;
      reqR(17) <= array_obj_ref_248_store_0_req_1;
      reqR(16) <= array_obj_ref_255_store_0_req_1;
      reqR(15) <= array_obj_ref_262_store_0_req_1;
      reqR(14) <= array_obj_ref_269_store_0_req_1;
      reqR(13) <= array_obj_ref_276_store_0_req_1;
      reqR(12) <= array_obj_ref_283_store_0_req_1;
      reqR(11) <= array_obj_ref_290_store_0_req_1;
      reqR(10) <= array_obj_ref_297_store_0_req_1;
      reqR(9) <= array_obj_ref_304_store_0_req_1;
      reqR(8) <= array_obj_ref_311_store_0_req_1;
      reqR(7) <= array_obj_ref_318_store_0_req_1;
      reqR(6) <= array_obj_ref_325_store_0_req_1;
      reqR(5) <= array_obj_ref_332_store_0_req_1;
      reqR(4) <= array_obj_ref_339_store_0_req_1;
      reqR(3) <= array_obj_ref_346_store_0_req_1;
      reqR(2) <= array_obj_ref_353_store_0_req_1;
      reqR(1) <= array_obj_ref_360_store_0_req_1;
      reqR(0) <= array_obj_ref_367_store_0_req_1;
      array_obj_ref_176_store_0_ack_1 <= ackR(27);
      array_obj_ref_185_store_0_ack_1 <= ackR(26);
      array_obj_ref_192_store_0_ack_1 <= ackR(25);
      array_obj_ref_199_store_0_ack_1 <= ackR(24);
      array_obj_ref_206_store_0_ack_1 <= ackR(23);
      array_obj_ref_213_store_0_ack_1 <= ackR(22);
      array_obj_ref_220_store_0_ack_1 <= ackR(21);
      array_obj_ref_227_store_0_ack_1 <= ackR(20);
      array_obj_ref_234_store_0_ack_1 <= ackR(19);
      array_obj_ref_241_store_0_ack_1 <= ackR(18);
      array_obj_ref_248_store_0_ack_1 <= ackR(17);
      array_obj_ref_255_store_0_ack_1 <= ackR(16);
      array_obj_ref_262_store_0_ack_1 <= ackR(15);
      array_obj_ref_269_store_0_ack_1 <= ackR(14);
      array_obj_ref_276_store_0_ack_1 <= ackR(13);
      array_obj_ref_283_store_0_ack_1 <= ackR(12);
      array_obj_ref_290_store_0_ack_1 <= ackR(11);
      array_obj_ref_297_store_0_ack_1 <= ackR(10);
      array_obj_ref_304_store_0_ack_1 <= ackR(9);
      array_obj_ref_311_store_0_ack_1 <= ackR(8);
      array_obj_ref_318_store_0_ack_1 <= ackR(7);
      array_obj_ref_325_store_0_ack_1 <= ackR(6);
      array_obj_ref_332_store_0_ack_1 <= ackR(5);
      array_obj_ref_339_store_0_ack_1 <= ackR(4);
      array_obj_ref_346_store_0_ack_1 <= ackR(3);
      array_obj_ref_353_store_0_ack_1 <= ackR(2);
      array_obj_ref_360_store_0_ack_1 <= ackR(1);
      array_obj_ref_367_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_176_word_address_0 & array_obj_ref_185_word_address_0 & array_obj_ref_192_word_address_0 & array_obj_ref_199_word_address_0 & array_obj_ref_206_word_address_0 & array_obj_ref_213_word_address_0 & array_obj_ref_220_word_address_0 & array_obj_ref_227_word_address_0 & array_obj_ref_234_word_address_0 & array_obj_ref_241_word_address_0 & array_obj_ref_248_word_address_0 & array_obj_ref_255_word_address_0 & array_obj_ref_262_word_address_0 & array_obj_ref_269_word_address_0 & array_obj_ref_276_word_address_0 & array_obj_ref_283_word_address_0 & array_obj_ref_290_word_address_0 & array_obj_ref_297_word_address_0 & array_obj_ref_304_word_address_0 & array_obj_ref_311_word_address_0 & array_obj_ref_318_word_address_0 & array_obj_ref_325_word_address_0 & array_obj_ref_332_word_address_0 & array_obj_ref_339_word_address_0 & array_obj_ref_346_word_address_0 & array_obj_ref_353_word_address_0 & array_obj_ref_360_word_address_0 & array_obj_ref_367_word_address_0;
      data_in <= array_obj_ref_176_data_0 & array_obj_ref_185_data_0 & array_obj_ref_192_data_0 & array_obj_ref_199_data_0 & array_obj_ref_206_data_0 & array_obj_ref_213_data_0 & array_obj_ref_220_data_0 & array_obj_ref_227_data_0 & array_obj_ref_234_data_0 & array_obj_ref_241_data_0 & array_obj_ref_248_data_0 & array_obj_ref_255_data_0 & array_obj_ref_262_data_0 & array_obj_ref_269_data_0 & array_obj_ref_276_data_0 & array_obj_ref_283_data_0 & array_obj_ref_290_data_0 & array_obj_ref_297_data_0 & array_obj_ref_304_data_0 & array_obj_ref_311_data_0 & array_obj_ref_318_data_0 & array_obj_ref_325_data_0 & array_obj_ref_332_data_0 & array_obj_ref_339_data_0 & array_obj_ref_346_data_0 & array_obj_ref_353_data_0 & array_obj_ref_360_data_0 & array_obj_ref_367_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 9,
        data_width => 8,
        num_reqs => 28,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(8 downto 0),
          mdata => memory_space_1_sr_data(7 downto 0),
          mtag => memory_space_1_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 28,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity GV_16_initializer_in_click_bc is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(4 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity GV_16_initializer_in_click_bc;
architecture Default of GV_16_initializer_in_click_bc is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal GV_16_initializer_in_click_bc_CP_591_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_376_gather_scatter_req_0 : boolean;
  signal array_obj_ref_376_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_376_store_0_req_0 : boolean;
  signal array_obj_ref_376_store_0_ack_0 : boolean;
  signal array_obj_ref_376_store_0_req_1 : boolean;
  signal array_obj_ref_376_store_0_ack_1 : boolean;
  signal array_obj_ref_388_gather_scatter_req_0 : boolean;
  signal array_obj_ref_388_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_388_store_0_req_0 : boolean;
  signal array_obj_ref_388_store_0_ack_0 : boolean;
  signal array_obj_ref_388_store_0_req_1 : boolean;
  signal array_obj_ref_388_store_0_ack_1 : boolean;
  signal array_obj_ref_395_gather_scatter_req_0 : boolean;
  signal array_obj_ref_395_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_395_store_0_req_0 : boolean;
  signal array_obj_ref_395_store_0_ack_0 : boolean;
  signal array_obj_ref_395_store_0_req_1 : boolean;
  signal array_obj_ref_395_store_0_ack_1 : boolean;
  signal array_obj_ref_402_gather_scatter_req_0 : boolean;
  signal array_obj_ref_402_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_402_store_0_req_0 : boolean;
  signal array_obj_ref_402_store_0_ack_0 : boolean;
  signal array_obj_ref_402_store_0_req_1 : boolean;
  signal array_obj_ref_402_store_0_ack_1 : boolean;
  signal array_obj_ref_410_gather_scatter_req_0 : boolean;
  signal array_obj_ref_410_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_410_store_0_req_0 : boolean;
  signal array_obj_ref_410_store_0_ack_0 : boolean;
  signal array_obj_ref_410_store_0_req_1 : boolean;
  signal array_obj_ref_410_store_0_ack_1 : boolean;
  signal array_obj_ref_417_gather_scatter_req_0 : boolean;
  signal array_obj_ref_417_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_417_store_0_req_0 : boolean;
  signal array_obj_ref_417_store_0_ack_0 : boolean;
  signal array_obj_ref_417_store_0_req_1 : boolean;
  signal array_obj_ref_417_store_0_ack_1 : boolean;
  signal array_obj_ref_423_gather_scatter_req_0 : boolean;
  signal array_obj_ref_423_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_423_store_0_req_0 : boolean;
  signal array_obj_ref_423_store_0_ack_0 : boolean;
  signal array_obj_ref_423_store_0_req_1 : boolean;
  signal array_obj_ref_423_store_0_ack_1 : boolean;
  signal array_obj_ref_430_gather_scatter_req_0 : boolean;
  signal array_obj_ref_430_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_430_store_0_req_0 : boolean;
  signal array_obj_ref_430_store_0_ack_0 : boolean;
  signal array_obj_ref_430_store_0_req_1 : boolean;
  signal array_obj_ref_430_store_0_ack_1 : boolean;
  signal array_obj_ref_438_gather_scatter_req_0 : boolean;
  signal array_obj_ref_438_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_0 : boolean;
  signal array_obj_ref_438_store_0_ack_0 : boolean;
  signal array_obj_ref_438_store_0_req_1 : boolean;
  signal array_obj_ref_438_store_0_ack_1 : boolean;
  signal array_obj_ref_445_gather_scatter_req_0 : boolean;
  signal array_obj_ref_445_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_445_store_0_req_0 : boolean;
  signal array_obj_ref_445_store_0_ack_0 : boolean;
  signal array_obj_ref_445_store_0_req_1 : boolean;
  signal array_obj_ref_445_store_0_ack_1 : boolean;
  signal array_obj_ref_451_gather_scatter_req_0 : boolean;
  signal array_obj_ref_451_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_451_store_0_req_0 : boolean;
  signal array_obj_ref_451_store_0_ack_0 : boolean;
  signal array_obj_ref_451_store_0_req_1 : boolean;
  signal array_obj_ref_451_store_0_ack_1 : boolean;
  signal array_obj_ref_458_gather_scatter_req_0 : boolean;
  signal array_obj_ref_458_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_0 : boolean;
  signal array_obj_ref_458_store_0_ack_0 : boolean;
  signal array_obj_ref_458_store_0_req_1 : boolean;
  signal array_obj_ref_458_store_0_ack_1 : boolean;
  signal array_obj_ref_466_gather_scatter_req_0 : boolean;
  signal array_obj_ref_466_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_0 : boolean;
  signal array_obj_ref_466_store_0_ack_0 : boolean;
  signal array_obj_ref_466_store_0_req_1 : boolean;
  signal array_obj_ref_466_store_0_ack_1 : boolean;
  signal array_obj_ref_473_gather_scatter_req_0 : boolean;
  signal array_obj_ref_473_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_473_store_0_req_0 : boolean;
  signal array_obj_ref_473_store_0_ack_0 : boolean;
  signal array_obj_ref_473_store_0_req_1 : boolean;
  signal array_obj_ref_473_store_0_ack_1 : boolean;
  signal array_obj_ref_479_gather_scatter_req_0 : boolean;
  signal array_obj_ref_479_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_479_store_0_req_0 : boolean;
  signal array_obj_ref_479_store_0_ack_0 : boolean;
  signal array_obj_ref_479_store_0_req_1 : boolean;
  signal array_obj_ref_479_store_0_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  GV_16_initializer_in_click_bc_CP_591: Block -- control-path 
    signal cp_elements: BooleanArray(45 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(45);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(45), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    split_req_603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => array_obj_ref_376_gather_scatter_req_0); -- 
    split_ack_604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_gather_scatter_ack_0, ack => cp_elements(1)); -- 
    rr_611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => array_obj_ref_376_store_0_req_0); -- 
    ra_612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_store_0_ack_0, ack => cp_elements(2)); -- 
    cr_613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => array_obj_ref_376_store_0_req_1); -- 
    ca_614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_376_store_0_ack_1, ack => cp_elements(3)); -- 
    split_req_624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => array_obj_ref_388_gather_scatter_req_0); -- 
    split_ack_625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_gather_scatter_ack_0, ack => cp_elements(4)); -- 
    rr_632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => array_obj_ref_388_store_0_req_0); -- 
    ra_633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_store_0_ack_0, ack => cp_elements(5)); -- 
    cr_634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => array_obj_ref_388_store_0_req_1); -- 
    ca_635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_388_store_0_ack_1, ack => cp_elements(6)); -- 
    split_req_645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => array_obj_ref_395_gather_scatter_req_0); -- 
    split_ack_646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_gather_scatter_ack_0, ack => cp_elements(7)); -- 
    rr_653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => array_obj_ref_395_store_0_req_0); -- 
    ra_654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_store_0_ack_0, ack => cp_elements(8)); -- 
    cr_655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => array_obj_ref_395_store_0_req_1); -- 
    ca_656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_395_store_0_ack_1, ack => cp_elements(9)); -- 
    split_req_666_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => array_obj_ref_402_gather_scatter_req_0); -- 
    split_ack_667_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => array_obj_ref_402_store_0_req_0); -- 
    ra_675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => array_obj_ref_402_store_0_req_1); -- 
    ca_677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_402_store_0_ack_1, ack => cp_elements(12)); -- 
    split_req_687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => array_obj_ref_410_gather_scatter_req_0); -- 
    split_ack_688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => array_obj_ref_410_store_0_req_0); -- 
    ra_696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_store_0_ack_0, ack => cp_elements(14)); -- 
    cr_697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => array_obj_ref_410_store_0_req_1); -- 
    ca_698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_410_store_0_ack_1, ack => cp_elements(15)); -- 
    split_req_708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => array_obj_ref_417_gather_scatter_req_0); -- 
    split_ack_709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_417_store_0_req_0); -- 
    ra_717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_store_0_ack_0, ack => cp_elements(17)); -- 
    cr_718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_417_store_0_req_1); -- 
    ca_719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_417_store_0_ack_1, ack => cp_elements(18)); -- 
    split_req_729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_423_gather_scatter_req_0); -- 
    split_ack_730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_gather_scatter_ack_0, ack => cp_elements(19)); -- 
    rr_737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => array_obj_ref_423_store_0_req_0); -- 
    ra_738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_0, ack => cp_elements(20)); -- 
    cr_739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => array_obj_ref_423_store_0_req_1); -- 
    ca_740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_423_store_0_ack_1, ack => cp_elements(21)); -- 
    split_req_750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_430_gather_scatter_req_0); -- 
    split_ack_751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_gather_scatter_ack_0, ack => cp_elements(22)); -- 
    rr_758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_430_store_0_req_0); -- 
    ra_759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_0, ack => cp_elements(23)); -- 
    cr_760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_430_store_0_req_1); -- 
    ca_761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_store_0_ack_1, ack => cp_elements(24)); -- 
    split_req_771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => array_obj_ref_438_gather_scatter_req_0); -- 
    split_ack_772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    rr_779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => array_obj_ref_438_store_0_req_0); -- 
    ra_780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_0, ack => cp_elements(26)); -- 
    cr_781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => array_obj_ref_438_store_0_req_1); -- 
    ca_782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_438_store_0_ack_1, ack => cp_elements(27)); -- 
    split_req_792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_445_gather_scatter_req_0); -- 
    split_ack_793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    rr_800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => array_obj_ref_445_store_0_req_0); -- 
    ra_801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_store_0_ack_0, ack => cp_elements(29)); -- 
    cr_802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_445_store_0_req_1); -- 
    ca_803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_445_store_0_ack_1, ack => cp_elements(30)); -- 
    split_req_813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_451_gather_scatter_req_0); -- 
    split_ack_814_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_gather_scatter_ack_0, ack => cp_elements(31)); -- 
    rr_821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_451_store_0_req_0); -- 
    ra_822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_store_0_ack_0, ack => cp_elements(32)); -- 
    cr_823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_451_store_0_req_1); -- 
    ca_824_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_store_0_ack_1, ack => cp_elements(33)); -- 
    split_req_834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_458_gather_scatter_req_0); -- 
    split_ack_835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_gather_scatter_ack_0, ack => cp_elements(34)); -- 
    rr_842_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_458_store_0_req_0); -- 
    ra_843_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_store_0_ack_0, ack => cp_elements(35)); -- 
    cr_844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_458_store_0_req_1); -- 
    ca_845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_458_store_0_ack_1, ack => cp_elements(36)); -- 
    split_req_855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_466_gather_scatter_req_0); -- 
    split_ack_856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_gather_scatter_ack_0, ack => cp_elements(37)); -- 
    rr_863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_466_store_0_req_0); -- 
    ra_864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_store_0_ack_0, ack => cp_elements(38)); -- 
    cr_865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_466_store_0_req_1); -- 
    ca_866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_466_store_0_ack_1, ack => cp_elements(39)); -- 
    split_req_876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => array_obj_ref_473_gather_scatter_req_0); -- 
    split_ack_877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_gather_scatter_ack_0, ack => cp_elements(40)); -- 
    rr_884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => array_obj_ref_473_store_0_req_0); -- 
    ra_885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_store_0_ack_0, ack => cp_elements(41)); -- 
    cr_886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => array_obj_ref_473_store_0_req_1); -- 
    ca_887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_473_store_0_ack_1, ack => cp_elements(42)); -- 
    split_req_897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => array_obj_ref_479_gather_scatter_req_0); -- 
    split_ack_898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_gather_scatter_ack_0, ack => cp_elements(43)); -- 
    rr_905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => array_obj_ref_479_store_0_req_0); -- 
    ra_906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_store_0_ack_0, ack => cp_elements(44)); -- 
    cr_907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => array_obj_ref_479_store_0_req_1); -- 
    ca_908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_479_store_0_ack_1, ack => cp_elements(45)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_376_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_376_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_388_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_388_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_395_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_395_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_402_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_402_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_410_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_410_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_417_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_417_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_423_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_423_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_430_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_430_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_438_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_438_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_445_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_445_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_451_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_451_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_458_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_458_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_466_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_466_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_473_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_473_word_address_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_479_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_479_word_address_0 : std_logic_vector(4 downto 0);
    signal expr_377_wire_constant : std_logic_vector(31 downto 0);
    signal expr_389_wire_constant : std_logic_vector(31 downto 0);
    signal expr_396_wire_constant : std_logic_vector(31 downto 0);
    signal expr_403_wire_constant : std_logic_vector(31 downto 0);
    signal expr_411_wire_constant : std_logic_vector(31 downto 0);
    signal expr_418_wire_constant : std_logic_vector(31 downto 0);
    signal expr_424_wire_constant : std_logic_vector(31 downto 0);
    signal expr_431_wire_constant : std_logic_vector(31 downto 0);
    signal expr_439_wire_constant : std_logic_vector(31 downto 0);
    signal expr_446_wire_constant : std_logic_vector(31 downto 0);
    signal expr_452_wire_constant : std_logic_vector(31 downto 0);
    signal expr_459_wire_constant : std_logic_vector(31 downto 0);
    signal expr_467_wire_constant : std_logic_vector(31 downto 0);
    signal expr_474_wire_constant : std_logic_vector(31 downto 0);
    signal expr_480_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_376_word_address_0 <= "00000";
    array_obj_ref_388_word_address_0 <= "00001";
    array_obj_ref_395_word_address_0 <= "00100";
    array_obj_ref_402_word_address_0 <= "00101";
    array_obj_ref_410_word_address_0 <= "00110";
    array_obj_ref_417_word_address_0 <= "01000";
    array_obj_ref_423_word_address_0 <= "01001";
    array_obj_ref_430_word_address_0 <= "01010";
    array_obj_ref_438_word_address_0 <= "01011";
    array_obj_ref_445_word_address_0 <= "01101";
    array_obj_ref_451_word_address_0 <= "01110";
    array_obj_ref_458_word_address_0 <= "01111";
    array_obj_ref_466_word_address_0 <= "10000";
    array_obj_ref_473_word_address_0 <= "10010";
    array_obj_ref_479_word_address_0 <= "10011";
    expr_377_wire_constant <= "00000000000000000001000010101100";
    expr_389_wire_constant <= "00000000111111111111111111111111";
    expr_396_wire_constant <= "01111111111111111111111111111111";
    expr_403_wire_constant <= "00000000000000010001000010101100";
    expr_411_wire_constant <= "00000000111111111111111111111111";
    expr_418_wire_constant <= "00000000000000000000000000000001";
    expr_424_wire_constant <= "01111111111111111111111111111111";
    expr_431_wire_constant <= "00000000000000100001000010101100";
    expr_439_wire_constant <= "00000000111111111111111111111111";
    expr_446_wire_constant <= "00000000000000000000000000000010";
    expr_452_wire_constant <= "01111111111111111111111111111111";
    expr_459_wire_constant <= "00000000000000110001000010101100";
    expr_467_wire_constant <= "00000000111111111111111111111111";
    expr_474_wire_constant <= "00000000000000000000000000000011";
    expr_480_wire_constant <= "01111111111111111111111111111111";
    array_obj_ref_376_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_376_gather_scatter_ack_0 <= array_obj_ref_376_gather_scatter_req_0;
      aggregated_sig <= expr_377_wire_constant;
      array_obj_ref_376_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_388_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_388_gather_scatter_ack_0 <= array_obj_ref_388_gather_scatter_req_0;
      aggregated_sig <= expr_389_wire_constant;
      array_obj_ref_388_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_395_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_395_gather_scatter_ack_0 <= array_obj_ref_395_gather_scatter_req_0;
      aggregated_sig <= expr_396_wire_constant;
      array_obj_ref_395_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_402_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_402_gather_scatter_ack_0 <= array_obj_ref_402_gather_scatter_req_0;
      aggregated_sig <= expr_403_wire_constant;
      array_obj_ref_402_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_410_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_410_gather_scatter_ack_0 <= array_obj_ref_410_gather_scatter_req_0;
      aggregated_sig <= expr_411_wire_constant;
      array_obj_ref_410_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_417_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_417_gather_scatter_ack_0 <= array_obj_ref_417_gather_scatter_req_0;
      aggregated_sig <= expr_418_wire_constant;
      array_obj_ref_417_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_423_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_423_gather_scatter_ack_0 <= array_obj_ref_423_gather_scatter_req_0;
      aggregated_sig <= expr_424_wire_constant;
      array_obj_ref_423_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_430_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_430_gather_scatter_ack_0 <= array_obj_ref_430_gather_scatter_req_0;
      aggregated_sig <= expr_431_wire_constant;
      array_obj_ref_430_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_438_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_438_gather_scatter_ack_0 <= array_obj_ref_438_gather_scatter_req_0;
      aggregated_sig <= expr_439_wire_constant;
      array_obj_ref_438_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_445_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_445_gather_scatter_ack_0 <= array_obj_ref_445_gather_scatter_req_0;
      aggregated_sig <= expr_446_wire_constant;
      array_obj_ref_445_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_451_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_451_gather_scatter_ack_0 <= array_obj_ref_451_gather_scatter_req_0;
      aggregated_sig <= expr_452_wire_constant;
      array_obj_ref_451_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_458_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_458_gather_scatter_ack_0 <= array_obj_ref_458_gather_scatter_req_0;
      aggregated_sig <= expr_459_wire_constant;
      array_obj_ref_458_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_466_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_466_gather_scatter_ack_0 <= array_obj_ref_466_gather_scatter_req_0;
      aggregated_sig <= expr_467_wire_constant;
      array_obj_ref_466_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_473_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_473_gather_scatter_ack_0 <= array_obj_ref_473_gather_scatter_req_0;
      aggregated_sig <= expr_474_wire_constant;
      array_obj_ref_473_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    array_obj_ref_479_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      array_obj_ref_479_gather_scatter_ack_0 <= array_obj_ref_479_gather_scatter_req_0;
      aggregated_sig <= expr_480_wire_constant;
      array_obj_ref_479_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if array_obj_ref_410_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_410_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_410_word_address_0) &  " data array_obj_ref_410_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_410_data_0) severity note; --
        end if;
        if array_obj_ref_417_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_417_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_417_word_address_0) &  " data array_obj_ref_417_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_417_data_0) severity note; --
        end if;
        if array_obj_ref_466_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_466_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_466_word_address_0) &  " data array_obj_ref_466_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_466_data_0) severity note; --
        end if;
        if array_obj_ref_458_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_458_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_458_word_address_0) &  " data array_obj_ref_458_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_458_data_0) severity note; --
        end if;
        if array_obj_ref_402_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_402_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_402_word_address_0) &  " data array_obj_ref_402_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_402_data_0) severity note; --
        end if;
        if array_obj_ref_451_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_451_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_451_word_address_0) &  " data array_obj_ref_451_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_451_data_0) severity note; --
        end if;
        if array_obj_ref_445_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_445_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_445_word_address_0) &  " data array_obj_ref_445_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_445_data_0) severity note; --
        end if;
        if array_obj_ref_395_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_395_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_395_word_address_0) &  " data array_obj_ref_395_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_395_data_0) severity note; --
        end if;
        if array_obj_ref_479_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_479_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_479_word_address_0) &  " data array_obj_ref_479_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_479_data_0) severity note; --
        end if;
        if array_obj_ref_438_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_438_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_438_word_address_0) &  " data array_obj_ref_438_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_438_data_0) severity note; --
        end if;
        if array_obj_ref_388_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_388_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_388_word_address_0) &  " data array_obj_ref_388_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_388_data_0) severity note; --
        end if;
        if array_obj_ref_430_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_430_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_430_word_address_0) &  " data array_obj_ref_430_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_430_data_0) severity note; --
        end if;
        if array_obj_ref_376_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_376_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_376_word_address_0) &  " data array_obj_ref_376_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_376_data_0) severity note; --
        end if;
        if array_obj_ref_423_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_423_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_423_word_address_0) &  " data array_obj_ref_423_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_423_data_0) severity note; --
        end if;
        if array_obj_ref_473_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_2 address array_obj_ref_473_word_address_0 ="  &  convert_slv_to_hex_string(array_obj_ref_473_word_address_0) &  " data array_obj_ref_473_data_0 ="  &  convert_slv_to_hex_string(array_obj_ref_473_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : array_obj_ref_410_store_0 array_obj_ref_417_store_0 array_obj_ref_466_store_0 array_obj_ref_458_store_0 array_obj_ref_402_store_0 array_obj_ref_451_store_0 array_obj_ref_445_store_0 array_obj_ref_395_store_0 array_obj_ref_479_store_0 array_obj_ref_438_store_0 array_obj_ref_388_store_0 array_obj_ref_430_store_0 array_obj_ref_376_store_0 array_obj_ref_423_store_0 array_obj_ref_473_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(74 downto 0);
      signal data_in: std_logic_vector(479 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= array_obj_ref_410_store_0_req_0;
      reqL(13) <= array_obj_ref_417_store_0_req_0;
      reqL(12) <= array_obj_ref_466_store_0_req_0;
      reqL(11) <= array_obj_ref_458_store_0_req_0;
      reqL(10) <= array_obj_ref_402_store_0_req_0;
      reqL(9) <= array_obj_ref_451_store_0_req_0;
      reqL(8) <= array_obj_ref_445_store_0_req_0;
      reqL(7) <= array_obj_ref_395_store_0_req_0;
      reqL(6) <= array_obj_ref_479_store_0_req_0;
      reqL(5) <= array_obj_ref_438_store_0_req_0;
      reqL(4) <= array_obj_ref_388_store_0_req_0;
      reqL(3) <= array_obj_ref_430_store_0_req_0;
      reqL(2) <= array_obj_ref_376_store_0_req_0;
      reqL(1) <= array_obj_ref_423_store_0_req_0;
      reqL(0) <= array_obj_ref_473_store_0_req_0;
      array_obj_ref_410_store_0_ack_0 <= ackL(14);
      array_obj_ref_417_store_0_ack_0 <= ackL(13);
      array_obj_ref_466_store_0_ack_0 <= ackL(12);
      array_obj_ref_458_store_0_ack_0 <= ackL(11);
      array_obj_ref_402_store_0_ack_0 <= ackL(10);
      array_obj_ref_451_store_0_ack_0 <= ackL(9);
      array_obj_ref_445_store_0_ack_0 <= ackL(8);
      array_obj_ref_395_store_0_ack_0 <= ackL(7);
      array_obj_ref_479_store_0_ack_0 <= ackL(6);
      array_obj_ref_438_store_0_ack_0 <= ackL(5);
      array_obj_ref_388_store_0_ack_0 <= ackL(4);
      array_obj_ref_430_store_0_ack_0 <= ackL(3);
      array_obj_ref_376_store_0_ack_0 <= ackL(2);
      array_obj_ref_423_store_0_ack_0 <= ackL(1);
      array_obj_ref_473_store_0_ack_0 <= ackL(0);
      reqR(14) <= array_obj_ref_410_store_0_req_1;
      reqR(13) <= array_obj_ref_417_store_0_req_1;
      reqR(12) <= array_obj_ref_466_store_0_req_1;
      reqR(11) <= array_obj_ref_458_store_0_req_1;
      reqR(10) <= array_obj_ref_402_store_0_req_1;
      reqR(9) <= array_obj_ref_451_store_0_req_1;
      reqR(8) <= array_obj_ref_445_store_0_req_1;
      reqR(7) <= array_obj_ref_395_store_0_req_1;
      reqR(6) <= array_obj_ref_479_store_0_req_1;
      reqR(5) <= array_obj_ref_438_store_0_req_1;
      reqR(4) <= array_obj_ref_388_store_0_req_1;
      reqR(3) <= array_obj_ref_430_store_0_req_1;
      reqR(2) <= array_obj_ref_376_store_0_req_1;
      reqR(1) <= array_obj_ref_423_store_0_req_1;
      reqR(0) <= array_obj_ref_473_store_0_req_1;
      array_obj_ref_410_store_0_ack_1 <= ackR(14);
      array_obj_ref_417_store_0_ack_1 <= ackR(13);
      array_obj_ref_466_store_0_ack_1 <= ackR(12);
      array_obj_ref_458_store_0_ack_1 <= ackR(11);
      array_obj_ref_402_store_0_ack_1 <= ackR(10);
      array_obj_ref_451_store_0_ack_1 <= ackR(9);
      array_obj_ref_445_store_0_ack_1 <= ackR(8);
      array_obj_ref_395_store_0_ack_1 <= ackR(7);
      array_obj_ref_479_store_0_ack_1 <= ackR(6);
      array_obj_ref_438_store_0_ack_1 <= ackR(5);
      array_obj_ref_388_store_0_ack_1 <= ackR(4);
      array_obj_ref_430_store_0_ack_1 <= ackR(3);
      array_obj_ref_376_store_0_ack_1 <= ackR(2);
      array_obj_ref_423_store_0_ack_1 <= ackR(1);
      array_obj_ref_473_store_0_ack_1 <= ackR(0);
      addr_in <= array_obj_ref_410_word_address_0 & array_obj_ref_417_word_address_0 & array_obj_ref_466_word_address_0 & array_obj_ref_458_word_address_0 & array_obj_ref_402_word_address_0 & array_obj_ref_451_word_address_0 & array_obj_ref_445_word_address_0 & array_obj_ref_395_word_address_0 & array_obj_ref_479_word_address_0 & array_obj_ref_438_word_address_0 & array_obj_ref_388_word_address_0 & array_obj_ref_430_word_address_0 & array_obj_ref_376_word_address_0 & array_obj_ref_423_word_address_0 & array_obj_ref_473_word_address_0;
      data_in <= array_obj_ref_410_data_0 & array_obj_ref_417_data_0 & array_obj_ref_466_data_0 & array_obj_ref_458_data_0 & array_obj_ref_402_data_0 & array_obj_ref_451_data_0 & array_obj_ref_445_data_0 & array_obj_ref_395_data_0 & array_obj_ref_479_data_0 & array_obj_ref_438_data_0 & array_obj_ref_388_data_0 & array_obj_ref_430_data_0 & array_obj_ref_376_data_0 & array_obj_ref_423_data_0 & array_obj_ref_473_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 5,
        data_width => 32,
        num_reqs => 15,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(4 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_bswap_i16 is -- 
  generic (tag_length : integer); 
  port ( -- 
    i : in  std_logic_vector(15 downto 0);
    ret_val_x_x : out  std_logic_vector(15 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_bswap_i16;
architecture Default of ahir_glue_bswap_i16 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ret_val_x_x_buffer :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_CP_969_start: Boolean;
  -- links between control-path and data-path
  signal binary_523_inst_ack_1 : boolean;
  signal binary_523_inst_ack_0 : boolean;
  signal binary_523_inst_req_1 : boolean;
  signal binary_528_inst_req_0 : boolean;
  signal binary_528_inst_ack_0 : boolean;
  signal binary_528_inst_req_1 : boolean;
  signal binary_528_inst_ack_1 : boolean;
  signal binary_523_inst_req_0 : boolean;
  signal binary_517_inst_ack_1 : boolean;
  signal binary_517_inst_req_1 : boolean;
  signal binary_517_inst_req_0 : boolean;
  signal binary_517_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  ret_val_x_x <= ret_val_x_x_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 3, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_bswap_i16_CP_969: Block -- control-path 
    signal cp_elements: BooleanArray(15 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(15);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(15), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cpelement_group_2 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(4));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => binary_517_inst_req_0); -- 
    cp_elements(3) <= cp_elements(1);
    cp_elements(4) <= cp_elements(1);
    ra_993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_517_inst_ack_0, ack => cp_elements(5)); -- 
    cr_994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => binary_517_inst_req_1); -- 
    ca_995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_517_inst_ack_1, ack => cp_elements(6)); -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => binary_523_inst_req_0); -- 
    cp_elements(8) <= cp_elements(1);
    cp_elements(9) <= cp_elements(1);
    ra_1005_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_523_inst_ack_0, ack => cp_elements(10)); -- 
    cr_1006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_523_inst_req_1); -- 
    ca_1007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_523_inst_ack_1, ack => cp_elements(11)); -- 
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(13) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => binary_528_inst_req_0); -- 
    cp_elements(13) <= cp_elements(1);
    ra_1018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_528_inst_ack_0, ack => cp_elements(14)); -- 
    cr_1019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => binary_528_inst_req_1); -- 
    ca_1020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_528_inst_ack_1, ack => cp_elements(15)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal tmp1_524 : std_logic_vector(15 downto 0);
    signal tmp_518 : std_logic_vector(15 downto 0);
    signal type_cast_516_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_522_wire_constant : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    type_cast_516_wire_constant <= "0000000000001000";
    type_cast_522_wire_constant <= "0000000000001000";
    -- shared split operator group (0) : binary_517_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i;
      tmp_518 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_517_inst_req_0,
          ackL => binary_517_inst_ack_0,
          reqR => binary_517_inst_req_1,
          ackR => binary_517_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_523_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= i;
      tmp1_524 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_523_inst_req_0,
          ackL => binary_523_inst_ack_0,
          reqR => binary_523_inst_req_1,
          ackR => binary_523_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_528_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_524 & tmp_518;
      ret_val_x_x_buffer <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_528_inst_req_0,
          ackL => binary_528_inst_ack_0,
          reqR => binary_528_inst_req_1,
          ackR => binary_528_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_chk is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_chk;
architecture Default of ahir_glue_chk is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_chk_CP_1029_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_569_load_1_req_0 : boolean;
  signal binary_633_inst_req_0 : boolean;
  signal binary_588_inst_req_1 : boolean;
  signal binary_633_inst_ack_0 : boolean;
  signal ptr_deref_569_load_1_ack_0 : boolean;
  signal ptr_deref_985_addr_0_ack_0 : boolean;
  signal ptr_deref_1085_store_2_ack_1 : boolean;
  signal simple_obj_ref_653_inst_ack_0 : boolean;
  signal if_stmt_645_branch_req_0 : boolean;
  signal binary_677_inst_ack_0 : boolean;
  signal if_stmt_679_branch_ack_0 : boolean;
  signal ptr_deref_621_addr_3_req_0 : boolean;
  signal binary_639_inst_req_1 : boolean;
  signal simple_obj_ref_687_inst_req_0 : boolean;
  signal phi_stmt_847_req_0 : boolean;
  signal ptr_deref_569_load_0_ack_1 : boolean;
  signal binary_610_inst_ack_1 : boolean;
  signal ptr_deref_621_load_0_req_0 : boolean;
  signal type_cast_577_inst_ack_0 : boolean;
  signal ptr_deref_621_load_3_ack_0 : boolean;
  signal binary_582_inst_req_0 : boolean;
  signal ptr_deref_985_addr_0_req_0 : boolean;
  signal ptr_deref_621_load_3_ack_1 : boolean;
  signal ptr_deref_985_store_0_req_0 : boolean;
  signal binary_588_inst_ack_0 : boolean;
  signal type_cast_617_inst_req_0 : boolean;
  signal type_cast_617_inst_ack_0 : boolean;
  signal binary_633_inst_req_1 : boolean;
  signal ptr_deref_569_load_2_req_0 : boolean;
  signal binary_588_inst_ack_1 : boolean;
  signal binary_991_inst_req_1 : boolean;
  signal binary_1008_inst_req_1 : boolean;
  signal if_stmt_993_branch_req_0 : boolean;
  signal ptr_deref_621_load_3_req_0 : boolean;
  signal ptr_deref_985_gather_scatter_ack_0 : boolean;
  signal ptr_deref_985_root_address_inst_ack_0 : boolean;
  signal ptr_deref_621_addr_0_req_0 : boolean;
  signal ptr_deref_569_load_1_req_1 : boolean;
  signal binary_1092_inst_req_0 : boolean;
  signal ptr_deref_569_load_1_ack_1 : boolean;
  signal ptr_deref_621_addr_0_ack_0 : boolean;
  signal ptr_deref_1085_addr_0_req_1 : boolean;
  signal ptr_deref_1085_store_2_req_1 : boolean;
  signal ptr_deref_569_load_2_ack_0 : boolean;
  signal type_cast_850_inst_ack_0 : boolean;
  signal ptr_deref_621_addr_0_req_1 : boolean;
  signal ptr_deref_985_gather_scatter_req_0 : boolean;
  signal binary_633_inst_ack_1 : boolean;
  signal ptr_deref_621_addr_0_ack_1 : boolean;
  signal ptr_deref_1085_store_0_ack_1 : boolean;
  signal ptr_deref_1085_store_0_req_1 : boolean;
  signal binary_627_inst_ack_0 : boolean;
  signal if_stmt_993_branch_ack_0 : boolean;
  signal binary_610_inst_req_1 : boolean;
  signal ptr_deref_569_load_0_req_0 : boolean;
  signal ptr_deref_985_addr_3_req_1 : boolean;
  signal ptr_deref_569_load_2_req_1 : boolean;
  signal ptr_deref_621_addr_1_req_0 : boolean;
  signal ptr_deref_569_load_2_ack_1 : boolean;
  signal binary_1092_inst_ack_0 : boolean;
  signal ptr_deref_621_addr_1_ack_0 : boolean;
  signal binary_1092_inst_req_1 : boolean;
  signal ptr_deref_621_addr_1_req_1 : boolean;
  signal ptr_deref_621_addr_3_ack_1 : boolean;
  signal ptr_deref_569_load_3_req_0 : boolean;
  signal binary_665_inst_req_0 : boolean;
  signal ptr_deref_1085_addr_1_req_0 : boolean;
  signal ptr_deref_569_load_0_req_1 : boolean;
  signal binary_665_inst_req_1 : boolean;
  signal binary_656_inst_req_0 : boolean;
  signal ptr_deref_1085_store_3_req_1 : boolean;
  signal ptr_deref_569_load_3_req_1 : boolean;
  signal binary_665_inst_ack_1 : boolean;
  signal ptr_deref_1085_addr_0_ack_1 : boolean;
  signal binary_656_inst_ack_0 : boolean;
  signal if_stmt_599_branch_req_0 : boolean;
  signal binary_665_inst_ack_0 : boolean;
  signal ptr_deref_621_base_resize_req_0 : boolean;
  signal ptr_deref_569_load_3_ack_1 : boolean;
  signal ptr_deref_569_load_3_ack_0 : boolean;
  signal ptr_deref_621_addr_1_ack_1 : boolean;
  signal binary_656_inst_req_1 : boolean;
  signal ptr_deref_621_base_resize_ack_0 : boolean;
  signal ptr_deref_621_addr_2_req_0 : boolean;
  signal ptr_deref_569_gather_scatter_req_0 : boolean;
  signal type_cast_898_inst_req_0 : boolean;
  signal binary_656_inst_ack_1 : boolean;
  signal ptr_deref_569_gather_scatter_ack_0 : boolean;
  signal ptr_deref_621_addr_2_ack_0 : boolean;
  signal ptr_deref_1085_addr_1_ack_0 : boolean;
  signal ptr_deref_621_addr_2_req_1 : boolean;
  signal ptr_deref_985_addr_3_ack_1 : boolean;
  signal binary_627_inst_req_0 : boolean;
  signal binary_1092_inst_ack_1 : boolean;
  signal type_cast_850_inst_req_0 : boolean;
  signal type_cast_573_inst_req_0 : boolean;
  signal type_cast_573_inst_ack_0 : boolean;
  signal if_stmt_599_branch_ack_0 : boolean;
  signal simple_obj_ref_607_inst_req_0 : boolean;
  signal ptr_deref_621_load_1_req_1 : boolean;
  signal ptr_deref_1085_root_address_inst_ack_0 : boolean;
  signal ptr_deref_621_gather_scatter_req_0 : boolean;
  signal binary_639_inst_ack_0 : boolean;
  signal binary_671_inst_req_1 : boolean;
  signal ptr_deref_621_addr_3_ack_0 : boolean;
  signal binary_627_inst_req_1 : boolean;
  signal ptr_deref_1085_base_resize_req_0 : boolean;
  signal type_cast_643_inst_req_0 : boolean;
  signal ptr_deref_1085_root_address_inst_req_0 : boolean;
  signal binary_610_inst_req_0 : boolean;
  signal simple_obj_ref_687_inst_ack_0 : boolean;
  signal ptr_deref_621_load_0_req_1 : boolean;
  signal binary_627_inst_ack_1 : boolean;
  signal binary_639_inst_ack_1 : boolean;
  signal ptr_deref_621_load_2_req_1 : boolean;
  signal ptr_deref_985_addr_3_ack_0 : boolean;
  signal binary_991_inst_ack_0 : boolean;
  signal binary_677_inst_req_1 : boolean;
  signal ptr_deref_569_load_0_ack_0 : boolean;
  signal ptr_deref_621_load_2_ack_1 : boolean;
  signal ptr_deref_621_load_3_req_1 : boolean;
  signal ptr_deref_621_load_0_ack_1 : boolean;
  signal if_stmt_993_branch_ack_1 : boolean;
  signal binary_588_inst_req_0 : boolean;
  signal binary_610_inst_ack_0 : boolean;
  signal ptr_deref_621_addr_3_req_1 : boolean;
  signal phi_stmt_754_req_1 : boolean;
  signal ptr_deref_1085_addr_1_req_1 : boolean;
  signal binary_597_inst_ack_1 : boolean;
  signal if_stmt_679_branch_req_0 : boolean;
  signal binary_1008_inst_ack_1 : boolean;
  signal type_cast_760_inst_req_0 : boolean;
  signal ptr_deref_621_load_2_ack_0 : boolean;
  signal binary_582_inst_ack_1 : boolean;
  signal ptr_deref_621_load_0_ack_0 : boolean;
  signal simple_obj_ref_653_inst_req_0 : boolean;
  signal binary_671_inst_req_0 : boolean;
  signal binary_582_inst_req_1 : boolean;
  signal binary_582_inst_ack_0 : boolean;
  signal ptr_deref_985_addr_3_req_0 : boolean;
  signal phi_stmt_895_req_1 : boolean;
  signal type_cast_898_inst_ack_0 : boolean;
  signal binary_677_inst_ack_1 : boolean;
  signal binary_671_inst_ack_1 : boolean;
  signal binary_690_inst_ack_0 : boolean;
  signal binary_690_inst_req_1 : boolean;
  signal ptr_deref_1085_addr_2_ack_0 : boolean;
  signal if_stmt_645_branch_ack_1 : boolean;
  signal ptr_deref_621_load_1_req_0 : boolean;
  signal ptr_deref_621_load_1_ack_0 : boolean;
  signal if_stmt_599_branch_ack_1 : boolean;
  signal type_cast_643_inst_ack_0 : boolean;
  signal ptr_deref_621_root_address_inst_req_0 : boolean;
  signal call_stmt_697_call_ack_0 : boolean;
  signal ptr_deref_1085_addr_0_ack_0 : boolean;
  signal if_stmt_1094_branch_req_0 : boolean;
  signal if_stmt_679_branch_ack_1 : boolean;
  signal ptr_deref_1085_addr_2_req_0 : boolean;
  signal binary_690_inst_ack_1 : boolean;
  signal call_stmt_697_call_req_0 : boolean;
  signal ptr_deref_1085_base_resize_ack_0 : boolean;
  signal type_cast_593_inst_req_0 : boolean;
  signal ptr_deref_621_addr_2_ack_1 : boolean;
  signal ptr_deref_985_addr_2_ack_1 : boolean;
  signal ptr_deref_1085_store_3_ack_1 : boolean;
  signal type_cast_593_inst_ack_0 : boolean;
  signal ptr_deref_621_load_2_req_0 : boolean;
  signal ptr_deref_621_root_address_inst_ack_0 : boolean;
  signal binary_639_inst_req_0 : boolean;
  signal binary_671_inst_ack_0 : boolean;
  signal ptr_deref_1085_addr_1_ack_1 : boolean;
  signal binary_677_inst_req_0 : boolean;
  signal call_stmt_697_call_ack_1 : boolean;
  signal binary_597_inst_req_0 : boolean;
  signal simple_obj_ref_607_inst_ack_0 : boolean;
  signal ptr_deref_621_gather_scatter_ack_0 : boolean;
  signal ptr_deref_621_load_1_ack_1 : boolean;
  signal if_stmt_645_branch_ack_0 : boolean;
  signal binary_991_inst_ack_1 : boolean;
  signal type_cast_700_inst_req_0 : boolean;
  signal type_cast_700_inst_ack_0 : boolean;
  signal binary_710_inst_req_1 : boolean;
  signal binary_710_inst_ack_1 : boolean;
  signal ptr_deref_1085_addr_2_ack_1 : boolean;
  signal binary_710_inst_req_0 : boolean;
  signal binary_710_inst_ack_0 : boolean;
  signal type_cast_767_inst_req_0 : boolean;
  signal type_cast_767_inst_ack_0 : boolean;
  signal binary_705_inst_req_0 : boolean;
  signal binary_705_inst_ack_0 : boolean;
  signal if_stmt_1094_branch_ack_1 : boolean;
  signal ptr_deref_1085_addr_2_req_1 : boolean;
  signal if_stmt_1094_branch_ack_0 : boolean;
  signal call_stmt_697_call_req_1 : boolean;
  signal binary_690_inst_req_0 : boolean;
  signal binary_597_inst_ack_0 : boolean;
  signal binary_597_inst_req_1 : boolean;
  signal binary_705_inst_req_1 : boolean;
  signal binary_705_inst_ack_1 : boolean;
  signal type_cast_760_inst_ack_0 : boolean;
  signal phi_stmt_761_req_1 : boolean;
  signal ptr_deref_1085_store_1_ack_1 : boolean;
  signal ptr_deref_985_store_0_ack_0 : boolean;
  signal ptr_deref_1085_addr_0_req_0 : boolean;
  signal type_cast_577_inst_req_0 : boolean;
  signal ptr_deref_985_addr_0_req_1 : boolean;
  signal ptr_deref_985_store_1_req_0 : boolean;
  signal ptr_deref_985_store_1_ack_0 : boolean;
  signal ptr_deref_985_addr_0_ack_1 : boolean;
  signal ptr_deref_1085_store_1_req_1 : boolean;
  signal array_obj_ref_1024_index_0_resize_req_0 : boolean;
  signal ternary_1014_inst_req_0 : boolean;
  signal ptr_deref_985_store_2_req_0 : boolean;
  signal array_obj_ref_1024_offset_inst_req_0 : boolean;
  signal array_obj_ref_1024_index_0_rename_ack_0 : boolean;
  signal binary_1020_inst_ack_1 : boolean;
  signal array_obj_ref_1024_index_0_rename_req_0 : boolean;
  signal ptr_deref_985_store_2_ack_0 : boolean;
  signal array_obj_ref_1024_index_0_resize_ack_0 : boolean;
  signal ternary_1014_inst_ack_0 : boolean;
  signal ptr_deref_985_store_3_req_0 : boolean;
  signal ptr_deref_985_store_3_ack_0 : boolean;
  signal ptr_deref_985_store_0_req_1 : boolean;
  signal ptr_deref_985_store_0_ack_1 : boolean;
  signal binary_1003_inst_req_0 : boolean;
  signal ptr_deref_985_base_resize_req_0 : boolean;
  signal binary_1003_inst_ack_0 : boolean;
  signal ptr_deref_985_addr_1_req_0 : boolean;
  signal simple_obj_ref_537_inst_req_0 : boolean;
  signal binary_1003_inst_req_1 : boolean;
  signal simple_obj_ref_537_inst_ack_0 : boolean;
  signal binary_1003_inst_ack_1 : boolean;
  signal ptr_deref_985_addr_1_ack_0 : boolean;
  signal type_cast_538_inst_req_0 : boolean;
  signal type_cast_538_inst_ack_0 : boolean;
  signal ptr_deref_985_addr_1_req_1 : boolean;
  signal ptr_deref_985_base_resize_ack_0 : boolean;
  signal ptr_deref_985_addr_1_ack_1 : boolean;
  signal ptr_deref_985_store_1_req_1 : boolean;
  signal type_cast_542_inst_req_0 : boolean;
  signal ptr_deref_985_store_1_ack_1 : boolean;
  signal type_cast_542_inst_ack_0 : boolean;
  signal ptr_deref_985_store_2_req_1 : boolean;
  signal ptr_deref_985_store_2_ack_1 : boolean;
  signal ptr_deref_985_store_3_req_1 : boolean;
  signal ptr_deref_985_store_3_ack_1 : boolean;
  signal array_obj_ref_549_base_resize_req_0 : boolean;
  signal array_obj_ref_549_base_resize_ack_0 : boolean;
  signal array_obj_ref_549_root_address_inst_req_0 : boolean;
  signal array_obj_ref_549_root_address_inst_ack_0 : boolean;
  signal binary_1008_inst_req_0 : boolean;
  signal array_obj_ref_549_root_address_inst_req_1 : boolean;
  signal array_obj_ref_549_root_address_inst_ack_1 : boolean;
  signal ptr_deref_985_addr_2_req_0 : boolean;
  signal array_obj_ref_549_final_reg_req_0 : boolean;
  signal array_obj_ref_549_final_reg_ack_0 : boolean;
  signal binary_1020_inst_req_0 : boolean;
  signal binary_1020_inst_ack_0 : boolean;
  signal ptr_deref_985_addr_2_ack_0 : boolean;
  signal binary_1008_inst_ack_0 : boolean;
  signal ptr_deref_985_root_address_inst_req_0 : boolean;
  signal binary_1020_inst_req_1 : boolean;
  signal ptr_deref_985_addr_2_req_1 : boolean;
  signal binary_991_inst_req_0 : boolean;
  signal ptr_deref_553_base_resize_req_0 : boolean;
  signal ptr_deref_553_base_resize_ack_0 : boolean;
  signal ptr_deref_553_root_address_inst_req_0 : boolean;
  signal ptr_deref_553_root_address_inst_ack_0 : boolean;
  signal ptr_deref_553_addr_0_req_0 : boolean;
  signal ptr_deref_553_addr_0_ack_0 : boolean;
  signal ptr_deref_553_addr_0_req_1 : boolean;
  signal ptr_deref_553_addr_0_ack_1 : boolean;
  signal ptr_deref_553_addr_1_req_0 : boolean;
  signal ptr_deref_553_addr_1_ack_0 : boolean;
  signal ptr_deref_553_addr_1_req_1 : boolean;
  signal ptr_deref_553_addr_1_ack_1 : boolean;
  signal ptr_deref_553_addr_2_req_0 : boolean;
  signal ptr_deref_553_addr_2_ack_0 : boolean;
  signal ptr_deref_553_addr_2_req_1 : boolean;
  signal ptr_deref_553_addr_2_ack_1 : boolean;
  signal ptr_deref_553_addr_3_req_0 : boolean;
  signal ptr_deref_553_addr_3_ack_0 : boolean;
  signal ptr_deref_553_addr_3_req_1 : boolean;
  signal ptr_deref_553_addr_3_ack_1 : boolean;
  signal ptr_deref_553_load_0_req_0 : boolean;
  signal ptr_deref_553_load_0_ack_0 : boolean;
  signal ptr_deref_553_load_1_req_0 : boolean;
  signal ptr_deref_553_load_1_ack_0 : boolean;
  signal ptr_deref_553_load_2_req_0 : boolean;
  signal ptr_deref_553_load_2_ack_0 : boolean;
  signal ptr_deref_553_load_3_req_0 : boolean;
  signal ptr_deref_553_load_3_ack_0 : boolean;
  signal ptr_deref_553_load_0_req_1 : boolean;
  signal ptr_deref_553_load_0_ack_1 : boolean;
  signal ptr_deref_553_load_1_req_1 : boolean;
  signal ptr_deref_553_load_1_ack_1 : boolean;
  signal ptr_deref_553_load_2_req_1 : boolean;
  signal ptr_deref_553_load_2_ack_1 : boolean;
  signal ptr_deref_553_load_3_req_1 : boolean;
  signal ptr_deref_553_load_3_ack_1 : boolean;
  signal ptr_deref_553_gather_scatter_req_0 : boolean;
  signal ptr_deref_553_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_558_base_resize_req_0 : boolean;
  signal array_obj_ref_558_base_resize_ack_0 : boolean;
  signal array_obj_ref_558_root_address_inst_req_0 : boolean;
  signal array_obj_ref_558_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_558_root_address_inst_req_1 : boolean;
  signal array_obj_ref_558_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_558_final_reg_req_0 : boolean;
  signal array_obj_ref_558_final_reg_ack_0 : boolean;
  signal array_obj_ref_565_base_resize_req_0 : boolean;
  signal array_obj_ref_565_base_resize_ack_0 : boolean;
  signal array_obj_ref_565_root_address_inst_req_0 : boolean;
  signal array_obj_ref_565_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_565_root_address_inst_req_1 : boolean;
  signal array_obj_ref_565_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_565_final_reg_req_0 : boolean;
  signal array_obj_ref_565_final_reg_ack_0 : boolean;
  signal ptr_deref_569_base_resize_req_0 : boolean;
  signal ptr_deref_569_base_resize_ack_0 : boolean;
  signal ptr_deref_569_root_address_inst_req_0 : boolean;
  signal ptr_deref_569_root_address_inst_ack_0 : boolean;
  signal ptr_deref_569_addr_0_req_0 : boolean;
  signal ptr_deref_569_addr_0_ack_0 : boolean;
  signal ptr_deref_569_addr_0_req_1 : boolean;
  signal ptr_deref_569_addr_0_ack_1 : boolean;
  signal ptr_deref_569_addr_1_req_0 : boolean;
  signal ptr_deref_569_addr_1_ack_0 : boolean;
  signal ptr_deref_569_addr_1_req_1 : boolean;
  signal ptr_deref_569_addr_1_ack_1 : boolean;
  signal ptr_deref_569_addr_2_req_0 : boolean;
  signal ptr_deref_569_addr_2_ack_0 : boolean;
  signal ptr_deref_569_addr_2_req_1 : boolean;
  signal ptr_deref_569_addr_2_ack_1 : boolean;
  signal ptr_deref_569_addr_3_req_0 : boolean;
  signal ptr_deref_569_addr_3_ack_0 : boolean;
  signal ptr_deref_569_addr_3_req_1 : boolean;
  signal ptr_deref_569_addr_3_ack_1 : boolean;
  signal binary_715_inst_req_0 : boolean;
  signal binary_715_inst_ack_0 : boolean;
  signal binary_715_inst_req_1 : boolean;
  signal binary_715_inst_ack_1 : boolean;
  signal phi_stmt_847_ack_0 : boolean;
  signal if_stmt_717_branch_req_0 : boolean;
  signal if_stmt_717_branch_ack_1 : boolean;
  signal phi_stmt_895_req_0 : boolean;
  signal phi_stmt_754_req_0 : boolean;
  signal if_stmt_717_branch_ack_0 : boolean;
  signal ptr_deref_1085_addr_3_req_0 : boolean;
  signal ptr_deref_1085_addr_3_ack_0 : boolean;
  signal binary_728_inst_req_0 : boolean;
  signal type_cast_857_inst_req_0 : boolean;
  signal binary_728_inst_ack_0 : boolean;
  signal ptr_deref_1085_addr_3_req_1 : boolean;
  signal binary_728_inst_req_1 : boolean;
  signal ptr_deref_1085_addr_3_ack_1 : boolean;
  signal binary_728_inst_ack_1 : boolean;
  signal simple_obj_ref_725_inst_req_0 : boolean;
  signal simple_obj_ref_725_inst_ack_0 : boolean;
  signal binary_737_inst_req_0 : boolean;
  signal binary_737_inst_ack_0 : boolean;
  signal binary_737_inst_req_1 : boolean;
  signal binary_737_inst_ack_1 : boolean;
  signal type_cast_857_inst_ack_0 : boolean;
  signal phi_stmt_854_ack_0 : boolean;
  signal if_stmt_739_branch_req_0 : boolean;
  signal if_stmt_739_branch_ack_1 : boolean;
  signal if_stmt_739_branch_ack_0 : boolean;
  signal phi_stmt_761_req_0 : boolean;
  signal phi_stmt_895_ack_0 : boolean;
  signal binary_750_inst_req_0 : boolean;
  signal binary_750_inst_ack_0 : boolean;
  signal binary_750_inst_req_1 : boolean;
  signal ptr_deref_1085_gather_scatter_req_0 : boolean;
  signal binary_750_inst_ack_1 : boolean;
  signal ptr_deref_1085_gather_scatter_ack_0 : boolean;
  signal phi_stmt_754_ack_0 : boolean;
  signal phi_stmt_761_ack_0 : boolean;
  signal binary_773_inst_req_0 : boolean;
  signal binary_773_inst_ack_0 : boolean;
  signal binary_773_inst_req_1 : boolean;
  signal binary_773_inst_ack_1 : boolean;
  signal ptr_deref_1085_store_0_req_0 : boolean;
  signal type_cast_900_inst_req_0 : boolean;
  signal binary_778_inst_req_0 : boolean;
  signal binary_778_inst_ack_0 : boolean;
  signal binary_778_inst_req_1 : boolean;
  signal ptr_deref_1085_store_0_ack_0 : boolean;
  signal binary_778_inst_ack_1 : boolean;
  signal phi_stmt_860_ack_0 : boolean;
  signal type_cast_1103_inst_req_0 : boolean;
  signal type_cast_1103_inst_ack_0 : boolean;
  signal binary_784_inst_req_0 : boolean;
  signal binary_784_inst_ack_0 : boolean;
  signal binary_784_inst_req_1 : boolean;
  signal binary_784_inst_ack_1 : boolean;
  signal binary_790_inst_req_0 : boolean;
  signal binary_790_inst_ack_0 : boolean;
  signal binary_790_inst_req_1 : boolean;
  signal binary_790_inst_ack_1 : boolean;
  signal phi_stmt_854_req_0 : boolean;
  signal array_obj_ref_794_index_0_resize_req_0 : boolean;
  signal array_obj_ref_794_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_794_index_0_rename_req_0 : boolean;
  signal array_obj_ref_794_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_794_offset_inst_req_0 : boolean;
  signal array_obj_ref_794_offset_inst_ack_0 : boolean;
  signal array_obj_ref_794_base_resize_req_0 : boolean;
  signal array_obj_ref_794_base_resize_ack_0 : boolean;
  signal ptr_deref_1085_store_1_req_0 : boolean;
  signal array_obj_ref_794_root_address_inst_req_0 : boolean;
  signal phi_stmt_847_req_1 : boolean;
  signal array_obj_ref_794_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_794_root_address_inst_req_1 : boolean;
  signal array_obj_ref_794_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1085_store_1_ack_0 : boolean;
  signal array_obj_ref_794_final_reg_req_0 : boolean;
  signal array_obj_ref_794_final_reg_ack_0 : boolean;
  signal type_cast_1107_inst_req_0 : boolean;
  signal type_cast_799_inst_req_0 : boolean;
  signal type_cast_1107_inst_ack_0 : boolean;
  signal type_cast_799_inst_ack_0 : boolean;
  signal ptr_deref_803_base_resize_req_0 : boolean;
  signal type_cast_863_inst_req_0 : boolean;
  signal ptr_deref_803_base_resize_ack_0 : boolean;
  signal type_cast_859_inst_req_0 : boolean;
  signal ptr_deref_1085_store_2_req_0 : boolean;
  signal ptr_deref_803_root_address_inst_req_0 : boolean;
  signal ptr_deref_803_root_address_inst_ack_0 : boolean;
  signal type_cast_859_inst_ack_0 : boolean;
  signal ptr_deref_803_addr_0_req_0 : boolean;
  signal ptr_deref_803_addr_0_ack_0 : boolean;
  signal phi_stmt_854_req_1 : boolean;
  signal ptr_deref_803_addr_0_req_1 : boolean;
  signal ptr_deref_803_addr_0_ack_1 : boolean;
  signal ptr_deref_803_addr_1_req_0 : boolean;
  signal type_cast_863_inst_ack_0 : boolean;
  signal ptr_deref_803_addr_1_ack_0 : boolean;
  signal ptr_deref_803_addr_1_req_1 : boolean;
  signal ptr_deref_1085_store_2_ack_0 : boolean;
  signal ptr_deref_803_addr_1_ack_1 : boolean;
  signal ptr_deref_803_load_0_req_0 : boolean;
  signal ptr_deref_803_load_0_ack_0 : boolean;
  signal ptr_deref_803_load_1_req_0 : boolean;
  signal ptr_deref_803_load_1_ack_0 : boolean;
  signal ptr_deref_803_load_0_req_1 : boolean;
  signal ptr_deref_803_load_0_ack_1 : boolean;
  signal ptr_deref_1085_store_3_req_0 : boolean;
  signal ptr_deref_803_load_1_req_1 : boolean;
  signal ptr_deref_803_load_1_ack_1 : boolean;
  signal ptr_deref_803_gather_scatter_req_0 : boolean;
  signal ptr_deref_1085_store_3_ack_0 : boolean;
  signal ptr_deref_803_gather_scatter_ack_0 : boolean;
  signal type_cast_807_inst_req_0 : boolean;
  signal type_cast_807_inst_ack_0 : boolean;
  signal simple_obj_ref_1105_inst_req_0 : boolean;
  signal simple_obj_ref_1105_inst_ack_0 : boolean;
  signal binary_812_inst_req_0 : boolean;
  signal binary_812_inst_ack_0 : boolean;
  signal binary_812_inst_req_1 : boolean;
  signal binary_812_inst_ack_1 : boolean;
  signal phi_stmt_860_req_0 : boolean;
  signal type_cast_865_inst_req_0 : boolean;
  signal type_cast_900_inst_ack_0 : boolean;
  signal type_cast_816_inst_req_0 : boolean;
  signal type_cast_865_inst_ack_0 : boolean;
  signal type_cast_816_inst_ack_0 : boolean;
  signal binary_820_inst_req_0 : boolean;
  signal binary_820_inst_ack_0 : boolean;
  signal binary_820_inst_req_1 : boolean;
  signal binary_820_inst_ack_1 : boolean;
  signal phi_stmt_860_req_1 : boolean;
  signal binary_826_inst_req_0 : boolean;
  signal binary_826_inst_ack_0 : boolean;
  signal binary_826_inst_req_1 : boolean;
  signal binary_826_inst_ack_1 : boolean;
  signal if_stmt_828_branch_req_0 : boolean;
  signal if_stmt_828_branch_ack_1 : boolean;
  signal if_stmt_828_branch_ack_0 : boolean;
  signal binary_839_inst_req_0 : boolean;
  signal binary_839_inst_ack_0 : boolean;
  signal binary_839_inst_req_1 : boolean;
  signal binary_839_inst_ack_1 : boolean;
  signal array_obj_ref_843_index_0_resize_req_0 : boolean;
  signal array_obj_ref_843_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_843_index_0_rename_req_0 : boolean;
  signal array_obj_ref_843_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_843_offset_inst_req_0 : boolean;
  signal array_obj_ref_843_offset_inst_ack_0 : boolean;
  signal array_obj_ref_843_base_resize_req_0 : boolean;
  signal array_obj_ref_843_base_resize_ack_0 : boolean;
  signal array_obj_ref_843_root_address_inst_req_0 : boolean;
  signal array_obj_ref_843_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_843_root_address_inst_req_1 : boolean;
  signal array_obj_ref_843_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_843_final_reg_req_0 : boolean;
  signal array_obj_ref_843_final_reg_ack_0 : boolean;
  signal binary_871_inst_req_0 : boolean;
  signal binary_871_inst_ack_0 : boolean;
  signal binary_871_inst_req_1 : boolean;
  signal binary_871_inst_ack_1 : boolean;
  signal if_stmt_873_branch_req_0 : boolean;
  signal if_stmt_873_branch_ack_1 : boolean;
  signal if_stmt_873_branch_ack_0 : boolean;
  signal ptr_deref_882_base_resize_req_0 : boolean;
  signal ptr_deref_882_base_resize_ack_0 : boolean;
  signal ptr_deref_882_root_address_inst_req_0 : boolean;
  signal ptr_deref_882_root_address_inst_ack_0 : boolean;
  signal ptr_deref_882_addr_0_req_0 : boolean;
  signal ptr_deref_882_addr_0_ack_0 : boolean;
  signal ptr_deref_882_load_0_req_0 : boolean;
  signal ptr_deref_882_load_0_ack_0 : boolean;
  signal ptr_deref_882_load_0_req_1 : boolean;
  signal ptr_deref_882_load_0_ack_1 : boolean;
  signal ptr_deref_882_gather_scatter_req_0 : boolean;
  signal ptr_deref_882_gather_scatter_ack_0 : boolean;
  signal type_cast_886_inst_req_0 : boolean;
  signal type_cast_886_inst_ack_0 : boolean;
  signal binary_891_inst_req_0 : boolean;
  signal binary_891_inst_ack_0 : boolean;
  signal binary_891_inst_req_1 : boolean;
  signal binary_891_inst_ack_1 : boolean;
  signal binary_906_inst_req_0 : boolean;
  signal binary_906_inst_ack_0 : boolean;
  signal binary_906_inst_req_1 : boolean;
  signal binary_906_inst_ack_1 : boolean;
  signal binary_912_inst_req_0 : boolean;
  signal binary_912_inst_ack_0 : boolean;
  signal binary_912_inst_req_1 : boolean;
  signal binary_912_inst_ack_1 : boolean;
  signal binary_917_inst_req_0 : boolean;
  signal binary_917_inst_ack_0 : boolean;
  signal binary_917_inst_req_1 : boolean;
  signal binary_917_inst_ack_1 : boolean;
  signal binary_923_inst_req_0 : boolean;
  signal binary_923_inst_ack_0 : boolean;
  signal binary_923_inst_req_1 : boolean;
  signal binary_923_inst_ack_1 : boolean;
  signal binary_928_inst_req_0 : boolean;
  signal binary_928_inst_ack_0 : boolean;
  signal binary_928_inst_req_1 : boolean;
  signal binary_928_inst_ack_1 : boolean;
  signal type_cast_932_inst_req_0 : boolean;
  signal type_cast_932_inst_ack_0 : boolean;
  signal binary_938_inst_req_0 : boolean;
  signal binary_938_inst_ack_0 : boolean;
  signal binary_938_inst_req_1 : boolean;
  signal binary_938_inst_ack_1 : boolean;
  signal if_stmt_940_branch_req_0 : boolean;
  signal if_stmt_940_branch_ack_1 : boolean;
  signal if_stmt_940_branch_ack_0 : boolean;
  signal binary_951_inst_req_0 : boolean;
  signal binary_951_inst_ack_0 : boolean;
  signal binary_951_inst_req_1 : boolean;
  signal binary_951_inst_ack_1 : boolean;
  signal simple_obj_ref_948_inst_req_0 : boolean;
  signal simple_obj_ref_948_inst_ack_0 : boolean;
  signal array_obj_ref_961_base_resize_req_0 : boolean;
  signal array_obj_ref_961_base_resize_ack_0 : boolean;
  signal array_obj_ref_961_root_address_inst_req_0 : boolean;
  signal array_obj_ref_961_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_961_root_address_inst_req_1 : boolean;
  signal array_obj_ref_961_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_961_final_reg_req_0 : boolean;
  signal array_obj_ref_961_final_reg_ack_0 : boolean;
  signal ptr_deref_964_base_resize_req_0 : boolean;
  signal ptr_deref_964_base_resize_ack_0 : boolean;
  signal ptr_deref_964_root_address_inst_req_0 : boolean;
  signal ptr_deref_964_root_address_inst_ack_0 : boolean;
  signal ptr_deref_964_addr_0_req_0 : boolean;
  signal ptr_deref_964_addr_0_ack_0 : boolean;
  signal ptr_deref_964_addr_0_req_1 : boolean;
  signal ptr_deref_964_addr_0_ack_1 : boolean;
  signal ptr_deref_964_addr_1_req_0 : boolean;
  signal ptr_deref_964_addr_1_ack_0 : boolean;
  signal ptr_deref_964_addr_1_req_1 : boolean;
  signal ptr_deref_964_addr_1_ack_1 : boolean;
  signal ptr_deref_964_addr_2_req_0 : boolean;
  signal ptr_deref_964_addr_2_ack_0 : boolean;
  signal ptr_deref_964_addr_2_req_1 : boolean;
  signal ptr_deref_964_addr_2_ack_1 : boolean;
  signal ptr_deref_964_addr_3_req_0 : boolean;
  signal ptr_deref_964_addr_3_ack_0 : boolean;
  signal ptr_deref_964_addr_3_req_1 : boolean;
  signal ptr_deref_964_addr_3_ack_1 : boolean;
  signal ptr_deref_964_gather_scatter_req_0 : boolean;
  signal ptr_deref_964_gather_scatter_ack_0 : boolean;
  signal ptr_deref_964_store_0_req_0 : boolean;
  signal ptr_deref_964_store_0_ack_0 : boolean;
  signal ptr_deref_964_store_1_req_0 : boolean;
  signal ptr_deref_964_store_1_ack_0 : boolean;
  signal ptr_deref_964_store_2_req_0 : boolean;
  signal ptr_deref_964_store_2_ack_0 : boolean;
  signal ptr_deref_964_store_3_req_0 : boolean;
  signal ptr_deref_964_store_3_ack_0 : boolean;
  signal ptr_deref_964_store_0_req_1 : boolean;
  signal ptr_deref_964_store_0_ack_1 : boolean;
  signal ptr_deref_964_store_1_req_1 : boolean;
  signal ptr_deref_964_store_1_ack_1 : boolean;
  signal ptr_deref_964_store_2_req_1 : boolean;
  signal ptr_deref_964_store_2_ack_1 : boolean;
  signal ptr_deref_964_store_3_req_1 : boolean;
  signal ptr_deref_964_store_3_ack_1 : boolean;
  signal binary_971_inst_req_0 : boolean;
  signal binary_971_inst_ack_0 : boolean;
  signal binary_971_inst_req_1 : boolean;
  signal binary_971_inst_ack_1 : boolean;
  signal array_obj_ref_975_index_0_resize_req_0 : boolean;
  signal array_obj_ref_975_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_975_index_0_rename_req_0 : boolean;
  signal array_obj_ref_975_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_975_offset_inst_req_0 : boolean;
  signal array_obj_ref_975_offset_inst_ack_0 : boolean;
  signal array_obj_ref_975_base_resize_req_0 : boolean;
  signal array_obj_ref_975_base_resize_ack_0 : boolean;
  signal array_obj_ref_975_root_address_inst_req_0 : boolean;
  signal array_obj_ref_975_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_975_root_address_inst_req_1 : boolean;
  signal array_obj_ref_975_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_975_final_reg_req_0 : boolean;
  signal array_obj_ref_975_final_reg_ack_0 : boolean;
  signal array_obj_ref_982_base_resize_req_0 : boolean;
  signal array_obj_ref_982_base_resize_ack_0 : boolean;
  signal array_obj_ref_982_root_address_inst_req_0 : boolean;
  signal array_obj_ref_982_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_982_root_address_inst_req_1 : boolean;
  signal array_obj_ref_982_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_982_final_reg_req_0 : boolean;
  signal array_obj_ref_982_final_reg_ack_0 : boolean;
  signal array_obj_ref_1024_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1024_base_resize_req_0 : boolean;
  signal array_obj_ref_1024_base_resize_ack_0 : boolean;
  signal array_obj_ref_1024_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1024_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1024_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1024_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1024_final_reg_req_0 : boolean;
  signal array_obj_ref_1024_final_reg_ack_0 : boolean;
  signal ptr_deref_1027_base_resize_req_0 : boolean;
  signal ptr_deref_1027_base_resize_ack_0 : boolean;
  signal ptr_deref_1027_root_address_inst_req_0 : boolean;
  signal ptr_deref_1027_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1027_addr_0_req_0 : boolean;
  signal ptr_deref_1027_addr_0_ack_0 : boolean;
  signal ptr_deref_1027_addr_0_req_1 : boolean;
  signal ptr_deref_1027_addr_0_ack_1 : boolean;
  signal ptr_deref_1027_addr_1_req_0 : boolean;
  signal ptr_deref_1027_addr_1_ack_0 : boolean;
  signal ptr_deref_1027_addr_1_req_1 : boolean;
  signal ptr_deref_1027_addr_1_ack_1 : boolean;
  signal ptr_deref_1027_addr_2_req_0 : boolean;
  signal ptr_deref_1027_addr_2_ack_0 : boolean;
  signal ptr_deref_1027_addr_2_req_1 : boolean;
  signal ptr_deref_1027_addr_2_ack_1 : boolean;
  signal ptr_deref_1027_addr_3_req_0 : boolean;
  signal ptr_deref_1027_addr_3_ack_0 : boolean;
  signal ptr_deref_1027_addr_3_req_1 : boolean;
  signal ptr_deref_1027_addr_3_ack_1 : boolean;
  signal ptr_deref_1027_gather_scatter_req_0 : boolean;
  signal ptr_deref_1027_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1027_store_0_req_0 : boolean;
  signal ptr_deref_1027_store_0_ack_0 : boolean;
  signal ptr_deref_1027_store_1_req_0 : boolean;
  signal ptr_deref_1027_store_1_ack_0 : boolean;
  signal ptr_deref_1027_store_2_req_0 : boolean;
  signal ptr_deref_1027_store_2_ack_0 : boolean;
  signal ptr_deref_1027_store_3_req_0 : boolean;
  signal ptr_deref_1027_store_3_ack_0 : boolean;
  signal ptr_deref_1027_store_0_req_1 : boolean;
  signal ptr_deref_1027_store_0_ack_1 : boolean;
  signal ptr_deref_1027_store_1_req_1 : boolean;
  signal ptr_deref_1027_store_1_ack_1 : boolean;
  signal ptr_deref_1027_store_2_req_1 : boolean;
  signal ptr_deref_1027_store_2_ack_1 : boolean;
  signal ptr_deref_1027_store_3_req_1 : boolean;
  signal ptr_deref_1027_store_3_ack_1 : boolean;
  signal array_obj_ref_1033_base_resize_req_0 : boolean;
  signal array_obj_ref_1033_base_resize_ack_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1033_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1033_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1033_final_reg_req_0 : boolean;
  signal array_obj_ref_1033_final_reg_ack_0 : boolean;
  signal type_cast_1037_inst_req_0 : boolean;
  signal type_cast_1037_inst_ack_0 : boolean;
  signal ptr_deref_1041_base_resize_req_0 : boolean;
  signal ptr_deref_1041_base_resize_ack_0 : boolean;
  signal ptr_deref_1041_root_address_inst_req_0 : boolean;
  signal ptr_deref_1041_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1041_addr_0_req_0 : boolean;
  signal ptr_deref_1041_addr_0_ack_0 : boolean;
  signal ptr_deref_1041_addr_0_req_1 : boolean;
  signal ptr_deref_1041_addr_0_ack_1 : boolean;
  signal ptr_deref_1041_addr_1_req_0 : boolean;
  signal ptr_deref_1041_addr_1_ack_0 : boolean;
  signal ptr_deref_1041_addr_1_req_1 : boolean;
  signal ptr_deref_1041_addr_1_ack_1 : boolean;
  signal ptr_deref_1041_addr_2_req_0 : boolean;
  signal ptr_deref_1041_addr_2_ack_0 : boolean;
  signal ptr_deref_1041_addr_2_req_1 : boolean;
  signal ptr_deref_1041_addr_2_ack_1 : boolean;
  signal ptr_deref_1041_addr_3_req_0 : boolean;
  signal ptr_deref_1041_addr_3_ack_0 : boolean;
  signal ptr_deref_1041_addr_3_req_1 : boolean;
  signal ptr_deref_1041_addr_3_ack_1 : boolean;
  signal ptr_deref_1041_load_0_req_0 : boolean;
  signal ptr_deref_1041_load_0_ack_0 : boolean;
  signal ptr_deref_1041_load_1_req_0 : boolean;
  signal ptr_deref_1041_load_1_ack_0 : boolean;
  signal ptr_deref_1041_load_2_req_0 : boolean;
  signal ptr_deref_1041_load_2_ack_0 : boolean;
  signal ptr_deref_1041_load_3_req_0 : boolean;
  signal ptr_deref_1041_load_3_ack_0 : boolean;
  signal ptr_deref_1041_load_0_req_1 : boolean;
  signal ptr_deref_1041_load_0_ack_1 : boolean;
  signal ptr_deref_1041_load_1_req_1 : boolean;
  signal ptr_deref_1041_load_1_ack_1 : boolean;
  signal ptr_deref_1041_load_2_req_1 : boolean;
  signal ptr_deref_1041_load_2_ack_1 : boolean;
  signal ptr_deref_1041_load_3_req_1 : boolean;
  signal ptr_deref_1041_load_3_ack_1 : boolean;
  signal ptr_deref_1041_gather_scatter_req_0 : boolean;
  signal ptr_deref_1041_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1048_base_resize_req_0 : boolean;
  signal array_obj_ref_1048_base_resize_ack_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1048_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1048_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1048_final_reg_req_0 : boolean;
  signal array_obj_ref_1048_final_reg_ack_0 : boolean;
  signal type_cast_1052_inst_req_0 : boolean;
  signal type_cast_1052_inst_ack_0 : boolean;
  signal ptr_deref_1055_base_resize_req_0 : boolean;
  signal ptr_deref_1055_base_resize_ack_0 : boolean;
  signal ptr_deref_1055_root_address_inst_req_0 : boolean;
  signal ptr_deref_1055_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1055_addr_0_req_0 : boolean;
  signal ptr_deref_1055_addr_0_ack_0 : boolean;
  signal ptr_deref_1055_addr_0_req_1 : boolean;
  signal ptr_deref_1055_addr_0_ack_1 : boolean;
  signal ptr_deref_1055_addr_1_req_0 : boolean;
  signal ptr_deref_1055_addr_1_ack_0 : boolean;
  signal ptr_deref_1055_addr_1_req_1 : boolean;
  signal ptr_deref_1055_addr_1_ack_1 : boolean;
  signal ptr_deref_1055_addr_2_req_0 : boolean;
  signal ptr_deref_1055_addr_2_ack_0 : boolean;
  signal ptr_deref_1055_addr_2_req_1 : boolean;
  signal ptr_deref_1055_addr_2_ack_1 : boolean;
  signal ptr_deref_1055_addr_3_req_0 : boolean;
  signal ptr_deref_1055_addr_3_ack_0 : boolean;
  signal ptr_deref_1055_addr_3_req_1 : boolean;
  signal ptr_deref_1055_addr_3_ack_1 : boolean;
  signal ptr_deref_1055_gather_scatter_req_0 : boolean;
  signal ptr_deref_1055_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1055_store_0_req_0 : boolean;
  signal ptr_deref_1055_store_0_ack_0 : boolean;
  signal ptr_deref_1055_store_1_req_0 : boolean;
  signal ptr_deref_1055_store_1_ack_0 : boolean;
  signal ptr_deref_1055_store_2_req_0 : boolean;
  signal ptr_deref_1055_store_2_ack_0 : boolean;
  signal ptr_deref_1055_store_3_req_0 : boolean;
  signal ptr_deref_1055_store_3_ack_0 : boolean;
  signal ptr_deref_1055_store_0_req_1 : boolean;
  signal ptr_deref_1055_store_0_ack_1 : boolean;
  signal ptr_deref_1055_store_1_req_1 : boolean;
  signal ptr_deref_1055_store_1_ack_1 : boolean;
  signal ptr_deref_1055_store_2_req_1 : boolean;
  signal ptr_deref_1055_store_2_ack_1 : boolean;
  signal ptr_deref_1055_store_3_req_1 : boolean;
  signal ptr_deref_1055_store_3_ack_1 : boolean;
  signal array_obj_ref_1063_base_resize_req_0 : boolean;
  signal array_obj_ref_1063_base_resize_ack_0 : boolean;
  signal array_obj_ref_1063_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1063_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1063_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1063_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1063_final_reg_req_0 : boolean;
  signal array_obj_ref_1063_final_reg_ack_0 : boolean;
  signal type_cast_1067_inst_req_0 : boolean;
  signal type_cast_1067_inst_ack_0 : boolean;
  signal ptr_deref_1071_base_resize_req_0 : boolean;
  signal ptr_deref_1071_base_resize_ack_0 : boolean;
  signal ptr_deref_1071_root_address_inst_req_0 : boolean;
  signal ptr_deref_1071_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1071_addr_0_req_0 : boolean;
  signal ptr_deref_1071_addr_0_ack_0 : boolean;
  signal ptr_deref_1071_addr_0_req_1 : boolean;
  signal ptr_deref_1071_addr_0_ack_1 : boolean;
  signal ptr_deref_1071_addr_1_req_0 : boolean;
  signal ptr_deref_1071_addr_1_ack_0 : boolean;
  signal ptr_deref_1071_addr_1_req_1 : boolean;
  signal ptr_deref_1071_addr_1_ack_1 : boolean;
  signal ptr_deref_1071_addr_2_req_0 : boolean;
  signal ptr_deref_1071_addr_2_ack_0 : boolean;
  signal ptr_deref_1071_addr_2_req_1 : boolean;
  signal ptr_deref_1071_addr_2_ack_1 : boolean;
  signal ptr_deref_1071_addr_3_req_0 : boolean;
  signal ptr_deref_1071_addr_3_ack_0 : boolean;
  signal ptr_deref_1071_addr_3_req_1 : boolean;
  signal ptr_deref_1071_addr_3_ack_1 : boolean;
  signal ptr_deref_1071_load_0_req_0 : boolean;
  signal ptr_deref_1071_load_0_ack_0 : boolean;
  signal ptr_deref_1071_load_1_req_0 : boolean;
  signal ptr_deref_1071_load_1_ack_0 : boolean;
  signal ptr_deref_1071_load_2_req_0 : boolean;
  signal ptr_deref_1071_load_2_ack_0 : boolean;
  signal ptr_deref_1071_load_3_req_0 : boolean;
  signal ptr_deref_1071_load_3_ack_0 : boolean;
  signal ptr_deref_1071_load_0_req_1 : boolean;
  signal ptr_deref_1071_load_0_ack_1 : boolean;
  signal ptr_deref_1071_load_1_req_1 : boolean;
  signal ptr_deref_1071_load_1_ack_1 : boolean;
  signal ptr_deref_1071_load_2_req_1 : boolean;
  signal ptr_deref_1071_load_2_ack_1 : boolean;
  signal ptr_deref_1071_load_3_req_1 : boolean;
  signal ptr_deref_1071_load_3_ack_1 : boolean;
  signal ptr_deref_1071_gather_scatter_req_0 : boolean;
  signal ptr_deref_1071_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1078_base_resize_req_0 : boolean;
  signal array_obj_ref_1078_base_resize_ack_0 : boolean;
  signal array_obj_ref_1078_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1078_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1078_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1078_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1078_final_reg_req_0 : boolean;
  signal array_obj_ref_1078_final_reg_ack_0 : boolean;
  signal type_cast_1082_inst_req_0 : boolean;
  signal type_cast_1082_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_chk_CP_1029: Block -- control-path 
    signal cp_elements: BooleanArray(979 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(979);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(979), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(141);
    cpelement_group_2 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(898));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(3) <= cp_elements(213);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(900));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(249) & cp_elements(902));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(287) & cp_elements(904));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(7) <= OrReduce(cp_elements(308) & cp_elements(906));
    cp_elements(8) <= cp_elements(921);
    cp_elements(9) <= cp_elements(391);
    cp_elements(10) <= OrReduce(cp_elements(400) & cp_elements(923));
    cp_elements(11) <= cp_elements(956);
    cp_elements(12) <= OrReduce(cp_elements(430) & cp_elements(958));
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(489) & cp_elements(971));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(14) <= cp_elements(606);
    cp_elements(15) <= OrReduce(cp_elements(613) & cp_elements(973));
    cp_elements(16) <= cp_elements(779);
    cp_elements(17) <= cp_elements(876);
    cp_elements(18) <= OrReduce(cp_elements(975) & cp_elements(977));
    cp_elements(19) <= cp_elements(0);
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(21) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_538_inst_req_0); -- 
    cp_elements(21) <= cp_elements(19);
    cp_elements(22) <= cp_elements(19);
    req_1156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => simple_obj_ref_537_inst_req_0); -- 
    ack_1157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_537_inst_ack_0, ack => cp_elements(23)); -- 
    ack_1162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_538_inst_ack_0, ack => cp_elements(24)); -- 
    cp_elements(25) <= cp_elements(24);
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => type_cast_542_inst_req_0); -- 
    cp_elements(27) <= cp_elements(25);
    cp_elements(28) <= cp_elements(25);
    cp_elements(29) <= type_cast_542_inst_ack_0;
    cp_elements(30) <= cp_elements(25);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1199_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_549_final_reg_req_0); -- 
    cp_elements(32) <= cp_elements(29);
    base_resize_req_1186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_549_base_resize_req_0); -- 
    base_resize_ack_1187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_base_resize_ack_0, ack => cp_elements(33)); -- 
    plus_base_rr_1192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_549_root_address_inst_req_0); -- 
    plus_base_ra_1193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_root_address_inst_ack_0, ack => cp_elements(34)); -- 
    plus_base_cr_1194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_549_root_address_inst_req_1); -- 
    plus_base_ca_1195_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_root_address_inst_ack_1, ack => cp_elements(35)); -- 
    final_reg_ack_1200_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_549_final_reg_ack_0, ack => cp_elements(36)); -- 
    base_resize_req_1213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_553_base_resize_req_0); -- 
    base_resize_ack_1214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_base_resize_ack_0, ack => cp_elements(37)); -- 
    sum_rename_req_1218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_553_root_address_inst_req_0); -- 
    cp_elements(38) <= ptr_deref_553_root_address_inst_ack_0;
    cp_elements(39) <= cp_elements(38);
    rr_1226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => ptr_deref_553_addr_0_req_0); -- 
    ra_1227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_0_ack_0, ack => cp_elements(40)); -- 
    cr_1228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_553_addr_0_req_1); -- 
    ca_1229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_0_ack_1, ack => cp_elements(41)); -- 
    cp_elements(42) <= cp_elements(38);
    rr_1233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_553_addr_1_req_0); -- 
    ra_1234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_1_ack_0, ack => cp_elements(43)); -- 
    cr_1235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_553_addr_1_req_1); -- 
    ca_1236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_1_ack_1, ack => cp_elements(44)); -- 
    cp_elements(45) <= cp_elements(38);
    rr_1240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_553_addr_2_req_0); -- 
    ra_1241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_2_ack_0, ack => cp_elements(46)); -- 
    cr_1242_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_553_addr_2_req_1); -- 
    ca_1243_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_2_ack_1, ack => cp_elements(47)); -- 
    cp_elements(48) <= cp_elements(38);
    rr_1247_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_553_addr_3_req_0); -- 
    ra_1248_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_3_ack_0, ack => cp_elements(49)); -- 
    cr_1249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_553_addr_3_req_1); -- 
    ca_1250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_addr_3_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(41) & cp_elements(44) & cp_elements(47) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(52) <= cp_elements(51);
    rr_1260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_553_load_0_req_0); -- 
    ra_1261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_0_ack_0, ack => cp_elements(53)); -- 
    cp_elements(54) <= cp_elements(51);
    rr_1265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_553_load_1_req_0); -- 
    ra_1266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_1_ack_0, ack => cp_elements(55)); -- 
    cp_elements(56) <= cp_elements(51);
    rr_1270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_553_load_2_req_0); -- 
    ra_1271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_2_ack_0, ack => cp_elements(57)); -- 
    cp_elements(58) <= cp_elements(51);
    rr_1275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_553_load_3_req_0); -- 
    ra_1276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_3_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(55) & cp_elements(57) & cp_elements(59));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(61) <= cp_elements(60);
    cr_1286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_553_load_0_req_1); -- 
    ca_1287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_0_ack_1, ack => cp_elements(62)); -- 
    cp_elements(63) <= cp_elements(60);
    cr_1291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_553_load_1_req_1); -- 
    ca_1292_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_1_ack_1, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(60);
    cr_1296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_553_load_2_req_1); -- 
    ca_1297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_2_ack_1, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(60);
    cr_1301_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_553_load_3_req_1); -- 
    ca_1302_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_553_load_3_ack_1, ack => cp_elements(68)); -- 
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(62) & cp_elements(64) & cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1303_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_553_gather_scatter_req_0); -- 
    cp_elements(70) <= ptr_deref_553_gather_scatter_ack_0;
    cp_elements(71) <= cp_elements(25);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_558_final_reg_req_0); -- 
    cp_elements(73) <= cp_elements(70);
    base_resize_req_1315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_558_base_resize_req_0); -- 
    base_resize_ack_1316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_base_resize_ack_0, ack => cp_elements(74)); -- 
    plus_base_rr_1321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_558_root_address_inst_req_0); -- 
    plus_base_ra_1322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_root_address_inst_ack_0, ack => cp_elements(75)); -- 
    plus_base_cr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_558_root_address_inst_req_1); -- 
    plus_base_ca_1324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_root_address_inst_ack_1, ack => cp_elements(76)); -- 
    final_reg_ack_1329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_558_final_reg_ack_0, ack => cp_elements(77)); -- 
    cp_elements(78) <= cp_elements(25);
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(83));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_1353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => array_obj_ref_565_final_reg_req_0); -- 
    cp_elements(80) <= cp_elements(29);
    base_resize_req_1340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => array_obj_ref_565_base_resize_req_0); -- 
    base_resize_ack_1341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_base_resize_ack_0, ack => cp_elements(81)); -- 
    plus_base_rr_1346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_565_root_address_inst_req_0); -- 
    plus_base_ra_1347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_root_address_inst_ack_0, ack => cp_elements(82)); -- 
    plus_base_cr_1348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_565_root_address_inst_req_1); -- 
    plus_base_ca_1349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_root_address_inst_ack_1, ack => cp_elements(83)); -- 
    final_reg_ack_1354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_565_final_reg_ack_0, ack => cp_elements(84)); -- 
    base_resize_req_1367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_569_base_resize_req_0); -- 
    base_resize_ack_1368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_base_resize_ack_0, ack => cp_elements(85)); -- 
    sum_rename_req_1372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_569_root_address_inst_req_0); -- 
    cp_elements(86) <= ptr_deref_569_root_address_inst_ack_0;
    cp_elements(87) <= cp_elements(86);
    rr_1380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => ptr_deref_569_addr_0_req_0); -- 
    ra_1381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_0_ack_0, ack => cp_elements(88)); -- 
    cr_1382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_569_addr_0_req_1); -- 
    ca_1383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_0_ack_1, ack => cp_elements(89)); -- 
    cp_elements(90) <= cp_elements(86);
    rr_1387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => ptr_deref_569_addr_1_req_0); -- 
    ra_1388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_1_ack_0, ack => cp_elements(91)); -- 
    cr_1389_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => ptr_deref_569_addr_1_req_1); -- 
    ca_1390_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_1_ack_1, ack => cp_elements(92)); -- 
    cp_elements(93) <= cp_elements(86);
    rr_1394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_569_addr_2_req_0); -- 
    ra_1395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_2_ack_0, ack => cp_elements(94)); -- 
    cr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_569_addr_2_req_1); -- 
    ca_1397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_2_ack_1, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(86);
    rr_1401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_569_addr_3_req_0); -- 
    ra_1402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_3_ack_0, ack => cp_elements(97)); -- 
    cr_1403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_569_addr_3_req_1); -- 
    ca_1404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_addr_3_ack_1, ack => cp_elements(98)); -- 
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(92) & cp_elements(95) & cp_elements(98));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(100) <= cp_elements(99);
    rr_1414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_569_load_0_req_0); -- 
    ra_1415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_0_ack_0, ack => cp_elements(101)); -- 
    cp_elements(102) <= cp_elements(99);
    rr_1419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => ptr_deref_569_load_1_req_0); -- 
    ra_1420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_1_ack_0, ack => cp_elements(103)); -- 
    cp_elements(104) <= cp_elements(99);
    rr_1424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_569_load_2_req_0); -- 
    ra_1425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_2_ack_0, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(99);
    rr_1429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_569_load_3_req_0); -- 
    ra_1430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_3_ack_0, ack => cp_elements(107)); -- 
    cpelement_group_108 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(101) & cp_elements(103) & cp_elements(105) & cp_elements(107));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(108),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(109) <= cp_elements(108);
    cr_1440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_569_load_0_req_1); -- 
    ca_1441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_0_ack_1, ack => cp_elements(110)); -- 
    cp_elements(111) <= cp_elements(108);
    cr_1445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_569_load_1_req_1); -- 
    ca_1446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_1_ack_1, ack => cp_elements(112)); -- 
    cp_elements(113) <= cp_elements(108);
    cr_1450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_569_load_2_req_1); -- 
    ca_1451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_2_ack_1, ack => cp_elements(114)); -- 
    cp_elements(115) <= cp_elements(108);
    cr_1455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_569_load_3_req_1); -- 
    ca_1456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_load_3_ack_1, ack => cp_elements(116)); -- 
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112) & cp_elements(114) & cp_elements(116));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_569_gather_scatter_req_0); -- 
    merge_ack_1458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_569_gather_scatter_ack_0, ack => cp_elements(118)); -- 
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(120));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => type_cast_573_inst_req_0); -- 
    cp_elements(120) <= cp_elements(25);
    ack_1468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_573_inst_ack_0, ack => cp_elements(121)); -- 
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(124));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => type_cast_577_inst_req_0); -- 
    cp_elements(123) <= cp_elements(25);
    cp_elements(124) <= cp_elements(70);
    ack_1478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_577_inst_ack_0, ack => cp_elements(125)); -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(121) & cp_elements(125) & cp_elements(127));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => binary_582_inst_req_0); -- 
    cp_elements(127) <= cp_elements(25);
    ra_1489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_582_inst_ack_0, ack => cp_elements(128)); -- 
    cr_1490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => binary_582_inst_req_1); -- 
    ca_1491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_582_inst_ack_1, ack => cp_elements(129)); -- 
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(129) & cp_elements(131));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => binary_588_inst_req_0); -- 
    cp_elements(131) <= cp_elements(25);
    ra_1501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_0, ack => cp_elements(132)); -- 
    cr_1502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => binary_588_inst_req_1); -- 
    ca_1503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_588_inst_ack_1, ack => cp_elements(133)); -- 
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(135) & cp_elements(138));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => binary_597_inst_req_0); -- 
    cp_elements(135) <= cp_elements(25);
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => type_cast_593_inst_req_0); -- 
    cp_elements(137) <= cp_elements(25);
    ack_1515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_593_inst_ack_0, ack => cp_elements(138)); -- 
    ra_1520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_597_inst_ack_0, ack => cp_elements(139)); -- 
    cr_1521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => binary_597_inst_req_1); -- 
    ca_1522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_597_inst_ack_1, ack => cp_elements(140)); -- 
    cpelement_group_141 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(77) & cp_elements(140));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(141),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(142) <= cp_elements(1);
    cp_elements(143) <= false;
    cp_elements(144) <= cp_elements(143);
    cp_elements(145) <= cp_elements(1);
    branch_req_1530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => if_stmt_599_branch_req_0); -- 
    cp_elements(146) <= cp_elements(145);
    cp_elements(147) <= cp_elements(146);
    if_choice_transition_1535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_599_branch_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    else_choice_transition_1539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_599_branch_ack_0, ack => cp_elements(150)); -- 
    cpelement_group_151 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(152) & cp_elements(153));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(151),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => binary_610_inst_req_0); -- 
    cp_elements(152) <= cp_elements(2);
    cp_elements(153) <= cp_elements(2);
    ra_1557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_610_inst_ack_0, ack => cp_elements(154)); -- 
    cr_1558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => binary_610_inst_req_1); -- 
    ca_1559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_610_inst_ack_1, ack => cp_elements(155)); -- 
    pipe_wreq_1564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => simple_obj_ref_607_inst_req_0); -- 
    pipe_wack_1565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_607_inst_ack_0, ack => cp_elements(156)); -- 
    cp_elements(157) <= cp_elements(150);
    cpelement_group_158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(159) & cp_elements(160));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => type_cast_617_inst_req_0); -- 
    cp_elements(159) <= cp_elements(157);
    cp_elements(160) <= cp_elements(157);
    ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_617_inst_ack_0, ack => cp_elements(161)); -- 
    base_resize_req_1591_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => ptr_deref_621_base_resize_req_0); -- 
    base_resize_ack_1592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_base_resize_ack_0, ack => cp_elements(162)); -- 
    sum_rename_req_1596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => ptr_deref_621_root_address_inst_req_0); -- 
    cp_elements(163) <= ptr_deref_621_root_address_inst_ack_0;
    cp_elements(164) <= cp_elements(163);
    rr_1604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => ptr_deref_621_addr_0_req_0); -- 
    ra_1605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_0_ack_0, ack => cp_elements(165)); -- 
    cr_1606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => ptr_deref_621_addr_0_req_1); -- 
    ca_1607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_0_ack_1, ack => cp_elements(166)); -- 
    cp_elements(167) <= cp_elements(163);
    rr_1611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => ptr_deref_621_addr_1_req_0); -- 
    ra_1612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_1_ack_0, ack => cp_elements(168)); -- 
    cr_1613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => ptr_deref_621_addr_1_req_1); -- 
    ca_1614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_1_ack_1, ack => cp_elements(169)); -- 
    cp_elements(170) <= cp_elements(163);
    rr_1618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => ptr_deref_621_addr_2_req_0); -- 
    ra_1619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_2_ack_0, ack => cp_elements(171)); -- 
    cr_1620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => ptr_deref_621_addr_2_req_1); -- 
    ca_1621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_2_ack_1, ack => cp_elements(172)); -- 
    cp_elements(173) <= cp_elements(163);
    rr_1625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => ptr_deref_621_addr_3_req_0); -- 
    ra_1626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_3_ack_0, ack => cp_elements(174)); -- 
    cr_1627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(174), ack => ptr_deref_621_addr_3_req_1); -- 
    ca_1628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_addr_3_ack_1, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(166) & cp_elements(169) & cp_elements(172) & cp_elements(175));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(177) <= cp_elements(176);
    rr_1638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => ptr_deref_621_load_0_req_0); -- 
    ra_1639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_0_ack_0, ack => cp_elements(178)); -- 
    cp_elements(179) <= cp_elements(176);
    rr_1643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => ptr_deref_621_load_1_req_0); -- 
    ra_1644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_1_ack_0, ack => cp_elements(180)); -- 
    cp_elements(181) <= cp_elements(176);
    rr_1648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => ptr_deref_621_load_2_req_0); -- 
    ra_1649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_2_ack_0, ack => cp_elements(182)); -- 
    cp_elements(183) <= cp_elements(176);
    rr_1653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => ptr_deref_621_load_3_req_0); -- 
    ra_1654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_3_ack_0, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(180) & cp_elements(182) & cp_elements(184));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(186) <= cp_elements(185);
    cr_1664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => ptr_deref_621_load_0_req_1); -- 
    ca_1665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_0_ack_1, ack => cp_elements(187)); -- 
    cp_elements(188) <= cp_elements(185);
    cr_1669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_621_load_1_req_1); -- 
    ca_1670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_1_ack_1, ack => cp_elements(189)); -- 
    cp_elements(190) <= cp_elements(185);
    cr_1674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_621_load_2_req_1); -- 
    ca_1675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_2_ack_1, ack => cp_elements(191)); -- 
    cp_elements(192) <= cp_elements(185);
    cr_1679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_621_load_3_req_1); -- 
    ca_1680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_621_load_3_ack_1, ack => cp_elements(193)); -- 
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(187) & cp_elements(189) & cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_1681_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => ptr_deref_621_gather_scatter_req_0); -- 
    cp_elements(195) <= ptr_deref_621_gather_scatter_ack_0;
    cpelement_group_196 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(197) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => binary_627_inst_req_0); -- 
    cp_elements(197) <= cp_elements(157);
    cp_elements(198) <= cp_elements(195);
    ra_1692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_627_inst_ack_0, ack => cp_elements(199)); -- 
    cr_1693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => binary_627_inst_req_1); -- 
    ca_1694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_627_inst_ack_1, ack => cp_elements(200)); -- 
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(202));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => binary_633_inst_req_0); -- 
    cp_elements(202) <= cp_elements(157);
    ra_1704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_633_inst_ack_0, ack => cp_elements(203)); -- 
    cr_1705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => binary_633_inst_req_1); -- 
    ca_1706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_633_inst_ack_1, ack => cp_elements(204)); -- 
    cpelement_group_205 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(206) & cp_elements(207));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(205),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1715_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => binary_639_inst_req_0); -- 
    cp_elements(206) <= cp_elements(157);
    cp_elements(207) <= cp_elements(195);
    ra_1716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_639_inst_ack_0, ack => cp_elements(208)); -- 
    cr_1717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => binary_639_inst_req_1); -- 
    ca_1718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_639_inst_ack_1, ack => cp_elements(209)); -- 
    cpelement_group_210 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(209) & cp_elements(211));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(210),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => type_cast_643_inst_req_0); -- 
    cp_elements(211) <= cp_elements(157);
    ack_1728_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_643_inst_ack_0, ack => cp_elements(212)); -- 
    cpelement_group_213 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(204) & cp_elements(212));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(213),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(214) <= cp_elements(3);
    cp_elements(215) <= false;
    cp_elements(216) <= cp_elements(215);
    cp_elements(217) <= cp_elements(3);
    branch_req_1736_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => if_stmt_645_branch_req_0); -- 
    cp_elements(218) <= cp_elements(217);
    cp_elements(219) <= cp_elements(218);
    if_choice_transition_1741_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_645_branch_ack_1, ack => cp_elements(220)); -- 
    cp_elements(221) <= cp_elements(218);
    else_choice_transition_1745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_645_branch_ack_0, ack => cp_elements(222)); -- 
    cpelement_group_223 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(224) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(223),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => binary_656_inst_req_0); -- 
    cp_elements(224) <= cp_elements(4);
    cp_elements(225) <= cp_elements(4);
    ra_1763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_656_inst_ack_0, ack => cp_elements(226)); -- 
    cr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => binary_656_inst_req_1); -- 
    ca_1765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_656_inst_ack_1, ack => cp_elements(227)); -- 
    pipe_wreq_1770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => simple_obj_ref_653_inst_req_0); -- 
    pipe_wack_1771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_653_inst_ack_0, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(220);
    cpelement_group_230 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(231) & cp_elements(232));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(230),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => binary_665_inst_req_0); -- 
    cp_elements(231) <= cp_elements(229);
    cp_elements(232) <= cp_elements(229);
    ra_1784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_665_inst_ack_0, ack => cp_elements(233)); -- 
    cr_1785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => binary_665_inst_req_1); -- 
    ca_1786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_665_inst_ack_1, ack => cp_elements(234)); -- 
    cpelement_group_235 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(234) & cp_elements(236));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(235),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => binary_671_inst_req_0); -- 
    cp_elements(236) <= cp_elements(229);
    ra_1796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_671_inst_ack_0, ack => cp_elements(237)); -- 
    cr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => binary_671_inst_req_1); -- 
    ca_1798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_671_inst_ack_1, ack => cp_elements(238)); -- 
    cpelement_group_239 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(240));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(239),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => binary_677_inst_req_0); -- 
    cp_elements(240) <= cp_elements(229);
    ra_1808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_677_inst_ack_0, ack => cp_elements(241)); -- 
    cr_1809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => binary_677_inst_req_1); -- 
    ca_1810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_677_inst_ack_1, ack => cp_elements(242)); -- 
    cp_elements(243) <= cp_elements(242);
    cp_elements(244) <= false;
    cp_elements(245) <= cp_elements(244);
    cp_elements(246) <= cp_elements(242);
    branch_req_1818_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => if_stmt_679_branch_req_0); -- 
    cp_elements(247) <= cp_elements(246);
    cp_elements(248) <= cp_elements(247);
    if_choice_transition_1823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_679_branch_ack_1, ack => cp_elements(249)); -- 
    cp_elements(250) <= cp_elements(247);
    else_choice_transition_1827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_679_branch_ack_0, ack => cp_elements(251)); -- 
    crr_1863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => call_stmt_697_call_req_0); -- 
    cpelement_group_252 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(253) & cp_elements(254));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(252),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => binary_690_inst_req_0); -- 
    cp_elements(253) <= cp_elements(5);
    cp_elements(254) <= cp_elements(5);
    ra_1845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_690_inst_ack_0, ack => cp_elements(255)); -- 
    cr_1846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => binary_690_inst_req_1); -- 
    ca_1847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_690_inst_ack_1, ack => cp_elements(256)); -- 
    pipe_wreq_1852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => simple_obj_ref_687_inst_req_0); -- 
    pipe_wack_1853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_687_inst_ack_0, ack => cp_elements(257)); -- 
    cra_1864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_697_call_ack_0, ack => cp_elements(258)); -- 
    ccr_1868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => call_stmt_697_call_req_1); -- 
    cca_1869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_697_call_ack_1, ack => cp_elements(259)); -- 
    cp_elements(260) <= cp_elements(259);
    cpelement_group_261 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(263));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(261),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_1883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => type_cast_700_inst_req_0); -- 
    cp_elements(262) <= cp_elements(260);
    cp_elements(263) <= cp_elements(260);
    cp_elements(264) <= type_cast_700_inst_ack_0;
    cpelement_group_265 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(266) & cp_elements(267) & cp_elements(268));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(265),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => binary_705_inst_req_0); -- 
    cp_elements(266) <= cp_elements(260);
    cp_elements(267) <= cp_elements(264);
    cp_elements(268) <= cp_elements(260);
    ra_1895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_705_inst_ack_0, ack => cp_elements(269)); -- 
    cr_1896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => binary_705_inst_req_1); -- 
    ca_1897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_705_inst_ack_1, ack => cp_elements(270)); -- 
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(272) & cp_elements(273) & cp_elements(274));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => binary_710_inst_req_0); -- 
    cp_elements(272) <= cp_elements(260);
    cp_elements(273) <= cp_elements(264);
    cp_elements(274) <= cp_elements(260);
    ra_1908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_710_inst_ack_0, ack => cp_elements(275)); -- 
    cr_1909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => binary_710_inst_req_1); -- 
    ca_1910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_710_inst_ack_1, ack => cp_elements(276)); -- 
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(270) & cp_elements(276) & cp_elements(278));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => binary_715_inst_req_0); -- 
    cp_elements(278) <= cp_elements(260);
    ra_1921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_715_inst_ack_0, ack => cp_elements(279)); -- 
    cr_1922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => binary_715_inst_req_1); -- 
    ca_1923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_715_inst_ack_1, ack => cp_elements(280)); -- 
    cp_elements(281) <= cp_elements(280);
    cp_elements(282) <= false;
    cp_elements(283) <= cp_elements(282);
    cp_elements(284) <= cp_elements(280);
    branch_req_1931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => if_stmt_717_branch_req_0); -- 
    cp_elements(285) <= cp_elements(284);
    cp_elements(286) <= cp_elements(285);
    if_choice_transition_1936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(285);
    else_choice_transition_1940_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_0, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(292));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => binary_728_inst_req_0); -- 
    cp_elements(291) <= cp_elements(6);
    cp_elements(292) <= cp_elements(6);
    ra_1958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_728_inst_ack_0, ack => cp_elements(293)); -- 
    cr_1959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => binary_728_inst_req_1); -- 
    ca_1960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_728_inst_ack_1, ack => cp_elements(294)); -- 
    pipe_wreq_1965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => simple_obj_ref_725_inst_req_0); -- 
    pipe_wack_1966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_725_inst_ack_0, ack => cp_elements(295)); -- 
    cp_elements(296) <= cp_elements(289);
    cpelement_group_297 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(298) & cp_elements(299));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(297),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_1978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => binary_737_inst_req_0); -- 
    cp_elements(298) <= cp_elements(296);
    cp_elements(299) <= cp_elements(296);
    ra_1979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_737_inst_ack_0, ack => cp_elements(300)); -- 
    cr_1980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => binary_737_inst_req_1); -- 
    ca_1981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_737_inst_ack_1, ack => cp_elements(301)); -- 
    cp_elements(302) <= cp_elements(301);
    cp_elements(303) <= false;
    cp_elements(304) <= cp_elements(303);
    cp_elements(305) <= cp_elements(301);
    branch_req_1989_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => if_stmt_739_branch_req_0); -- 
    cp_elements(306) <= cp_elements(305);
    cp_elements(307) <= cp_elements(306);
    if_choice_transition_1994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_739_branch_ack_1, ack => cp_elements(308)); -- 
    cp_elements(309) <= cp_elements(306);
    else_choice_transition_1998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_739_branch_ack_0, ack => cp_elements(310)); -- 
    cp_elements(311) <= cp_elements(7);
    cpelement_group_312 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(314));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(312),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => binary_750_inst_req_0); -- 
    cp_elements(313) <= cp_elements(311);
    cp_elements(314) <= cp_elements(311);
    ra_2013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_750_inst_ack_0, ack => cp_elements(315)); -- 
    cr_2014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => binary_750_inst_req_1); -- 
    ca_2015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_750_inst_ack_1, ack => cp_elements(316)); -- 
    cp_elements(317) <= cp_elements(8);
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(320));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => binary_773_inst_req_0); -- 
    cp_elements(319) <= cp_elements(317);
    cp_elements(320) <= cp_elements(317);
    ra_2028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_773_inst_ack_0, ack => cp_elements(321)); -- 
    cr_2029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => binary_773_inst_req_1); -- 
    ca_2030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_773_inst_ack_1, ack => cp_elements(322)); -- 
    cpelement_group_323 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(322) & cp_elements(324) & cp_elements(325));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(323),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => binary_778_inst_req_0); -- 
    cp_elements(324) <= cp_elements(317);
    cp_elements(325) <= cp_elements(317);
    ra_2041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_778_inst_ack_0, ack => cp_elements(326)); -- 
    cr_2042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => binary_778_inst_req_1); -- 
    ca_2043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_778_inst_ack_1, ack => cp_elements(327)); -- 
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(330));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2052_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => binary_784_inst_req_0); -- 
    cp_elements(329) <= cp_elements(317);
    cp_elements(330) <= cp_elements(317);
    ra_2053_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_784_inst_ack_0, ack => cp_elements(331)); -- 
    cr_2054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => binary_784_inst_req_1); -- 
    ca_2055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_784_inst_ack_1, ack => cp_elements(332)); -- 
    cpelement_group_333 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(332) & cp_elements(334));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(333),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => binary_790_inst_req_0); -- 
    cp_elements(334) <= cp_elements(317);
    ra_2065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_790_inst_ack_0, ack => cp_elements(335)); -- 
    cr_2066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => binary_790_inst_req_1); -- 
    ca_2067_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_790_inst_ack_1, ack => cp_elements(336)); -- 
    index_resize_req_2082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => array_obj_ref_794_index_0_resize_req_0); -- 
    cp_elements(337) <= cp_elements(317);
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(337) & cp_elements(346));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => array_obj_ref_794_final_reg_req_0); -- 
    cp_elements(339) <= cp_elements(317);
    base_resize_req_2098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => array_obj_ref_794_base_resize_req_0); -- 
    index_resize_ack_2083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_index_0_resize_ack_0, ack => cp_elements(340)); -- 
    scale_rename_req_2087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => array_obj_ref_794_index_0_rename_req_0); -- 
    scale_rename_ack_2088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_index_0_rename_ack_0, ack => cp_elements(341)); -- 
    final_index_req_2092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => array_obj_ref_794_offset_inst_req_0); -- 
    final_index_ack_2093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_offset_inst_ack_0, ack => cp_elements(342)); -- 
    base_resize_ack_2099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_base_resize_ack_0, ack => cp_elements(343)); -- 
    cpelement_group_344 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(342) & cp_elements(343));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(344), ack => array_obj_ref_794_root_address_inst_req_0); -- 
    plus_base_ra_2105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_root_address_inst_ack_0, ack => cp_elements(345)); -- 
    plus_base_cr_2106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => array_obj_ref_794_root_address_inst_req_1); -- 
    plus_base_ca_2107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_root_address_inst_ack_1, ack => cp_elements(346)); -- 
    final_reg_ack_2112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_794_final_reg_ack_0, ack => cp_elements(347)); -- 
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => type_cast_799_inst_req_0); -- 
    cp_elements(349) <= cp_elements(317);
    ack_2122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_799_inst_ack_0, ack => cp_elements(350)); -- 
    base_resize_req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => ptr_deref_803_base_resize_req_0); -- 
    base_resize_ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_base_resize_ack_0, ack => cp_elements(351)); -- 
    sum_rename_req_2140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => ptr_deref_803_root_address_inst_req_0); -- 
    cp_elements(352) <= ptr_deref_803_root_address_inst_ack_0;
    cp_elements(353) <= cp_elements(352);
    rr_2148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => ptr_deref_803_addr_0_req_0); -- 
    ra_2149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_addr_0_ack_0, ack => cp_elements(354)); -- 
    cr_2150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(354), ack => ptr_deref_803_addr_0_req_1); -- 
    ca_2151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_addr_0_ack_1, ack => cp_elements(355)); -- 
    cp_elements(356) <= cp_elements(352);
    rr_2155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => ptr_deref_803_addr_1_req_0); -- 
    ra_2156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_addr_1_ack_0, ack => cp_elements(357)); -- 
    cr_2157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => ptr_deref_803_addr_1_req_1); -- 
    ca_2158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_addr_1_ack_1, ack => cp_elements(358)); -- 
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(355) & cp_elements(358));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(360) <= cp_elements(359);
    rr_2168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => ptr_deref_803_load_0_req_0); -- 
    ra_2169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_0_ack_0, ack => cp_elements(361)); -- 
    cp_elements(362) <= cp_elements(359);
    rr_2173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => ptr_deref_803_load_1_req_0); -- 
    ra_2174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_1_ack_0, ack => cp_elements(363)); -- 
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(363));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(365) <= cp_elements(364);
    cr_2184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(365), ack => ptr_deref_803_load_0_req_1); -- 
    ca_2185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_0_ack_1, ack => cp_elements(366)); -- 
    cp_elements(367) <= cp_elements(364);
    cr_2189_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(367), ack => ptr_deref_803_load_1_req_1); -- 
    ca_2190_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_load_1_ack_1, ack => cp_elements(368)); -- 
    cpelement_group_369 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(366) & cp_elements(368));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(369),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_2191_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(369), ack => ptr_deref_803_gather_scatter_req_0); -- 
    merge_ack_2192_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_803_gather_scatter_ack_0, ack => cp_elements(370)); -- 
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(370) & cp_elements(372));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => type_cast_807_inst_req_0); -- 
    cp_elements(372) <= cp_elements(317);
    ack_2202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_807_inst_ack_0, ack => cp_elements(373)); -- 
    cpelement_group_374 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(373) & cp_elements(375) & cp_elements(376));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2212_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(374), ack => binary_812_inst_req_0); -- 
    cp_elements(375) <= cp_elements(317);
    cp_elements(376) <= cp_elements(317);
    ra_2213_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_812_inst_ack_0, ack => cp_elements(377)); -- 
    cr_2214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(377), ack => binary_812_inst_req_1); -- 
    ca_2215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_812_inst_ack_1, ack => cp_elements(378)); -- 
    cpelement_group_379 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(380) & cp_elements(383));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(379),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => binary_820_inst_req_0); -- 
    cp_elements(380) <= cp_elements(317);
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(327) & cp_elements(382));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2226_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => type_cast_816_inst_req_0); -- 
    cp_elements(382) <= cp_elements(317);
    ack_2227_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_816_inst_ack_0, ack => cp_elements(383)); -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_820_inst_ack_0, ack => cp_elements(384)); -- 
    cr_2233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => binary_820_inst_req_1); -- 
    ca_2234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_820_inst_ack_1, ack => cp_elements(385)); -- 
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(387) & cp_elements(388));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => binary_826_inst_req_0); -- 
    cp_elements(387) <= cp_elements(317);
    cp_elements(388) <= cp_elements(317);
    ra_2244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_826_inst_ack_0, ack => cp_elements(389)); -- 
    cr_2245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(389), ack => binary_826_inst_req_1); -- 
    ca_2246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_826_inst_ack_1, ack => cp_elements(390)); -- 
    cpelement_group_391 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(378) & cp_elements(385) & cp_elements(390));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(391),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(392) <= cp_elements(9);
    cp_elements(393) <= false;
    cp_elements(394) <= cp_elements(393);
    cp_elements(395) <= cp_elements(9);
    branch_req_2254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(395), ack => if_stmt_828_branch_req_0); -- 
    cp_elements(396) <= cp_elements(395);
    cp_elements(397) <= cp_elements(396);
    if_choice_transition_2259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_828_branch_ack_1, ack => cp_elements(398)); -- 
    cp_elements(399) <= cp_elements(396);
    else_choice_transition_2263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_828_branch_ack_0, ack => cp_elements(400)); -- 
    cp_elements(401) <= cp_elements(10);
    cpelement_group_402 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(403) & cp_elements(404));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(402),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => binary_839_inst_req_0); -- 
    cp_elements(403) <= cp_elements(401);
    cp_elements(404) <= cp_elements(401);
    ra_2278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_839_inst_ack_0, ack => cp_elements(405)); -- 
    cr_2279_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(405), ack => binary_839_inst_req_1); -- 
    ca_2280_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_839_inst_ack_1, ack => cp_elements(406)); -- 
    index_resize_req_2295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => array_obj_ref_843_index_0_resize_req_0); -- 
    cp_elements(407) <= cp_elements(401);
    cpelement_group_408 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(407) & cp_elements(416));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(408),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(408), ack => array_obj_ref_843_final_reg_req_0); -- 
    cp_elements(409) <= cp_elements(401);
    base_resize_req_2311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(409), ack => array_obj_ref_843_base_resize_req_0); -- 
    index_resize_ack_2296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_index_0_resize_ack_0, ack => cp_elements(410)); -- 
    scale_rename_req_2300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(410), ack => array_obj_ref_843_index_0_rename_req_0); -- 
    scale_rename_ack_2301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_index_0_rename_ack_0, ack => cp_elements(411)); -- 
    final_index_req_2305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => array_obj_ref_843_offset_inst_req_0); -- 
    final_index_ack_2306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_offset_inst_ack_0, ack => cp_elements(412)); -- 
    base_resize_ack_2312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_base_resize_ack_0, ack => cp_elements(413)); -- 
    cpelement_group_414 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(412) & cp_elements(413));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(414),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => array_obj_ref_843_root_address_inst_req_0); -- 
    plus_base_ra_2318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_root_address_inst_ack_0, ack => cp_elements(415)); -- 
    plus_base_cr_2319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(415), ack => array_obj_ref_843_root_address_inst_req_1); -- 
    plus_base_ca_2320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_root_address_inst_ack_1, ack => cp_elements(416)); -- 
    final_reg_ack_2325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_843_final_reg_ack_0, ack => cp_elements(417)); -- 
    cp_elements(418) <= cp_elements(11);
    cpelement_group_419 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(420) & cp_elements(421));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(419),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2337_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(419), ack => binary_871_inst_req_0); -- 
    cp_elements(420) <= cp_elements(418);
    cp_elements(421) <= cp_elements(418);
    ra_2338_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_871_inst_ack_0, ack => cp_elements(422)); -- 
    cr_2339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(422), ack => binary_871_inst_req_1); -- 
    ca_2340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_871_inst_ack_1, ack => cp_elements(423)); -- 
    cp_elements(424) <= cp_elements(423);
    cp_elements(425) <= false;
    cp_elements(426) <= cp_elements(425);
    cp_elements(427) <= cp_elements(423);
    branch_req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(427), ack => if_stmt_873_branch_req_0); -- 
    cp_elements(428) <= cp_elements(427);
    cp_elements(429) <= cp_elements(428);
    if_choice_transition_2353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_873_branch_ack_1, ack => cp_elements(430)); -- 
    cp_elements(431) <= cp_elements(428);
    cp_elements(432) <= if_stmt_873_branch_ack_0;
    cp_elements(433) <= cp_elements(12);
    cp_elements(434) <= cp_elements(433);
    base_resize_req_2375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(434), ack => ptr_deref_882_base_resize_req_0); -- 
    base_resize_ack_2376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_base_resize_ack_0, ack => cp_elements(435)); -- 
    sum_rename_req_2380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => ptr_deref_882_root_address_inst_req_0); -- 
    sum_rename_ack_2381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_root_address_inst_ack_0, ack => cp_elements(436)); -- 
    root_rename_req_2385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => ptr_deref_882_addr_0_req_0); -- 
    root_rename_ack_2386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_addr_0_ack_0, ack => cp_elements(437)); -- 
    rr_2396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(437), ack => ptr_deref_882_load_0_req_0); -- 
    ra_2397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_load_0_ack_0, ack => cp_elements(438)); -- 
    cr_2407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => ptr_deref_882_load_0_req_1); -- 
    ca_2408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_load_0_ack_1, ack => cp_elements(439)); -- 
    merge_req_2409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(439), ack => ptr_deref_882_gather_scatter_req_0); -- 
    merge_ack_2410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_882_gather_scatter_ack_0, ack => cp_elements(440)); -- 
    cpelement_group_441 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(440) & cp_elements(442));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(441),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => type_cast_886_inst_req_0); -- 
    cp_elements(442) <= cp_elements(433);
    ack_2420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_886_inst_ack_0, ack => cp_elements(443)); -- 
    cpelement_group_444 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(443) & cp_elements(445) & cp_elements(446));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(444),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => binary_891_inst_req_0); -- 
    cp_elements(445) <= cp_elements(433);
    cp_elements(446) <= cp_elements(433);
    ra_2431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_891_inst_ack_0, ack => cp_elements(447)); -- 
    cr_2432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(447), ack => binary_891_inst_req_1); -- 
    cp_elements(448) <= binary_891_inst_ack_1;
    cp_elements(449) <= cp_elements(969);
    cpelement_group_450 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(452));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(450),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(450), ack => binary_906_inst_req_0); -- 
    cp_elements(451) <= cp_elements(449);
    cp_elements(452) <= cp_elements(449);
    ra_2446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_906_inst_ack_0, ack => cp_elements(453)); -- 
    cr_2447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(453), ack => binary_906_inst_req_1); -- 
    ca_2448_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_906_inst_ack_1, ack => cp_elements(454)); -- 
    cpelement_group_455 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(456) & cp_elements(457));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(455),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => binary_912_inst_req_0); -- 
    cp_elements(456) <= cp_elements(449);
    cp_elements(457) <= cp_elements(449);
    ra_2458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_912_inst_ack_0, ack => cp_elements(458)); -- 
    cr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => binary_912_inst_req_1); -- 
    ca_2460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_912_inst_ack_1, ack => cp_elements(459)); -- 
    cpelement_group_460 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(454) & cp_elements(459) & cp_elements(461));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(460),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => binary_917_inst_req_0); -- 
    cp_elements(461) <= cp_elements(449);
    ra_2471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_917_inst_ack_0, ack => cp_elements(462)); -- 
    cr_2472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => binary_917_inst_req_1); -- 
    cp_elements(463) <= binary_917_inst_ack_1;
    cpelement_group_464 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(465) & cp_elements(466));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(464),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(464), ack => binary_923_inst_req_0); -- 
    cp_elements(465) <= cp_elements(449);
    cp_elements(466) <= cp_elements(463);
    ra_2483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_923_inst_ack_0, ack => cp_elements(467)); -- 
    cr_2484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => binary_923_inst_req_1); -- 
    ca_2485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_923_inst_ack_1, ack => cp_elements(468)); -- 
    cpelement_group_469 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(470) & cp_elements(471));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(469),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => binary_928_inst_req_0); -- 
    cp_elements(470) <= cp_elements(449);
    cp_elements(471) <= cp_elements(463);
    ra_2496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_928_inst_ack_0, ack => cp_elements(472)); -- 
    cr_2497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(472), ack => binary_928_inst_req_1); -- 
    ca_2498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_928_inst_ack_1, ack => cp_elements(473)); -- 
    cpelement_group_474 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(473) & cp_elements(475));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(474),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(474), ack => type_cast_932_inst_req_0); -- 
    cp_elements(475) <= cp_elements(449);
    ack_2508_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_932_inst_ack_0, ack => cp_elements(476)); -- 
    cpelement_group_477 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(476) & cp_elements(478));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(477),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => binary_938_inst_req_0); -- 
    cp_elements(478) <= cp_elements(449);
    ra_2518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_938_inst_ack_0, ack => cp_elements(479)); -- 
    cr_2519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(479), ack => binary_938_inst_req_1); -- 
    ca_2520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_938_inst_ack_1, ack => cp_elements(480)); -- 
    cp_elements(481) <= cp_elements(480);
    cp_elements(482) <= false;
    cp_elements(483) <= cp_elements(482);
    cp_elements(484) <= cp_elements(480);
    branch_req_2528_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => if_stmt_940_branch_req_0); -- 
    cp_elements(485) <= cp_elements(484);
    cp_elements(486) <= cp_elements(485);
    if_choice_transition_2533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_940_branch_ack_1, ack => cp_elements(487)); -- 
    cp_elements(488) <= cp_elements(485);
    else_choice_transition_2537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_940_branch_ack_0, ack => cp_elements(489)); -- 
    cpelement_group_490 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(491) & cp_elements(492));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(490),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => binary_951_inst_req_0); -- 
    cp_elements(491) <= cp_elements(13);
    cp_elements(492) <= cp_elements(13);
    ra_2555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_951_inst_ack_0, ack => cp_elements(493)); -- 
    cr_2556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(493), ack => binary_951_inst_req_1); -- 
    ca_2557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_951_inst_ack_1, ack => cp_elements(494)); -- 
    pipe_wreq_2562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(494), ack => simple_obj_ref_948_inst_req_0); -- 
    pipe_wack_2563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_948_inst_ack_0, ack => cp_elements(495)); -- 
    cp_elements(496) <= cp_elements(487);
    cp_elements(497) <= cp_elements(496);
    cpelement_group_498 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(497) & cp_elements(502));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(498),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(498), ack => array_obj_ref_961_final_reg_req_0); -- 
    cp_elements(499) <= cp_elements(496);
    base_resize_req_2577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => array_obj_ref_961_base_resize_req_0); -- 
    base_resize_ack_2578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_961_base_resize_ack_0, ack => cp_elements(500)); -- 
    plus_base_rr_2583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => array_obj_ref_961_root_address_inst_req_0); -- 
    plus_base_ra_2584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_961_root_address_inst_ack_0, ack => cp_elements(501)); -- 
    plus_base_cr_2585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => array_obj_ref_961_root_address_inst_req_1); -- 
    plus_base_ca_2586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_961_root_address_inst_ack_1, ack => cp_elements(502)); -- 
    final_reg_ack_2591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_961_final_reg_ack_0, ack => cp_elements(503)); -- 
    base_resize_req_2605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => ptr_deref_964_base_resize_req_0); -- 
    cp_elements(504) <= cp_elements(496);
    cpelement_group_505 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(504) & cp_elements(520));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(505),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => ptr_deref_964_gather_scatter_req_0); -- 
    base_resize_ack_2606_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_base_resize_ack_0, ack => cp_elements(506)); -- 
    sum_rename_req_2610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_964_root_address_inst_req_0); -- 
    cp_elements(507) <= ptr_deref_964_root_address_inst_ack_0;
    cp_elements(508) <= cp_elements(507);
    rr_2618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(508), ack => ptr_deref_964_addr_0_req_0); -- 
    ra_2619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_0_ack_0, ack => cp_elements(509)); -- 
    cr_2620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ptr_deref_964_addr_0_req_1); -- 
    ca_2621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_0_ack_1, ack => cp_elements(510)); -- 
    cp_elements(511) <= cp_elements(507);
    rr_2625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(511), ack => ptr_deref_964_addr_1_req_0); -- 
    ra_2626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_1_ack_0, ack => cp_elements(512)); -- 
    cr_2627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(512), ack => ptr_deref_964_addr_1_req_1); -- 
    ca_2628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_1_ack_1, ack => cp_elements(513)); -- 
    cp_elements(514) <= cp_elements(507);
    rr_2632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => ptr_deref_964_addr_2_req_0); -- 
    ra_2633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_2_ack_0, ack => cp_elements(515)); -- 
    cr_2634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => ptr_deref_964_addr_2_req_1); -- 
    ca_2635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_2_ack_1, ack => cp_elements(516)); -- 
    cp_elements(517) <= cp_elements(507);
    rr_2639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => ptr_deref_964_addr_3_req_0); -- 
    ra_2640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_3_ack_0, ack => cp_elements(518)); -- 
    cr_2641_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(518), ack => ptr_deref_964_addr_3_req_1); -- 
    ca_2642_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_addr_3_ack_1, ack => cp_elements(519)); -- 
    cpelement_group_520 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(510) & cp_elements(513) & cp_elements(516) & cp_elements(519));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(520),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(521) <= ptr_deref_964_gather_scatter_ack_0;
    cp_elements(522) <= cp_elements(521);
    rr_2654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(522), ack => ptr_deref_964_store_0_req_0); -- 
    ra_2655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_0_ack_0, ack => cp_elements(523)); -- 
    cp_elements(524) <= cp_elements(521);
    rr_2659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => ptr_deref_964_store_1_req_0); -- 
    ra_2660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_1_ack_0, ack => cp_elements(525)); -- 
    cp_elements(526) <= cp_elements(521);
    rr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(526), ack => ptr_deref_964_store_2_req_0); -- 
    ra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_2_ack_0, ack => cp_elements(527)); -- 
    cp_elements(528) <= cp_elements(521);
    rr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => ptr_deref_964_store_3_req_0); -- 
    ra_2670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_3_ack_0, ack => cp_elements(529)); -- 
    cpelement_group_530 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(523) & cp_elements(525) & cp_elements(527) & cp_elements(529));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(530),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(531) <= cp_elements(530);
    cp_elements(532) <= cp_elements(531);
    cr_2680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => ptr_deref_964_store_0_req_1); -- 
    ca_2681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_0_ack_1, ack => cp_elements(533)); -- 
    cp_elements(534) <= cp_elements(531);
    cr_2685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => ptr_deref_964_store_1_req_1); -- 
    ca_2686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_1_ack_1, ack => cp_elements(535)); -- 
    cp_elements(536) <= cp_elements(531);
    cr_2690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(536), ack => ptr_deref_964_store_2_req_1); -- 
    ca_2691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_2_ack_1, ack => cp_elements(537)); -- 
    cp_elements(538) <= cp_elements(531);
    cr_2695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => ptr_deref_964_store_3_req_1); -- 
    ca_2696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_964_store_3_ack_1, ack => cp_elements(539)); -- 
    cpelement_group_540 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(533) & cp_elements(535) & cp_elements(537) & cp_elements(539));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(540),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_541 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(542) & cp_elements(543));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(541),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => binary_971_inst_req_0); -- 
    cp_elements(542) <= cp_elements(496);
    cp_elements(543) <= cp_elements(496);
    ra_2706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_971_inst_ack_0, ack => cp_elements(544)); -- 
    cr_2707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(544), ack => binary_971_inst_req_1); -- 
    ca_2708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_971_inst_ack_1, ack => cp_elements(545)); -- 
    index_resize_req_2723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => array_obj_ref_975_index_0_resize_req_0); -- 
    cp_elements(546) <= cp_elements(496);
    cpelement_group_547 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(546) & cp_elements(555));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(547),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => array_obj_ref_975_final_reg_req_0); -- 
    cp_elements(548) <= cp_elements(496);
    base_resize_req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => array_obj_ref_975_base_resize_req_0); -- 
    index_resize_ack_2724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_index_0_resize_ack_0, ack => cp_elements(549)); -- 
    scale_rename_req_2728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => array_obj_ref_975_index_0_rename_req_0); -- 
    scale_rename_ack_2729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_index_0_rename_ack_0, ack => cp_elements(550)); -- 
    final_index_req_2733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => array_obj_ref_975_offset_inst_req_0); -- 
    final_index_ack_2734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_offset_inst_ack_0, ack => cp_elements(551)); -- 
    base_resize_ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_base_resize_ack_0, ack => cp_elements(552)); -- 
    cpelement_group_553 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(551) & cp_elements(552));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(553),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_2745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(553), ack => array_obj_ref_975_root_address_inst_req_0); -- 
    plus_base_ra_2746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_root_address_inst_ack_0, ack => cp_elements(554)); -- 
    plus_base_cr_2747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => array_obj_ref_975_root_address_inst_req_1); -- 
    plus_base_ca_2748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_root_address_inst_ack_1, ack => cp_elements(555)); -- 
    final_reg_ack_2753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_975_final_reg_ack_0, ack => cp_elements(556)); -- 
    cp_elements(557) <= cp_elements(496);
    cpelement_group_558 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(557) & cp_elements(562));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(558),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_2777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(558), ack => array_obj_ref_982_final_reg_req_0); -- 
    cp_elements(559) <= cp_elements(496);
    base_resize_req_2764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => array_obj_ref_982_base_resize_req_0); -- 
    base_resize_ack_2765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_982_base_resize_ack_0, ack => cp_elements(560)); -- 
    plus_base_rr_2770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(560), ack => array_obj_ref_982_root_address_inst_req_0); -- 
    plus_base_ra_2771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_982_root_address_inst_ack_0, ack => cp_elements(561)); -- 
    plus_base_cr_2772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => array_obj_ref_982_root_address_inst_req_1); -- 
    plus_base_ca_2773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_982_root_address_inst_ack_1, ack => cp_elements(562)); -- 
    cp_elements(563) <= array_obj_ref_982_final_reg_ack_0;
    cpelement_group_564 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(530) & cp_elements(556) & cp_elements(563) & cp_elements(580));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(564),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_2833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => ptr_deref_985_gather_scatter_req_0); -- 
    cp_elements(565) <= cp_elements(563);
    base_resize_req_2792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => ptr_deref_985_base_resize_req_0); -- 
    base_resize_ack_2793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_base_resize_ack_0, ack => cp_elements(566)); -- 
    sum_rename_req_2797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => ptr_deref_985_root_address_inst_req_0); -- 
    cp_elements(567) <= ptr_deref_985_root_address_inst_ack_0;
    cp_elements(568) <= cp_elements(567);
    rr_2805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_985_addr_0_req_0); -- 
    ra_2806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_0_ack_0, ack => cp_elements(569)); -- 
    cr_2807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => ptr_deref_985_addr_0_req_1); -- 
    ca_2808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_0_ack_1, ack => cp_elements(570)); -- 
    cp_elements(571) <= cp_elements(567);
    rr_2812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => ptr_deref_985_addr_1_req_0); -- 
    ra_2813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_1_ack_0, ack => cp_elements(572)); -- 
    cr_2814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(572), ack => ptr_deref_985_addr_1_req_1); -- 
    ca_2815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_1_ack_1, ack => cp_elements(573)); -- 
    cp_elements(574) <= cp_elements(567);
    rr_2819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => ptr_deref_985_addr_2_req_0); -- 
    ra_2820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_2_ack_0, ack => cp_elements(575)); -- 
    cr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => ptr_deref_985_addr_2_req_1); -- 
    ca_2822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_2_ack_1, ack => cp_elements(576)); -- 
    cp_elements(577) <= cp_elements(567);
    rr_2826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => ptr_deref_985_addr_3_req_0); -- 
    ra_2827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_3_ack_0, ack => cp_elements(578)); -- 
    cr_2828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => ptr_deref_985_addr_3_req_1); -- 
    ca_2829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_addr_3_ack_1, ack => cp_elements(579)); -- 
    cpelement_group_580 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(570) & cp_elements(573) & cp_elements(576) & cp_elements(579));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(580),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(581) <= ptr_deref_985_gather_scatter_ack_0;
    cp_elements(582) <= cp_elements(581);
    rr_2841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(582), ack => ptr_deref_985_store_0_req_0); -- 
    ra_2842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_0_ack_0, ack => cp_elements(583)); -- 
    cp_elements(584) <= cp_elements(581);
    rr_2846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => ptr_deref_985_store_1_req_0); -- 
    ra_2847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_1_ack_0, ack => cp_elements(585)); -- 
    cp_elements(586) <= cp_elements(581);
    rr_2851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ptr_deref_985_store_2_req_0); -- 
    ra_2852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_2_ack_0, ack => cp_elements(587)); -- 
    cp_elements(588) <= cp_elements(581);
    rr_2856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(588), ack => ptr_deref_985_store_3_req_0); -- 
    ra_2857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_3_ack_0, ack => cp_elements(589)); -- 
    cpelement_group_590 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(583) & cp_elements(585) & cp_elements(587) & cp_elements(589));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(590),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(591) <= cp_elements(590);
    cr_2867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => ptr_deref_985_store_0_req_1); -- 
    ca_2868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_0_ack_1, ack => cp_elements(592)); -- 
    cp_elements(593) <= cp_elements(590);
    cr_2872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_985_store_1_req_1); -- 
    ca_2873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_1_ack_1, ack => cp_elements(594)); -- 
    cp_elements(595) <= cp_elements(590);
    cr_2877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => ptr_deref_985_store_2_req_1); -- 
    ca_2878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_2_ack_1, ack => cp_elements(596)); -- 
    cp_elements(597) <= cp_elements(590);
    cr_2882_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(597), ack => ptr_deref_985_store_3_req_1); -- 
    ca_2883_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_985_store_3_ack_1, ack => cp_elements(598)); -- 
    cpelement_group_599 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(592) & cp_elements(594) & cp_elements(596) & cp_elements(598));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(599),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_600 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(601) & cp_elements(602) & cp_elements(603));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => binary_991_inst_req_0); -- 
    cp_elements(601) <= cp_elements(496);
    cp_elements(602) <= cp_elements(496);
    cp_elements(603) <= cp_elements(496);
    ra_2894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_991_inst_ack_0, ack => cp_elements(604)); -- 
    cr_2895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => binary_991_inst_req_1); -- 
    ca_2896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_991_inst_ack_1, ack => cp_elements(605)); -- 
    cpelement_group_606 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(540) & cp_elements(599) & cp_elements(605));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(606),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(607) <= cp_elements(14);
    cp_elements(608) <= false;
    cp_elements(609) <= cp_elements(608);
    cp_elements(610) <= cp_elements(14);
    branch_req_2904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(610), ack => if_stmt_993_branch_req_0); -- 
    cp_elements(611) <= cp_elements(610);
    cp_elements(612) <= cp_elements(611);
    if_choice_transition_2909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_993_branch_ack_1, ack => cp_elements(613)); -- 
    cp_elements(614) <= cp_elements(611);
    else_choice_transition_2913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_993_branch_ack_0, ack => cp_elements(615)); -- 
    cp_elements(616) <= cp_elements(15);
    cpelement_group_617 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(618) & cp_elements(619) & cp_elements(620));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(617),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(617), ack => binary_1003_inst_req_0); -- 
    cp_elements(618) <= cp_elements(616);
    cp_elements(619) <= cp_elements(616);
    cp_elements(620) <= cp_elements(616);
    ra_2929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1003_inst_ack_0, ack => cp_elements(621)); -- 
    cr_2930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => binary_1003_inst_req_1); -- 
    cp_elements(622) <= binary_1003_inst_ack_1;
    cpelement_group_623 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(624) & cp_elements(625) & cp_elements(626));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(623),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(623), ack => binary_1008_inst_req_0); -- 
    cp_elements(624) <= cp_elements(616);
    cp_elements(625) <= cp_elements(616);
    cp_elements(626) <= cp_elements(622);
    ra_2942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1008_inst_ack_0, ack => cp_elements(627)); -- 
    cr_2943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => binary_1008_inst_req_1); -- 
    ca_2944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1008_inst_ack_1, ack => cp_elements(628)); -- 
    cp_elements(629) <= cp_elements(616);
    cpelement_group_630 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(628) & cp_elements(629) & cp_elements(631) & cp_elements(632));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(630),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_2955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => ternary_1014_inst_req_0); -- 
    cp_elements(631) <= cp_elements(616);
    cp_elements(632) <= cp_elements(622);
    ack_2956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ternary_1014_inst_ack_0, ack => cp_elements(633)); -- 
    cpelement_group_634 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(633) & cp_elements(635));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(634),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_2965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(634), ack => binary_1020_inst_req_0); -- 
    cp_elements(635) <= cp_elements(616);
    ra_2966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1020_inst_ack_0, ack => cp_elements(636)); -- 
    cr_2967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => binary_1020_inst_req_1); -- 
    ca_2968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1020_inst_ack_1, ack => cp_elements(637)); -- 
    index_resize_req_2983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(637), ack => array_obj_ref_1024_index_0_resize_req_0); -- 
    cp_elements(638) <= cp_elements(616);
    cpelement_group_639 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(638) & cp_elements(647));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(639),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => array_obj_ref_1024_final_reg_req_0); -- 
    cp_elements(640) <= cp_elements(616);
    base_resize_req_2999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => array_obj_ref_1024_base_resize_req_0); -- 
    index_resize_ack_2984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_index_0_resize_ack_0, ack => cp_elements(641)); -- 
    scale_rename_req_2988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(641), ack => array_obj_ref_1024_index_0_rename_req_0); -- 
    scale_rename_ack_2989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_index_0_rename_ack_0, ack => cp_elements(642)); -- 
    final_index_req_2993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => array_obj_ref_1024_offset_inst_req_0); -- 
    final_index_ack_2994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_offset_inst_ack_0, ack => cp_elements(643)); -- 
    base_resize_ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_base_resize_ack_0, ack => cp_elements(644)); -- 
    cpelement_group_645 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(643) & cp_elements(644));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(645),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_3005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => array_obj_ref_1024_root_address_inst_req_0); -- 
    plus_base_ra_3006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_root_address_inst_ack_0, ack => cp_elements(646)); -- 
    plus_base_cr_3007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(646), ack => array_obj_ref_1024_root_address_inst_req_1); -- 
    plus_base_ca_3008_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_root_address_inst_ack_1, ack => cp_elements(647)); -- 
    final_reg_ack_3013_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1024_final_reg_ack_0, ack => cp_elements(648)); -- 
    cpelement_group_649 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(648) & cp_elements(650) & cp_elements(666));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(649),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(649), ack => ptr_deref_1027_gather_scatter_req_0); -- 
    cp_elements(650) <= cp_elements(616);
    cp_elements(651) <= cp_elements(650);
    base_resize_req_3027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(651), ack => ptr_deref_1027_base_resize_req_0); -- 
    base_resize_ack_3028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_base_resize_ack_0, ack => cp_elements(652)); -- 
    sum_rename_req_3032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_1027_root_address_inst_req_0); -- 
    cp_elements(653) <= ptr_deref_1027_root_address_inst_ack_0;
    cp_elements(654) <= cp_elements(653);
    rr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_1027_addr_0_req_0); -- 
    ra_3041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_0_ack_0, ack => cp_elements(655)); -- 
    cr_3042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => ptr_deref_1027_addr_0_req_1); -- 
    ca_3043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_0_ack_1, ack => cp_elements(656)); -- 
    cp_elements(657) <= cp_elements(653);
    rr_3047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(657), ack => ptr_deref_1027_addr_1_req_0); -- 
    ra_3048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_1_ack_0, ack => cp_elements(658)); -- 
    cr_3049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => ptr_deref_1027_addr_1_req_1); -- 
    ca_3050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_1_ack_1, ack => cp_elements(659)); -- 
    cp_elements(660) <= cp_elements(653);
    rr_3054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => ptr_deref_1027_addr_2_req_0); -- 
    ra_3055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_2_ack_0, ack => cp_elements(661)); -- 
    cr_3056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(661), ack => ptr_deref_1027_addr_2_req_1); -- 
    ca_3057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_2_ack_1, ack => cp_elements(662)); -- 
    cp_elements(663) <= cp_elements(653);
    rr_3061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => ptr_deref_1027_addr_3_req_0); -- 
    ra_3062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_3_ack_0, ack => cp_elements(664)); -- 
    cr_3063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(664), ack => ptr_deref_1027_addr_3_req_1); -- 
    ca_3064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_addr_3_ack_1, ack => cp_elements(665)); -- 
    cpelement_group_666 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(656) & cp_elements(659) & cp_elements(662) & cp_elements(665));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(666),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(667) <= ptr_deref_1027_gather_scatter_ack_0;
    cp_elements(668) <= cp_elements(667);
    rr_3076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => ptr_deref_1027_store_0_req_0); -- 
    ra_3077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_0_ack_0, ack => cp_elements(669)); -- 
    cp_elements(670) <= cp_elements(667);
    rr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(670), ack => ptr_deref_1027_store_1_req_0); -- 
    ra_3082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_1_ack_0, ack => cp_elements(671)); -- 
    cp_elements(672) <= cp_elements(667);
    rr_3086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(672), ack => ptr_deref_1027_store_2_req_0); -- 
    ra_3087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_2_ack_0, ack => cp_elements(673)); -- 
    cp_elements(674) <= cp_elements(667);
    rr_3091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(674), ack => ptr_deref_1027_store_3_req_0); -- 
    ra_3092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_3_ack_0, ack => cp_elements(675)); -- 
    cpelement_group_676 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(669) & cp_elements(671) & cp_elements(673) & cp_elements(675));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(676),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(677) <= cp_elements(676);
    cp_elements(678) <= cp_elements(677);
    cr_3102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => ptr_deref_1027_store_0_req_1); -- 
    ca_3103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_0_ack_1, ack => cp_elements(679)); -- 
    cp_elements(680) <= cp_elements(677);
    cr_3107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => ptr_deref_1027_store_1_req_1); -- 
    ca_3108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_1_ack_1, ack => cp_elements(681)); -- 
    cp_elements(682) <= cp_elements(677);
    cr_3112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => ptr_deref_1027_store_2_req_1); -- 
    ca_3113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_2_ack_1, ack => cp_elements(683)); -- 
    cp_elements(684) <= cp_elements(677);
    cr_3117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_1027_store_3_req_1); -- 
    ca_3118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1027_store_3_ack_1, ack => cp_elements(685)); -- 
    cpelement_group_686 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(679) & cp_elements(681) & cp_elements(683) & cp_elements(685));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(686),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(687) <= cp_elements(616);
    cpelement_group_688 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(687) & cp_elements(692));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(688), ack => array_obj_ref_1033_final_reg_req_0); -- 
    cp_elements(689) <= cp_elements(616);
    base_resize_req_3129_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(689), ack => array_obj_ref_1033_base_resize_req_0); -- 
    base_resize_ack_3130_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1033_base_resize_ack_0, ack => cp_elements(690)); -- 
    plus_base_rr_3135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => array_obj_ref_1033_root_address_inst_req_0); -- 
    plus_base_ra_3136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1033_root_address_inst_ack_0, ack => cp_elements(691)); -- 
    plus_base_cr_3137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(691), ack => array_obj_ref_1033_root_address_inst_req_1); -- 
    plus_base_ca_3138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1033_root_address_inst_ack_1, ack => cp_elements(692)); -- 
    final_reg_ack_3143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1033_final_reg_ack_0, ack => cp_elements(693)); -- 
    cpelement_group_694 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(693) & cp_elements(695));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(694),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => type_cast_1037_inst_req_0); -- 
    cp_elements(695) <= cp_elements(616);
    cp_elements(696) <= type_cast_1037_inst_ack_0;
    cpelement_group_697 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(676) & cp_elements(696) & cp_elements(713));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(697),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(698) <= cp_elements(696);
    base_resize_req_3166_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(698), ack => ptr_deref_1041_base_resize_req_0); -- 
    base_resize_ack_3167_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_base_resize_ack_0, ack => cp_elements(699)); -- 
    sum_rename_req_3171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_1041_root_address_inst_req_0); -- 
    cp_elements(700) <= ptr_deref_1041_root_address_inst_ack_0;
    cp_elements(701) <= cp_elements(700);
    rr_3179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_1041_addr_0_req_0); -- 
    ra_3180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_0_ack_0, ack => cp_elements(702)); -- 
    cr_3181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => ptr_deref_1041_addr_0_req_1); -- 
    ca_3182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_0_ack_1, ack => cp_elements(703)); -- 
    cp_elements(704) <= cp_elements(700);
    rr_3186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(704), ack => ptr_deref_1041_addr_1_req_0); -- 
    ra_3187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_1_ack_0, ack => cp_elements(705)); -- 
    cr_3188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => ptr_deref_1041_addr_1_req_1); -- 
    ca_3189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_1_ack_1, ack => cp_elements(706)); -- 
    cp_elements(707) <= cp_elements(700);
    rr_3193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => ptr_deref_1041_addr_2_req_0); -- 
    ra_3194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_2_ack_0, ack => cp_elements(708)); -- 
    cr_3195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => ptr_deref_1041_addr_2_req_1); -- 
    ca_3196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_2_ack_1, ack => cp_elements(709)); -- 
    cp_elements(710) <= cp_elements(700);
    rr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => ptr_deref_1041_addr_3_req_0); -- 
    ra_3201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_3_ack_0, ack => cp_elements(711)); -- 
    cr_3202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => ptr_deref_1041_addr_3_req_1); -- 
    ca_3203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_addr_3_ack_1, ack => cp_elements(712)); -- 
    cpelement_group_713 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(703) & cp_elements(706) & cp_elements(709) & cp_elements(712));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(713),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(714) <= cp_elements(697);
    rr_3213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(714), ack => ptr_deref_1041_load_0_req_0); -- 
    ra_3214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_0_ack_0, ack => cp_elements(715)); -- 
    cp_elements(716) <= cp_elements(697);
    rr_3218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(716), ack => ptr_deref_1041_load_1_req_0); -- 
    ra_3219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_1_ack_0, ack => cp_elements(717)); -- 
    cp_elements(718) <= cp_elements(697);
    rr_3223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(718), ack => ptr_deref_1041_load_2_req_0); -- 
    ra_3224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_2_ack_0, ack => cp_elements(719)); -- 
    cp_elements(720) <= cp_elements(697);
    rr_3228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => ptr_deref_1041_load_3_req_0); -- 
    ra_3229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_3_ack_0, ack => cp_elements(721)); -- 
    cpelement_group_722 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(715) & cp_elements(717) & cp_elements(719) & cp_elements(721));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(722),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(723) <= cp_elements(722);
    cr_3239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(723), ack => ptr_deref_1041_load_0_req_1); -- 
    ca_3240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_0_ack_1, ack => cp_elements(724)); -- 
    cp_elements(725) <= cp_elements(722);
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => ptr_deref_1041_load_1_req_1); -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_1_ack_1, ack => cp_elements(726)); -- 
    cp_elements(727) <= cp_elements(722);
    cr_3249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => ptr_deref_1041_load_2_req_1); -- 
    ca_3250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_2_ack_1, ack => cp_elements(728)); -- 
    cp_elements(729) <= cp_elements(722);
    cr_3254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => ptr_deref_1041_load_3_req_1); -- 
    ca_3255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_load_3_ack_1, ack => cp_elements(730)); -- 
    cpelement_group_731 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(724) & cp_elements(726) & cp_elements(728) & cp_elements(730));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(731),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_3256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(731), ack => ptr_deref_1041_gather_scatter_req_0); -- 
    merge_ack_3257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1041_gather_scatter_ack_0, ack => cp_elements(732)); -- 
    cp_elements(733) <= cp_elements(616);
    cpelement_group_734 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(733) & cp_elements(738));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(734),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => array_obj_ref_1048_final_reg_req_0); -- 
    cp_elements(735) <= cp_elements(616);
    base_resize_req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => array_obj_ref_1048_base_resize_req_0); -- 
    base_resize_ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_base_resize_ack_0, ack => cp_elements(736)); -- 
    plus_base_rr_3274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => array_obj_ref_1048_root_address_inst_req_0); -- 
    plus_base_ra_3275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_root_address_inst_ack_0, ack => cp_elements(737)); -- 
    plus_base_cr_3276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => array_obj_ref_1048_root_address_inst_req_1); -- 
    plus_base_ca_3277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_root_address_inst_ack_1, ack => cp_elements(738)); -- 
    final_reg_ack_3282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1048_final_reg_ack_0, ack => cp_elements(739)); -- 
    cpelement_group_740 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(739) & cp_elements(741));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(740),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => type_cast_1052_inst_req_0); -- 
    cp_elements(741) <= cp_elements(616);
    cp_elements(742) <= type_cast_1052_inst_ack_0;
    cpelement_group_743 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(732) & cp_elements(742) & cp_elements(759));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(743),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => ptr_deref_1055_gather_scatter_req_0); -- 
    cp_elements(744) <= cp_elements(742);
    base_resize_req_3306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => ptr_deref_1055_base_resize_req_0); -- 
    base_resize_ack_3307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_base_resize_ack_0, ack => cp_elements(745)); -- 
    sum_rename_req_3311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => ptr_deref_1055_root_address_inst_req_0); -- 
    cp_elements(746) <= ptr_deref_1055_root_address_inst_ack_0;
    cp_elements(747) <= cp_elements(746);
    rr_3319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(747), ack => ptr_deref_1055_addr_0_req_0); -- 
    ra_3320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_0_ack_0, ack => cp_elements(748)); -- 
    cr_3321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(748), ack => ptr_deref_1055_addr_0_req_1); -- 
    ca_3322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_0_ack_1, ack => cp_elements(749)); -- 
    cp_elements(750) <= cp_elements(746);
    rr_3326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(750), ack => ptr_deref_1055_addr_1_req_0); -- 
    ra_3327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_1_ack_0, ack => cp_elements(751)); -- 
    cr_3328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(751), ack => ptr_deref_1055_addr_1_req_1); -- 
    ca_3329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_1_ack_1, ack => cp_elements(752)); -- 
    cp_elements(753) <= cp_elements(746);
    rr_3333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ptr_deref_1055_addr_2_req_0); -- 
    ra_3334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_2_ack_0, ack => cp_elements(754)); -- 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(754), ack => ptr_deref_1055_addr_2_req_1); -- 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_2_ack_1, ack => cp_elements(755)); -- 
    cp_elements(756) <= cp_elements(746);
    rr_3340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => ptr_deref_1055_addr_3_req_0); -- 
    ra_3341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_3_ack_0, ack => cp_elements(757)); -- 
    cr_3342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => ptr_deref_1055_addr_3_req_1); -- 
    ca_3343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_addr_3_ack_1, ack => cp_elements(758)); -- 
    cpelement_group_759 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(749) & cp_elements(752) & cp_elements(755) & cp_elements(758));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(759),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(760) <= ptr_deref_1055_gather_scatter_ack_0;
    cp_elements(761) <= cp_elements(760);
    rr_3355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => ptr_deref_1055_store_0_req_0); -- 
    ra_3356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_0_ack_0, ack => cp_elements(762)); -- 
    cp_elements(763) <= cp_elements(760);
    rr_3360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => ptr_deref_1055_store_1_req_0); -- 
    ra_3361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_1_ack_0, ack => cp_elements(764)); -- 
    cp_elements(765) <= cp_elements(760);
    rr_3365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => ptr_deref_1055_store_2_req_0); -- 
    ra_3366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_2_ack_0, ack => cp_elements(766)); -- 
    cp_elements(767) <= cp_elements(760);
    rr_3370_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => ptr_deref_1055_store_3_req_0); -- 
    ra_3371_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_3_ack_0, ack => cp_elements(768)); -- 
    cpelement_group_769 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(762) & cp_elements(764) & cp_elements(766) & cp_elements(768));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(769),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(770) <= cp_elements(769);
    cr_3381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => ptr_deref_1055_store_0_req_1); -- 
    ca_3382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_0_ack_1, ack => cp_elements(771)); -- 
    cp_elements(772) <= cp_elements(769);
    cr_3386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => ptr_deref_1055_store_1_req_1); -- 
    ca_3387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_1_ack_1, ack => cp_elements(773)); -- 
    cp_elements(774) <= cp_elements(769);
    cr_3391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => ptr_deref_1055_store_2_req_1); -- 
    ca_3392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_2_ack_1, ack => cp_elements(775)); -- 
    cp_elements(776) <= cp_elements(769);
    cr_3396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => ptr_deref_1055_store_3_req_1); -- 
    ca_3397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1055_store_3_ack_1, ack => cp_elements(777)); -- 
    cpelement_group_778 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(771) & cp_elements(773) & cp_elements(775) & cp_elements(777));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(778),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_779 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(686) & cp_elements(778));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(779),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(780) <= cp_elements(615);
    cp_elements(781) <= cp_elements(780);
    cpelement_group_782 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(781) & cp_elements(786));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(782),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(782), ack => array_obj_ref_1063_final_reg_req_0); -- 
    cp_elements(783) <= cp_elements(780);
    base_resize_req_3411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => array_obj_ref_1063_base_resize_req_0); -- 
    base_resize_ack_3412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_base_resize_ack_0, ack => cp_elements(784)); -- 
    plus_base_rr_3417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => array_obj_ref_1063_root_address_inst_req_0); -- 
    plus_base_ra_3418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_root_address_inst_ack_0, ack => cp_elements(785)); -- 
    plus_base_cr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => array_obj_ref_1063_root_address_inst_req_1); -- 
    plus_base_ca_3420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_root_address_inst_ack_1, ack => cp_elements(786)); -- 
    final_reg_ack_3425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1063_final_reg_ack_0, ack => cp_elements(787)); -- 
    cpelement_group_788 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(787) & cp_elements(789));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(788),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => type_cast_1067_inst_req_0); -- 
    cp_elements(789) <= cp_elements(780);
    ack_3435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1067_inst_ack_0, ack => cp_elements(790)); -- 
    base_resize_req_3448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => ptr_deref_1071_base_resize_req_0); -- 
    base_resize_ack_3449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_base_resize_ack_0, ack => cp_elements(791)); -- 
    sum_rename_req_3453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => ptr_deref_1071_root_address_inst_req_0); -- 
    cp_elements(792) <= ptr_deref_1071_root_address_inst_ack_0;
    cp_elements(793) <= cp_elements(792);
    rr_3461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => ptr_deref_1071_addr_0_req_0); -- 
    ra_3462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_0_ack_0, ack => cp_elements(794)); -- 
    cr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => ptr_deref_1071_addr_0_req_1); -- 
    ca_3464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_0_ack_1, ack => cp_elements(795)); -- 
    cp_elements(796) <= cp_elements(792);
    rr_3468_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => ptr_deref_1071_addr_1_req_0); -- 
    ra_3469_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_1_ack_0, ack => cp_elements(797)); -- 
    cr_3470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => ptr_deref_1071_addr_1_req_1); -- 
    ca_3471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_1_ack_1, ack => cp_elements(798)); -- 
    cp_elements(799) <= cp_elements(792);
    rr_3475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => ptr_deref_1071_addr_2_req_0); -- 
    ra_3476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_2_ack_0, ack => cp_elements(800)); -- 
    cr_3477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => ptr_deref_1071_addr_2_req_1); -- 
    ca_3478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_2_ack_1, ack => cp_elements(801)); -- 
    cp_elements(802) <= cp_elements(792);
    rr_3482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(802), ack => ptr_deref_1071_addr_3_req_0); -- 
    ra_3483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_3_ack_0, ack => cp_elements(803)); -- 
    cr_3484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => ptr_deref_1071_addr_3_req_1); -- 
    ca_3485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_addr_3_ack_1, ack => cp_elements(804)); -- 
    cpelement_group_805 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(795) & cp_elements(798) & cp_elements(801) & cp_elements(804));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(805),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(806) <= cp_elements(805);
    rr_3495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_1071_load_0_req_0); -- 
    ra_3496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_0_ack_0, ack => cp_elements(807)); -- 
    cp_elements(808) <= cp_elements(805);
    rr_3500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => ptr_deref_1071_load_1_req_0); -- 
    ra_3501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_1_ack_0, ack => cp_elements(809)); -- 
    cp_elements(810) <= cp_elements(805);
    rr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => ptr_deref_1071_load_2_req_0); -- 
    ra_3506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_2_ack_0, ack => cp_elements(811)); -- 
    cp_elements(812) <= cp_elements(805);
    rr_3510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => ptr_deref_1071_load_3_req_0); -- 
    ra_3511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_3_ack_0, ack => cp_elements(813)); -- 
    cpelement_group_814 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(807) & cp_elements(809) & cp_elements(811) & cp_elements(813));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(814),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(815) <= cp_elements(814);
    cr_3521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => ptr_deref_1071_load_0_req_1); -- 
    ca_3522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_0_ack_1, ack => cp_elements(816)); -- 
    cp_elements(817) <= cp_elements(814);
    cr_3526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(817), ack => ptr_deref_1071_load_1_req_1); -- 
    ca_3527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_1_ack_1, ack => cp_elements(818)); -- 
    cp_elements(819) <= cp_elements(814);
    cr_3531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => ptr_deref_1071_load_2_req_1); -- 
    ca_3532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_2_ack_1, ack => cp_elements(820)); -- 
    cp_elements(821) <= cp_elements(814);
    cr_3536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => ptr_deref_1071_load_3_req_1); -- 
    ca_3537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_load_3_ack_1, ack => cp_elements(822)); -- 
    cpelement_group_823 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(816) & cp_elements(818) & cp_elements(820) & cp_elements(822));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(823),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_3538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => ptr_deref_1071_gather_scatter_req_0); -- 
    merge_ack_3539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1071_gather_scatter_ack_0, ack => cp_elements(824)); -- 
    cp_elements(825) <= cp_elements(780);
    cpelement_group_826 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(825) & cp_elements(830));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(826),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_3563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => array_obj_ref_1078_final_reg_req_0); -- 
    cp_elements(827) <= cp_elements(780);
    base_resize_req_3550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => array_obj_ref_1078_base_resize_req_0); -- 
    base_resize_ack_3551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_base_resize_ack_0, ack => cp_elements(828)); -- 
    plus_base_rr_3556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => array_obj_ref_1078_root_address_inst_req_0); -- 
    plus_base_ra_3557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_root_address_inst_ack_0, ack => cp_elements(829)); -- 
    plus_base_cr_3558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(829), ack => array_obj_ref_1078_root_address_inst_req_1); -- 
    plus_base_ca_3559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_root_address_inst_ack_1, ack => cp_elements(830)); -- 
    final_reg_ack_3564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1078_final_reg_ack_0, ack => cp_elements(831)); -- 
    cpelement_group_832 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(831) & cp_elements(833));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(832),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3573_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(832), ack => type_cast_1082_inst_req_0); -- 
    cp_elements(833) <= cp_elements(780);
    cp_elements(834) <= type_cast_1082_inst_ack_0;
    cpelement_group_835 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(824) & cp_elements(834) & cp_elements(851));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_3629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => ptr_deref_1085_gather_scatter_req_0); -- 
    cp_elements(836) <= cp_elements(834);
    base_resize_req_3588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(836), ack => ptr_deref_1085_base_resize_req_0); -- 
    base_resize_ack_3589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_base_resize_ack_0, ack => cp_elements(837)); -- 
    sum_rename_req_3593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(837), ack => ptr_deref_1085_root_address_inst_req_0); -- 
    cp_elements(838) <= ptr_deref_1085_root_address_inst_ack_0;
    cp_elements(839) <= cp_elements(838);
    rr_3601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(839), ack => ptr_deref_1085_addr_0_req_0); -- 
    ra_3602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_0_ack_0, ack => cp_elements(840)); -- 
    cr_3603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => ptr_deref_1085_addr_0_req_1); -- 
    ca_3604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_0_ack_1, ack => cp_elements(841)); -- 
    cp_elements(842) <= cp_elements(838);
    rr_3608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(842), ack => ptr_deref_1085_addr_1_req_0); -- 
    ra_3609_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_1_ack_0, ack => cp_elements(843)); -- 
    cr_3610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => ptr_deref_1085_addr_1_req_1); -- 
    ca_3611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_1_ack_1, ack => cp_elements(844)); -- 
    cp_elements(845) <= cp_elements(838);
    rr_3615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => ptr_deref_1085_addr_2_req_0); -- 
    ra_3616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_2_ack_0, ack => cp_elements(846)); -- 
    cr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(846), ack => ptr_deref_1085_addr_2_req_1); -- 
    ca_3618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_2_ack_1, ack => cp_elements(847)); -- 
    cp_elements(848) <= cp_elements(838);
    rr_3622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => ptr_deref_1085_addr_3_req_0); -- 
    ra_3623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_3_ack_0, ack => cp_elements(849)); -- 
    cr_3624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(849), ack => ptr_deref_1085_addr_3_req_1); -- 
    ca_3625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_addr_3_ack_1, ack => cp_elements(850)); -- 
    cpelement_group_851 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(841) & cp_elements(844) & cp_elements(847) & cp_elements(850));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(851),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(852) <= ptr_deref_1085_gather_scatter_ack_0;
    cp_elements(853) <= cp_elements(852);
    rr_3637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => ptr_deref_1085_store_0_req_0); -- 
    ra_3638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_0_ack_0, ack => cp_elements(854)); -- 
    cp_elements(855) <= cp_elements(852);
    rr_3642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(855), ack => ptr_deref_1085_store_1_req_0); -- 
    ra_3643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_1_ack_0, ack => cp_elements(856)); -- 
    cp_elements(857) <= cp_elements(852);
    rr_3647_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => ptr_deref_1085_store_2_req_0); -- 
    ra_3648_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_2_ack_0, ack => cp_elements(858)); -- 
    cp_elements(859) <= cp_elements(852);
    rr_3652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(859), ack => ptr_deref_1085_store_3_req_0); -- 
    ra_3653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_3_ack_0, ack => cp_elements(860)); -- 
    cpelement_group_861 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(854) & cp_elements(856) & cp_elements(858) & cp_elements(860));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(861),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(862) <= cp_elements(861);
    cr_3663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(862), ack => ptr_deref_1085_store_0_req_1); -- 
    ca_3664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_0_ack_1, ack => cp_elements(863)); -- 
    cp_elements(864) <= cp_elements(861);
    cr_3668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(864), ack => ptr_deref_1085_store_1_req_1); -- 
    ca_3669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_1_ack_1, ack => cp_elements(865)); -- 
    cp_elements(866) <= cp_elements(861);
    cr_3673_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(866), ack => ptr_deref_1085_store_2_req_1); -- 
    ca_3674_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_2_ack_1, ack => cp_elements(867)); -- 
    cp_elements(868) <= cp_elements(861);
    cr_3678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => ptr_deref_1085_store_3_req_1); -- 
    ca_3679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1085_store_3_ack_1, ack => cp_elements(869)); -- 
    cpelement_group_870 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(863) & cp_elements(865) & cp_elements(867) & cp_elements(869));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(870),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_871 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(872) & cp_elements(873));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(871),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_3688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => binary_1092_inst_req_0); -- 
    cp_elements(872) <= cp_elements(780);
    cp_elements(873) <= cp_elements(780);
    ra_3689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1092_inst_ack_0, ack => cp_elements(874)); -- 
    cr_3690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => binary_1092_inst_req_1); -- 
    ca_3691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1092_inst_ack_1, ack => cp_elements(875)); -- 
    cpelement_group_876 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(870) & cp_elements(875));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(876),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(877) <= cp_elements(17);
    cp_elements(878) <= false;
    cp_elements(879) <= cp_elements(878);
    cp_elements(880) <= cp_elements(17);
    branch_req_3699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(880), ack => if_stmt_1094_branch_req_0); -- 
    cp_elements(881) <= cp_elements(880);
    cp_elements(882) <= cp_elements(881);
    if_choice_transition_3704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1094_branch_ack_1, ack => cp_elements(883)); -- 
    cp_elements(884) <= cp_elements(881);
    else_choice_transition_3708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1094_branch_ack_0, ack => cp_elements(885)); -- 
    cp_elements(886) <= cp_elements(18);
    cpelement_group_887 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(888) & cp_elements(889));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(887),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(887), ack => type_cast_1103_inst_req_0); -- 
    cp_elements(888) <= cp_elements(886);
    cp_elements(889) <= cp_elements(886);
    ack_3723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1103_inst_ack_0, ack => cp_elements(890)); -- 
    cp_elements(891) <= cp_elements(890);
    cpelement_group_892 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(893) & cp_elements(894));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(892),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_3735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(892), ack => type_cast_1107_inst_req_0); -- 
    cp_elements(893) <= cp_elements(891);
    cp_elements(894) <= cp_elements(891);
    ack_3736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1107_inst_ack_0, ack => cp_elements(895)); -- 
    pipe_wreq_3741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(895), ack => simple_obj_ref_1105_inst_req_0); -- 
    pipe_wack_3742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1105_inst_ack_0, ack => cp_elements(896)); -- 
    cp_elements(897) <= false;
    cp_elements(898) <= cp_elements(897);
    cp_elements(899) <= false;
    cp_elements(900) <= cp_elements(899);
    cp_elements(901) <= false;
    cp_elements(902) <= cp_elements(901);
    cp_elements(903) <= false;
    cp_elements(904) <= cp_elements(903);
    cp_elements(905) <= false;
    cp_elements(906) <= cp_elements(905);
    cp_elements(907) <= cp_elements(398);
    cp_elements(908) <= cp_elements(907);
    req_3847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(908), ack => type_cast_760_inst_req_0); -- 
    ack_3848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_760_inst_ack_0, ack => cp_elements(909)); -- 
    phi_stmt_754_req_3849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => phi_stmt_754_req_1); -- 
    cp_elements(910) <= cp_elements(907);
    req_3859_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(910), ack => type_cast_767_inst_req_0); -- 
    ack_3860_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_767_inst_ack_0, ack => cp_elements(911)); -- 
    phi_stmt_761_req_3861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => phi_stmt_761_req_1); -- 
    cpelement_group_912 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(909) & cp_elements(911));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(912),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(913) <= cp_elements(316);
    cp_elements(914) <= cp_elements(913);
    phi_stmt_754_req_3876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(914), ack => phi_stmt_754_req_0); -- 
    cp_elements(915) <= cp_elements(913);
    phi_stmt_761_req_3888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(915), ack => phi_stmt_761_req_0); -- 
    cpelement_group_916 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(914) & cp_elements(915));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(916),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(917) <= OrReduce(cp_elements(912) & cp_elements(916));
    cp_elements(918) <= cp_elements(917);
    phi_stmt_754_ack_3893_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_754_ack_0, ack => cp_elements(919)); -- 
    phi_stmt_761_ack_3894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_761_ack_0, ack => cp_elements(920)); -- 
    cpelement_group_921 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(919) & cp_elements(920));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(921),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(922) <= false;
    cp_elements(923) <= cp_elements(922);
    cp_elements(924) <= cp_elements(310);
    cp_elements(925) <= cp_elements(924);
    phi_stmt_847_req_3921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(925), ack => phi_stmt_847_req_1); -- 
    cp_elements(926) <= cp_elements(924);
    cp_elements(927) <= cp_elements(926);
    cp_elements(928) <= cp_elements(926);
    req_3936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(928), ack => type_cast_859_inst_req_0); -- 
    ack_3937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_859_inst_ack_0, ack => cp_elements(929)); -- 
    cpelement_group_930 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(927) & cp_elements(929));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(930),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_854_req_3938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(930), ack => phi_stmt_854_req_1); -- 
    cp_elements(931) <= cp_elements(924);
    cp_elements(932) <= cp_elements(931);
    cp_elements(933) <= cp_elements(931);
    req_3953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(933), ack => type_cast_865_inst_req_0); -- 
    ack_3954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_865_inst_ack_0, ack => cp_elements(934)); -- 
    cpelement_group_935 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(932) & cp_elements(934));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(935),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_860_req_3955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => phi_stmt_860_req_1); -- 
    cpelement_group_936 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(925) & cp_elements(930) & cp_elements(935));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(936),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(937) <= cp_elements(417);
    cp_elements(938) <= cp_elements(937);
    req_3968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(938), ack => type_cast_850_inst_req_0); -- 
    ack_3969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_850_inst_ack_0, ack => cp_elements(939)); -- 
    phi_stmt_847_req_3970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => phi_stmt_847_req_0); -- 
    cp_elements(940) <= cp_elements(937);
    cp_elements(941) <= cp_elements(940);
    req_3980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(941), ack => type_cast_857_inst_req_0); -- 
    ack_3981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_857_inst_ack_0, ack => cp_elements(942)); -- 
    cp_elements(943) <= cp_elements(940);
    cpelement_group_944 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(942) & cp_elements(943));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(944),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_854_req_3987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => phi_stmt_854_req_0); -- 
    cp_elements(945) <= cp_elements(937);
    cp_elements(946) <= cp_elements(945);
    req_3997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(946), ack => type_cast_863_inst_req_0); -- 
    ack_3998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_863_inst_ack_0, ack => cp_elements(947)); -- 
    cp_elements(948) <= cp_elements(945);
    cpelement_group_949 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(947) & cp_elements(948));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(949),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_860_req_4004_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => phi_stmt_860_req_0); -- 
    cpelement_group_950 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(939) & cp_elements(944) & cp_elements(949));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(950),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(951) <= OrReduce(cp_elements(936) & cp_elements(950));
    cp_elements(952) <= cp_elements(951);
    phi_stmt_847_ack_4009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_847_ack_0, ack => cp_elements(953)); -- 
    phi_stmt_854_ack_4010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_854_ack_0, ack => cp_elements(954)); -- 
    phi_stmt_860_ack_4011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_860_ack_0, ack => cp_elements(955)); -- 
    cpelement_group_956 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(953) & cp_elements(954) & cp_elements(955));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(956),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(957) <= false;
    cp_elements(958) <= cp_elements(957);
    cp_elements(959) <= cp_elements(432);
    cp_elements(960) <= cp_elements(432);
    req_4041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(960), ack => type_cast_900_inst_req_0); -- 
    ack_4042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_900_inst_ack_0, ack => cp_elements(961)); -- 
    cpelement_group_962 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(959) & cp_elements(961));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(962),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_895_req_4043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => phi_stmt_895_req_1); -- 
    cp_elements(963) <= cp_elements(448);
    req_4056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(963), ack => type_cast_898_inst_req_0); -- 
    ack_4057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_898_inst_ack_0, ack => cp_elements(964)); -- 
    cp_elements(965) <= cp_elements(448);
    cpelement_group_966 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(964) & cp_elements(965));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(966),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_895_req_4063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(966), ack => phi_stmt_895_req_0); -- 
    cp_elements(967) <= OrReduce(cp_elements(962) & cp_elements(966));
    cp_elements(968) <= cp_elements(967);
    phi_stmt_895_ack_4068_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_895_ack_0, ack => cp_elements(969)); -- 
    cp_elements(970) <= false;
    cp_elements(971) <= cp_elements(970);
    cp_elements(972) <= false;
    cp_elements(973) <= cp_elements(972);
    cp_elements(974) <= false;
    cp_elements(975) <= cp_elements(974);
    cp_elements(976) <= OrReduce(cp_elements(16) & cp_elements(885));
    cp_elements(977) <= cp_elements(976);
    cp_elements(978) <= OrReduce(cp_elements(156) & cp_elements(228) & cp_elements(257) & cp_elements(295) & cp_elements(495) & cp_elements(883) & cp_elements(896));
    cp_elements(979) <= cp_elements(978);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1024_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1024_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1024_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1024_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1033_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1033_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1033_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1048_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1063_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1063_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1063_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1078_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1078_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1078_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_549_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_558_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_565_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_794_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_794_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_794_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_794_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_843_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_843_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_843_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_843_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_961_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_961_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_961_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_975_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_975_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_975_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_975_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_982_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_982_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_982_root_address : std_logic_vector(15 downto 0);
    signal binary_610_wire : std_logic_vector(31 downto 0);
    signal binary_656_wire : std_logic_vector(31 downto 0);
    signal binary_690_wire : std_logic_vector(31 downto 0);
    signal binary_728_wire : std_logic_vector(31 downto 0);
    signal binary_951_wire : std_logic_vector(31 downto 0);
    signal elt5x_xi11_1038 : std_logic_vector(31 downto 0);
    signal elt5x_xi_1068 : std_logic_vector(31 downto 0);
    signal expr_609_wire_constant : std_logic_vector(31 downto 0);
    signal expr_655_wire_constant : std_logic_vector(31 downto 0);
    signal expr_689_wire_constant : std_logic_vector(31 downto 0);
    signal expr_727_wire_constant : std_logic_vector(31 downto 0);
    signal expr_950_wire_constant : std_logic_vector(31 downto 0);
    signal indvarx_xi12x_xi_754 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xi14x_xi_827 : std_logic_vector(31 downto 0);
    signal orx_xcondx_xi_716 : std_logic_vector(0 downto 0);
    signal ptr_deref_1027_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1027_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1027_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1027_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1027_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1027_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1027_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1041_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1041_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1041_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1041_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1041_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1055_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1055_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1055_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1055_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1055_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1055_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1071_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1071_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1071_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1071_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1071_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1085_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1085_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1085_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1085_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1085_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1085_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_553_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_553_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_553_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_569_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_569_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_569_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_621_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_621_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_621_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_621_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_621_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_621_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_803_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_803_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_803_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_803_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_803_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_803_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_803_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_803_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_882_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_882_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_882_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_882_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_882_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_964_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_964_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_964_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_964_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_964_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_964_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_964_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_964_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_985_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_985_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_985_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_985_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_985_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_985_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_985_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_985_word_offset_3 : std_logic_vector(15 downto 0);
    signal scevgep12x_xix_xi_800 : std_logic_vector(31 downto 0);
    signal scevgep14x_xix_xi_844 : std_logic_vector(31 downto 0);
    signal scevgep_795 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1023_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1023_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_537_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_793_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_793_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_842_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_842_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_974_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_974_scaled : std_logic_vector(15 downto 0);
    signal tmp13_539 : std_logic_vector(31 downto 0);
    signal tmp14_543 : std_logic_vector(31 downto 0);
    signal tmp15_550 : std_logic_vector(31 downto 0);
    signal tmp16_554 : std_logic_vector(31 downto 0);
    signal tmp17_559 : std_logic_vector(31 downto 0);
    signal tmp17x_xix_xi_779 : std_logic_vector(31 downto 0);
    signal tmp18_566 : std_logic_vector(31 downto 0);
    signal tmp19_570 : std_logic_vector(31 downto 0);
    signal tmp20_574 : std_logic_vector(31 downto 0);
    signal tmp21_578 : std_logic_vector(31 downto 0);
    signal tmp22_583 : std_logic_vector(31 downto 0);
    signal tmp23_589 : std_logic_vector(31 downto 0);
    signal tmp24_598 : std_logic_vector(0 downto 0);
    signal tmp25_618 : std_logic_vector(31 downto 0);
    signal tmp26_622 : std_logic_vector(31 downto 0);
    signal tmp27_628 : std_logic_vector(31 downto 0);
    signal tmp28_634 : std_logic_vector(0 downto 0);
    signal tmp29_666 : std_logic_vector(31 downto 0);
    signal tmp30_672 : std_logic_vector(31 downto 0);
    signal tmp31_678 : std_logic_vector(0 downto 0);
    signal tmp32_697 : std_logic_vector(15 downto 0);
    signal tmp33_701 : std_logic_vector(31 downto 0);
    signal tmp34_706 : std_logic_vector(0 downto 0);
    signal tmp34x_xi_640 : std_logic_vector(31 downto 0);
    signal tmp35_711 : std_logic_vector(0 downto 0);
    signal tmp35x_xi_644 : std_logic_vector(15 downto 0);
    signal tmp36_738 : std_logic_vector(0 downto 0);
    signal tmp37_761 : std_logic_vector(31 downto 0);
    signal tmp38_804 : std_logic_vector(15 downto 0);
    signal tmp39_808 : std_logic_vector(31 downto 0);
    signal tmp40_813 : std_logic_vector(31 downto 0);
    signal tmp41_821 : std_logic_vector(0 downto 0);
    signal tmp42_872 : std_logic_vector(0 downto 0);
    signal tmp43_883 : std_logic_vector(7 downto 0);
    signal tmp44_887 : std_logic_vector(31 downto 0);
    signal tmp45_892 : std_logic_vector(31 downto 0);
    signal tmp46_895 : std_logic_vector(31 downto 0);
    signal tmp47_907 : std_logic_vector(31 downto 0);
    signal tmp48_913 : std_logic_vector(31 downto 0);
    signal tmp49_918 : std_logic_vector(31 downto 0);
    signal tmp50_924 : std_logic_vector(31 downto 0);
    signal tmp51_929 : std_logic_vector(31 downto 0);
    signal tmp52_933 : std_logic_vector(15 downto 0);
    signal tmp53_939 : std_logic_vector(0 downto 0);
    signal tmp54_962 : std_logic_vector(31 downto 0);
    signal tmp55_976 : std_logic_vector(31 downto 0);
    signal tmp56_983 : std_logic_vector(31 downto 0);
    signal tmp57_992 : std_logic_vector(0 downto 0);
    signal tmp58_1004 : std_logic_vector(31 downto 0);
    signal tmp59_1009 : std_logic_vector(0 downto 0);
    signal tmp5_751 : std_logic_vector(31 downto 0);
    signal tmp60_1015 : std_logic_vector(31 downto 0);
    signal tmp61_1021 : std_logic_vector(31 downto 0);
    signal tmp62_1025 : std_logic_vector(31 downto 0);
    signal tmp63_1034 : std_logic_vector(31 downto 0);
    signal tmp64_1049 : std_logic_vector(31 downto 0);
    signal tmp65_1053 : std_logic_vector(31 downto 0);
    signal tmp66_1064 : std_logic_vector(31 downto 0);
    signal tmp67_1079 : std_logic_vector(31 downto 0);
    signal tmp68_1083 : std_logic_vector(31 downto 0);
    signal tmp69_1093 : std_logic_vector(0 downto 0);
    signal tmp70_1104 : std_logic_vector(31 downto 0);
    signal tmp8_791 : std_logic_vector(31 downto 0);
    signal tmp_774 : std_logic_vector(31 downto 0);
    signal tmpx_xix_xi_785 : std_logic_vector(31 downto 0);
    signal type_cast_1018_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1091_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1107_wire : std_logic_vector(31 downto 0);
    signal type_cast_587_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_593_wire : std_logic_vector(31 downto 0);
    signal type_cast_596_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_626_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_632_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_638_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_664_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_670_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_676_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_736_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_749_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_758_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_760_wire : std_logic_vector(31 downto 0);
    signal type_cast_765_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_767_wire : std_logic_vector(31 downto 0);
    signal type_cast_772_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_783_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_789_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_816_wire : std_logic_vector(31 downto 0);
    signal type_cast_819_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_825_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_838_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_850_wire : std_logic_vector(31 downto 0);
    signal type_cast_853_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_857_wire : std_logic_vector(31 downto 0);
    signal type_cast_859_wire : std_logic_vector(31 downto 0);
    signal type_cast_863_wire : std_logic_vector(31 downto 0);
    signal type_cast_865_wire : std_logic_vector(31 downto 0);
    signal type_cast_870_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_898_wire : std_logic_vector(31 downto 0);
    signal type_cast_900_wire : std_logic_vector(31 downto 0);
    signal type_cast_905_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_911_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_937_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_970_wire_constant : std_logic_vector(31 downto 0);
    signal val6x_xi12_1042 : std_logic_vector(31 downto 0);
    signal val6x_xi_1072 : std_logic_vector(31 downto 0);
    signal xx_xinx_xlcssax_xix_xi_854 : std_logic_vector(31 downto 0);
    signal xx_xlcssa5x_xix_xi_847 : std_logic_vector(31 downto 0);
    signal xx_xlcssax_xix_xi_860 : std_logic_vector(31 downto 0);
    signal xx_xsum20x_xi_840 : std_logic_vector(31 downto 0);
    signal xx_xsumx_xi_972 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1024_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1033_final_offset <= "0000000000011110";
    array_obj_ref_1048_final_offset <= "0000000000011100";
    array_obj_ref_1063_final_offset <= "0000000000011110";
    array_obj_ref_1078_final_offset <= "0000000000011100";
    array_obj_ref_549_final_offset <= "0000000000001100";
    array_obj_ref_558_final_offset <= "0000000000001110";
    array_obj_ref_565_final_offset <= "0000000000010000";
    array_obj_ref_794_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_843_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_961_final_offset <= "0000000001010000";
    array_obj_ref_975_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_982_final_offset <= "0000000001010100";
    expr_609_wire_constant <= "11111111111111111111100000000000";
    expr_655_wire_constant <= "11111111111111111111100000000000";
    expr_689_wire_constant <= "11111111111111111111100000000000";
    expr_727_wire_constant <= "11111111111111111111100000000000";
    expr_950_wire_constant <= "11111111111111111111100000000000";
    ptr_deref_1027_word_offset_0 <= "0000000000000000";
    ptr_deref_1027_word_offset_1 <= "0000000000000001";
    ptr_deref_1027_word_offset_2 <= "0000000000000010";
    ptr_deref_1027_word_offset_3 <= "0000000000000011";
    ptr_deref_1041_word_offset_0 <= "0000000000000000";
    ptr_deref_1041_word_offset_1 <= "0000000000000001";
    ptr_deref_1041_word_offset_2 <= "0000000000000010";
    ptr_deref_1041_word_offset_3 <= "0000000000000011";
    ptr_deref_1055_word_offset_0 <= "0000000000000000";
    ptr_deref_1055_word_offset_1 <= "0000000000000001";
    ptr_deref_1055_word_offset_2 <= "0000000000000010";
    ptr_deref_1055_word_offset_3 <= "0000000000000011";
    ptr_deref_1071_word_offset_0 <= "0000000000000000";
    ptr_deref_1071_word_offset_1 <= "0000000000000001";
    ptr_deref_1071_word_offset_2 <= "0000000000000010";
    ptr_deref_1071_word_offset_3 <= "0000000000000011";
    ptr_deref_1085_word_offset_0 <= "0000000000000000";
    ptr_deref_1085_word_offset_1 <= "0000000000000001";
    ptr_deref_1085_word_offset_2 <= "0000000000000010";
    ptr_deref_1085_word_offset_3 <= "0000000000000011";
    ptr_deref_553_word_offset_0 <= "0000000000000000";
    ptr_deref_553_word_offset_1 <= "0000000000000001";
    ptr_deref_553_word_offset_2 <= "0000000000000010";
    ptr_deref_553_word_offset_3 <= "0000000000000011";
    ptr_deref_569_word_offset_0 <= "0000000000000000";
    ptr_deref_569_word_offset_1 <= "0000000000000001";
    ptr_deref_569_word_offset_2 <= "0000000000000010";
    ptr_deref_569_word_offset_3 <= "0000000000000011";
    ptr_deref_621_word_offset_0 <= "0000000000000000";
    ptr_deref_621_word_offset_1 <= "0000000000000001";
    ptr_deref_621_word_offset_2 <= "0000000000000010";
    ptr_deref_621_word_offset_3 <= "0000000000000011";
    ptr_deref_803_word_offset_0 <= "0000000000000000";
    ptr_deref_803_word_offset_1 <= "0000000000000001";
    ptr_deref_882_word_offset_0 <= "0000000000000000";
    ptr_deref_964_word_offset_0 <= "0000000000000000";
    ptr_deref_964_word_offset_1 <= "0000000000000001";
    ptr_deref_964_word_offset_2 <= "0000000000000010";
    ptr_deref_964_word_offset_3 <= "0000000000000011";
    ptr_deref_985_word_offset_0 <= "0000000000000000";
    ptr_deref_985_word_offset_1 <= "0000000000000001";
    ptr_deref_985_word_offset_2 <= "0000000000000010";
    ptr_deref_985_word_offset_3 <= "0000000000000011";
    type_cast_1018_wire_constant <= "00000000000000000000000000000000";
    type_cast_1091_wire_constant <= "11111111111111111111111111111111";
    type_cast_587_wire_constant <= "11111111111111111111111111110010";
    type_cast_596_wire_constant <= "00000000000000000000000000010100";
    type_cast_626_wire_constant <= "00000000000000000000000011110000";
    type_cast_632_wire_constant <= "00000000000000000000000001000000";
    type_cast_638_wire_constant <= "00000000000000000000000000010000";
    type_cast_664_wire_constant <= "00000000000000000000000000000010";
    type_cast_670_wire_constant <= "00000000000000000000000000111100";
    type_cast_676_wire_constant <= "00000000000000000000000000010100";
    type_cast_736_wire_constant <= "00000000000000000000000000000001";
    type_cast_749_wire_constant <= "11111111111111111111111111111110";
    type_cast_758_wire_constant <= "00000000000000000000000000000000";
    type_cast_765_wire_constant <= "00000000000000000000000000000000";
    type_cast_772_wire_constant <= "11111111111111111111111111111110";
    type_cast_783_wire_constant <= "00000000000000000000000000000001";
    type_cast_789_wire_constant <= "00000000000000000000000000001110";
    type_cast_819_wire_constant <= "00000000000000000000000000000001";
    type_cast_825_wire_constant <= "00000000000000000000000000000001";
    type_cast_838_wire_constant <= "00000000000000000000000000010000";
    type_cast_853_wire_constant <= "00000000000000000000000000000000";
    type_cast_870_wire_constant <= "00000000000000000000000000000001";
    type_cast_905_wire_constant <= "00000000000000001111111111111111";
    type_cast_911_wire_constant <= "00000000000000000000000000010000";
    type_cast_922_wire_constant <= "00000000000000000000000000010000";
    type_cast_937_wire_constant <= "1111111111111111";
    type_cast_970_wire_constant <= "00000000000000000000000000001110";
    phi_stmt_754: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_758_wire_constant & type_cast_760_wire;
      req <= phi_stmt_754_req_0 & phi_stmt_754_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_754_ack_0,
          idata => idata,
          odata => indvarx_xi12x_xi_754,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_754
    phi_stmt_761: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_765_wire_constant & type_cast_767_wire;
      req <= phi_stmt_761_req_0 & phi_stmt_761_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_761_ack_0,
          idata => idata,
          odata => tmp37_761,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_761
    phi_stmt_847: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_850_wire & type_cast_853_wire_constant;
      req <= phi_stmt_847_req_0 & phi_stmt_847_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_847_ack_0,
          idata => idata,
          odata => xx_xlcssa5x_xix_xi_847,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_847
    phi_stmt_854: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_857_wire & type_cast_859_wire;
      req <= phi_stmt_854_req_0 & phi_stmt_854_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_854_ack_0,
          idata => idata,
          odata => xx_xinx_xlcssax_xix_xi_854,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_854
    phi_stmt_860: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_863_wire & type_cast_865_wire;
      req <= phi_stmt_860_req_0 & phi_stmt_860_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_860_ack_0,
          idata => idata,
          odata => xx_xlcssax_xix_xi_860,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_860
    phi_stmt_895: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_898_wire & type_cast_900_wire;
      req <= phi_stmt_895_req_0 & phi_stmt_895_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_895_ack_0,
          idata => idata,
          odata => tmp46_895,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_895
    ternary_1014_inst: SelectBase generic map(data_width => 32) -- 
      port map( x => tmp22_583, y => tmp58_1004, sel => tmp59_1009, z => tmp60_1015, req => ternary_1014_inst_req_0, ack => ternary_1014_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1024_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp19_570, dout => array_obj_ref_1024_resized_base_address, req => array_obj_ref_1024_base_resize_req_0, ack => array_obj_ref_1024_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1024_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1024_root_address, dout => tmp62_1025, req => array_obj_ref_1024_final_reg_req_0, ack => array_obj_ref_1024_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1024_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp61_1021, dout => simple_obj_ref_1023_resized, req => array_obj_ref_1024_index_0_resize_req_0, ack => array_obj_ref_1024_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1024_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1023_scaled, dout => array_obj_ref_1024_final_offset, req => array_obj_ref_1024_offset_inst_req_0, ack => array_obj_ref_1024_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1033_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_1033_resized_base_address, req => array_obj_ref_1033_base_resize_req_0, ack => array_obj_ref_1033_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1033_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1033_root_address, dout => tmp63_1034, req => array_obj_ref_1033_final_reg_req_0, ack => array_obj_ref_1033_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1048_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_1048_resized_base_address, req => array_obj_ref_1048_base_resize_req_0, ack => array_obj_ref_1048_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1048_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1048_root_address, dout => tmp64_1049, req => array_obj_ref_1048_final_reg_req_0, ack => array_obj_ref_1048_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1063_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_1063_resized_base_address, req => array_obj_ref_1063_base_resize_req_0, ack => array_obj_ref_1063_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1063_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1063_root_address, dout => tmp66_1064, req => array_obj_ref_1063_final_reg_req_0, ack => array_obj_ref_1063_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1078_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_1078_resized_base_address, req => array_obj_ref_1078_base_resize_req_0, ack => array_obj_ref_1078_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1078_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1078_root_address, dout => tmp67_1079, req => array_obj_ref_1078_final_reg_req_0, ack => array_obj_ref_1078_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_549_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_549_resized_base_address, req => array_obj_ref_549_base_resize_req_0, ack => array_obj_ref_549_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_549_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_549_root_address, dout => tmp15_550, req => array_obj_ref_549_final_reg_req_0, ack => array_obj_ref_549_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_558_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_558_resized_base_address, req => array_obj_ref_558_base_resize_req_0, ack => array_obj_ref_558_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_558_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_558_root_address, dout => tmp17_559, req => array_obj_ref_558_final_reg_req_0, ack => array_obj_ref_558_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_565_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_565_resized_base_address, req => array_obj_ref_565_base_resize_req_0, ack => array_obj_ref_565_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_565_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_565_root_address, dout => tmp18_566, req => array_obj_ref_565_final_reg_req_0, ack => array_obj_ref_565_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_794_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_794_resized_base_address, req => array_obj_ref_794_base_resize_req_0, ack => array_obj_ref_794_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_794_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_794_root_address, dout => scevgep_795, req => array_obj_ref_794_final_reg_req_0, ack => array_obj_ref_794_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_794_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_791, dout => simple_obj_ref_793_resized, req => array_obj_ref_794_index_0_resize_req_0, ack => array_obj_ref_794_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_794_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_793_scaled, dout => array_obj_ref_794_final_offset, req => array_obj_ref_794_offset_inst_req_0, ack => array_obj_ref_794_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_843_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_843_resized_base_address, req => array_obj_ref_843_base_resize_req_0, ack => array_obj_ref_843_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_843_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_843_root_address, dout => scevgep14x_xix_xi_844, req => array_obj_ref_843_final_reg_req_0, ack => array_obj_ref_843_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_843_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsum20x_xi_840, dout => simple_obj_ref_842_resized, req => array_obj_ref_843_index_0_resize_req_0, ack => array_obj_ref_843_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_843_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_842_scaled, dout => array_obj_ref_843_final_offset, req => array_obj_ref_843_offset_inst_req_0, ack => array_obj_ref_843_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_961_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_961_resized_base_address, req => array_obj_ref_961_base_resize_req_0, ack => array_obj_ref_961_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_961_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_961_root_address, dout => tmp54_962, req => array_obj_ref_961_final_reg_req_0, ack => array_obj_ref_961_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_975_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_554, dout => array_obj_ref_975_resized_base_address, req => array_obj_ref_975_base_resize_req_0, ack => array_obj_ref_975_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_975_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_975_root_address, dout => tmp55_976, req => array_obj_ref_975_final_reg_req_0, ack => array_obj_ref_975_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_975_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsumx_xi_972, dout => simple_obj_ref_974_resized, req => array_obj_ref_975_index_0_resize_req_0, ack => array_obj_ref_975_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_975_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_974_scaled, dout => array_obj_ref_975_final_offset, req => array_obj_ref_975_offset_inst_req_0, ack => array_obj_ref_975_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_982_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_543, dout => array_obj_ref_982_resized_base_address, req => array_obj_ref_982_base_resize_req_0, ack => array_obj_ref_982_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_982_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_982_root_address, dout => tmp56_983, req => array_obj_ref_982_final_reg_req_0, ack => array_obj_ref_982_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1027_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_566, dout => ptr_deref_1027_resized_base_address, req => ptr_deref_1027_base_resize_req_0, ack => ptr_deref_1027_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1041_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi11_1038, dout => ptr_deref_1041_resized_base_address, req => ptr_deref_1041_base_resize_req_0, ack => ptr_deref_1041_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1055_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp65_1053, dout => ptr_deref_1055_resized_base_address, req => ptr_deref_1055_base_resize_req_0, ack => ptr_deref_1055_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1071_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi_1068, dout => ptr_deref_1071_resized_base_address, req => ptr_deref_1071_base_resize_req_0, ack => ptr_deref_1071_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1085_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp68_1083, dout => ptr_deref_1085_resized_base_address, req => ptr_deref_1085_base_resize_req_0, ack => ptr_deref_1085_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_553_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp15_550, dout => ptr_deref_553_resized_base_address, req => ptr_deref_553_base_resize_req_0, ack => ptr_deref_553_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_569_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_566, dout => ptr_deref_569_resized_base_address, req => ptr_deref_569_base_resize_req_0, ack => ptr_deref_569_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_621_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp25_618, dout => ptr_deref_621_resized_base_address, req => ptr_deref_621_base_resize_req_0, ack => ptr_deref_621_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_803_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => scevgep12x_xix_xi_800, dout => ptr_deref_803_resized_base_address, req => ptr_deref_803_base_resize_req_0, ack => ptr_deref_803_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_882_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xinx_xlcssax_xix_xi_854, dout => ptr_deref_882_resized_base_address, req => ptr_deref_882_base_resize_req_0, ack => ptr_deref_882_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_964_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp54_962, dout => ptr_deref_964_resized_base_address, req => ptr_deref_964_base_resize_req_0, ack => ptr_deref_964_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_985_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp56_983, dout => ptr_deref_985_resized_base_address, req => ptr_deref_985_base_resize_req_0, ack => ptr_deref_985_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1037_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp63_1034, dout => elt5x_xi11_1038, req => type_cast_1037_inst_req_0, ack => type_cast_1037_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1052_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp64_1049, dout => tmp65_1053, req => type_cast_1052_inst_req_0, ack => type_cast_1052_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1067_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp66_1064, dout => elt5x_xi_1068, req => type_cast_1067_inst_req_0, ack => type_cast_1067_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1082_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp67_1079, dout => tmp68_1083, req => type_cast_1082_inst_req_0, ack => type_cast_1082_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1103_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp14_543, dout => tmp70_1104, req => type_cast_1103_inst_req_0, ack => type_cast_1103_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1107_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp70_1104, dout => type_cast_1107_wire, req => type_cast_1107_inst_req_0, ack => type_cast_1107_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_538_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_537_wire, dout => tmp13_539, req => type_cast_538_inst_req_0, ack => type_cast_538_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_542_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_539, dout => tmp14_543, req => type_cast_542_inst_req_0, ack => type_cast_542_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_573_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp19_570, dout => tmp20_574, req => type_cast_573_inst_req_0, ack => type_cast_573_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_577_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp16_554, dout => tmp21_578, req => type_cast_577_inst_req_0, ack => type_cast_577_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_593_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp23_589, dout => type_cast_593_wire, req => type_cast_593_inst_req_0, ack => type_cast_593_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_617_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_559, dout => tmp25_618, req => type_cast_617_inst_req_0, ack => type_cast_617_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_643_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp34x_xi_640, dout => tmp35x_xi_644, req => type_cast_643_inst_req_0, ack => type_cast_643_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_700_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp32_697, dout => tmp33_701, req => type_cast_700_inst_req_0, ack => type_cast_700_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_760_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnextx_xi14x_xi_827, dout => type_cast_760_wire, req => type_cast_760_inst_req_0, ack => type_cast_760_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_767_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_813, dout => type_cast_767_wire, req => type_cast_767_inst_req_0, ack => type_cast_767_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_799_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => scevgep_795, dout => scevgep12x_xix_xi_800, req => type_cast_799_inst_req_0, ack => type_cast_799_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_807_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp38_804, dout => tmp39_808, req => type_cast_807_inst_req_0, ack => type_cast_807_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_816_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_779, dout => type_cast_816_wire, req => type_cast_816_inst_req_0, ack => type_cast_816_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_850_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_813, dout => type_cast_850_wire, req => type_cast_850_inst_req_0, ack => type_cast_850_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_857_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => scevgep14x_xix_xi_844, dout => type_cast_857_wire, req => type_cast_857_inst_req_0, ack => type_cast_857_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_859_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17_559, dout => type_cast_859_wire, req => type_cast_859_inst_req_0, ack => type_cast_859_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_863_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_779, dout => type_cast_863_wire, req => type_cast_863_inst_req_0, ack => type_cast_863_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_865_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp30_672, dout => type_cast_865_wire, req => type_cast_865_inst_req_0, ack => type_cast_865_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_886_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp43_883, dout => tmp44_887, req => type_cast_886_inst_req_0, ack => type_cast_886_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_898_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp45_892, dout => type_cast_898_wire, req => type_cast_898_inst_req_0, ack => type_cast_898_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_900_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => xx_xlcssa5x_xix_xi_847, dout => type_cast_900_wire, req => type_cast_900_inst_req_0, ack => type_cast_900_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_932_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp51_929, dout => tmp52_933, req => type_cast_932_inst_req_0, ack => type_cast_932_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1024_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1024_index_0_rename_ack_0 <= array_obj_ref_1024_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1023_resized;
      simple_obj_ref_1023_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_794_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_794_index_0_rename_ack_0 <= array_obj_ref_794_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_793_resized;
      simple_obj_ref_793_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_843_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_843_index_0_rename_ack_0 <= array_obj_ref_843_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_842_resized;
      simple_obj_ref_842_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_975_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_975_index_0_rename_ack_0 <= array_obj_ref_975_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_974_resized;
      simple_obj_ref_974_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1027_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1027_gather_scatter_ack_0 <= ptr_deref_1027_gather_scatter_req_0;
      aggregated_sig <= tmp62_1025;
      ptr_deref_1027_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1027_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1027_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1027_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1027_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1027_root_address_inst_ack_0 <= ptr_deref_1027_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1027_resized_base_address;
      ptr_deref_1027_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1041_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1041_gather_scatter_ack_0 <= ptr_deref_1041_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1041_data_3 & ptr_deref_1041_data_2 & ptr_deref_1041_data_1 & ptr_deref_1041_data_0;
      val6x_xi12_1042 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1041_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1041_root_address_inst_ack_0 <= ptr_deref_1041_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1041_resized_base_address;
      ptr_deref_1041_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1055_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1055_gather_scatter_ack_0 <= ptr_deref_1055_gather_scatter_req_0;
      aggregated_sig <= val6x_xi12_1042;
      ptr_deref_1055_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1055_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1055_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1055_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1055_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1055_root_address_inst_ack_0 <= ptr_deref_1055_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1055_resized_base_address;
      ptr_deref_1055_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1071_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1071_gather_scatter_ack_0 <= ptr_deref_1071_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1071_data_3 & ptr_deref_1071_data_2 & ptr_deref_1071_data_1 & ptr_deref_1071_data_0;
      val6x_xi_1072 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1071_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1071_root_address_inst_ack_0 <= ptr_deref_1071_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1071_resized_base_address;
      ptr_deref_1071_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1085_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1085_gather_scatter_ack_0 <= ptr_deref_1085_gather_scatter_req_0;
      aggregated_sig <= val6x_xi_1072;
      ptr_deref_1085_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1085_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1085_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1085_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1085_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1085_root_address_inst_ack_0 <= ptr_deref_1085_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1085_resized_base_address;
      ptr_deref_1085_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_553_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_553_gather_scatter_ack_0 <= ptr_deref_553_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_553_data_3 & ptr_deref_553_data_2 & ptr_deref_553_data_1 & ptr_deref_553_data_0;
      tmp16_554 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_553_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_553_root_address_inst_ack_0 <= ptr_deref_553_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_553_resized_base_address;
      ptr_deref_553_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_569_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_569_gather_scatter_ack_0 <= ptr_deref_569_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_569_data_3 & ptr_deref_569_data_2 & ptr_deref_569_data_1 & ptr_deref_569_data_0;
      tmp19_570 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_569_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_569_root_address_inst_ack_0 <= ptr_deref_569_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_569_resized_base_address;
      ptr_deref_569_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_621_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_621_gather_scatter_ack_0 <= ptr_deref_621_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_621_data_3 & ptr_deref_621_data_2 & ptr_deref_621_data_1 & ptr_deref_621_data_0;
      tmp26_622 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_621_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_621_root_address_inst_ack_0 <= ptr_deref_621_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_621_resized_base_address;
      ptr_deref_621_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_803_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_803_gather_scatter_ack_0 <= ptr_deref_803_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_803_data_1 & ptr_deref_803_data_0;
      tmp38_804 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_803_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_803_root_address_inst_ack_0 <= ptr_deref_803_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_803_resized_base_address;
      ptr_deref_803_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_882_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_882_addr_0_ack_0 <= ptr_deref_882_addr_0_req_0;
      aggregated_sig <= ptr_deref_882_root_address;
      ptr_deref_882_word_address_0 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_882_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_882_gather_scatter_ack_0 <= ptr_deref_882_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_882_data_0;
      tmp43_883 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_882_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_882_root_address_inst_ack_0 <= ptr_deref_882_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_882_resized_base_address;
      ptr_deref_882_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_964_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_964_gather_scatter_ack_0 <= ptr_deref_964_gather_scatter_req_0;
      aggregated_sig <= tmp17_559;
      ptr_deref_964_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_964_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_964_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_964_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_964_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_964_root_address_inst_ack_0 <= ptr_deref_964_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_964_resized_base_address;
      ptr_deref_964_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_985_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_985_gather_scatter_ack_0 <= ptr_deref_985_gather_scatter_req_0;
      aggregated_sig <= tmp55_976;
      ptr_deref_985_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_985_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_985_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_985_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_985_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_985_root_address_inst_ack_0 <= ptr_deref_985_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_985_resized_base_address;
      ptr_deref_985_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_1094_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp69_1093;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1094_branch_req_0,
          ack0 => if_stmt_1094_branch_ack_0,
          ack1 => if_stmt_1094_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_599_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp24_598;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_599_branch_req_0,
          ack0 => if_stmt_599_branch_ack_0,
          ack1 => if_stmt_599_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_645_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp28_634;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_645_branch_req_0,
          ack0 => if_stmt_645_branch_ack_0,
          ack1 => if_stmt_645_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_679_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp31_678;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_679_branch_req_0,
          ack0 => if_stmt_679_branch_ack_0,
          ack1 => if_stmt_679_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_717_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xi_716;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_717_branch_req_0,
          ack0 => if_stmt_717_branch_ack_0,
          ack1 => if_stmt_717_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_739_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_738;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_739_branch_req_0,
          ack0 => if_stmt_739_branch_ack_0,
          ack1 => if_stmt_739_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_828_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp41_821;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_828_branch_req_0,
          ack0 => if_stmt_828_branch_ack_0,
          ack1 => if_stmt_828_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_873_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp42_872;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_873_branch_req_0,
          ack0 => if_stmt_873_branch_ack_0,
          ack1 => if_stmt_873_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_940_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp53_939;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_940_branch_req_0,
          ack0 => if_stmt_940_branch_ack_0,
          ack1 => if_stmt_940_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_993_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp57_992;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_993_branch_req_0,
          ack0 => if_stmt_993_branch_ack_0,
          ack1 => if_stmt_993_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1024_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1024_final_offset & array_obj_ref_1024_resized_base_address;
      array_obj_ref_1024_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1024_root_address_inst_req_0,
          ackL => array_obj_ref_1024_root_address_inst_ack_0,
          reqR => array_obj_ref_1024_root_address_inst_req_1,
          ackR => array_obj_ref_1024_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1033_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1033_resized_base_address;
      array_obj_ref_1033_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1033_root_address_inst_req_0,
          ackL => array_obj_ref_1033_root_address_inst_ack_0,
          reqR => array_obj_ref_1033_root_address_inst_req_1,
          ackR => array_obj_ref_1033_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1048_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1048_resized_base_address;
      array_obj_ref_1048_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1048_root_address_inst_req_0,
          ackL => array_obj_ref_1048_root_address_inst_ack_0,
          reqR => array_obj_ref_1048_root_address_inst_req_1,
          ackR => array_obj_ref_1048_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1063_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1063_resized_base_address;
      array_obj_ref_1063_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1063_root_address_inst_req_0,
          ackL => array_obj_ref_1063_root_address_inst_ack_0,
          reqR => array_obj_ref_1063_root_address_inst_req_1,
          ackR => array_obj_ref_1063_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1078_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1078_resized_base_address;
      array_obj_ref_1078_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1078_root_address_inst_req_0,
          ackL => array_obj_ref_1078_root_address_inst_ack_0,
          reqR => array_obj_ref_1078_root_address_inst_req_1,
          ackR => array_obj_ref_1078_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_549_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_549_resized_base_address;
      array_obj_ref_549_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_549_root_address_inst_req_0,
          ackL => array_obj_ref_549_root_address_inst_ack_0,
          reqR => array_obj_ref_549_root_address_inst_req_1,
          ackR => array_obj_ref_549_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_558_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_558_resized_base_address;
      array_obj_ref_558_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_558_root_address_inst_req_0,
          ackL => array_obj_ref_558_root_address_inst_ack_0,
          reqR => array_obj_ref_558_root_address_inst_req_1,
          ackR => array_obj_ref_558_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_565_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_565_resized_base_address;
      array_obj_ref_565_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_565_root_address_inst_req_0,
          ackL => array_obj_ref_565_root_address_inst_ack_0,
          reqR => array_obj_ref_565_root_address_inst_req_1,
          ackR => array_obj_ref_565_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_794_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_794_final_offset & array_obj_ref_794_resized_base_address;
      array_obj_ref_794_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_794_root_address_inst_req_0,
          ackL => array_obj_ref_794_root_address_inst_ack_0,
          reqR => array_obj_ref_794_root_address_inst_req_1,
          ackR => array_obj_ref_794_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_843_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_843_final_offset & array_obj_ref_843_resized_base_address;
      array_obj_ref_843_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_843_root_address_inst_req_0,
          ackL => array_obj_ref_843_root_address_inst_ack_0,
          reqR => array_obj_ref_843_root_address_inst_req_1,
          ackR => array_obj_ref_843_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_961_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_961_resized_base_address;
      array_obj_ref_961_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_961_root_address_inst_req_0,
          ackL => array_obj_ref_961_root_address_inst_ack_0,
          reqR => array_obj_ref_961_root_address_inst_req_1,
          ackR => array_obj_ref_961_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_975_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_975_final_offset & array_obj_ref_975_resized_base_address;
      array_obj_ref_975_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_975_root_address_inst_req_0,
          ackL => array_obj_ref_975_root_address_inst_ack_0,
          reqR => array_obj_ref_975_root_address_inst_req_1,
          ackR => array_obj_ref_975_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_982_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_982_resized_base_address;
      array_obj_ref_982_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_982_root_address_inst_req_0,
          ackL => array_obj_ref_982_root_address_inst_ack_0,
          reqR => array_obj_ref_982_root_address_inst_req_1,
          ackR => array_obj_ref_982_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_1003_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp23_589 & tmp33_701;
      tmp58_1004 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1003_inst_req_0,
          ackL => binary_1003_inst_ack_0,
          reqR => binary_1003_inst_req_1,
          ackR => binary_1003_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_710_inst binary_1008_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_701 & tmp30_672 & tmp22_583 & tmp58_1004;
      tmp35_711 <= data_out(1 downto 1);
      tmp59_1009 <= data_out(0 downto 0);
      reqL(1) <= binary_710_inst_req_0;
      reqL(0) <= binary_1008_inst_req_0;
      binary_710_inst_ack_0 <= ackL(1);
      binary_1008_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_710_inst_req_1;
      reqR(0) <= binary_1008_inst_req_1;
      binary_710_inst_ack_1 <= ackR(1);
      binary_1008_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1020_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1018_wire_constant & tmp60_1015;
      tmp61_1021 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1020_inst_req_0,
          ackL => binary_1020_inst_ack_0,
          reqR => binary_1020_inst_req_1,
          ackR => binary_1020_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1092_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp14_543;
      tmp69_1093 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1092_inst_req_0,
          ackL => binary_1092_inst_ack_0,
          reqR => binary_1092_inst_req_1,
          ackR => binary_1092_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_582_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_574 & tmp21_578;
      tmp22_583 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_582_inst_req_0,
          ackL => binary_582_inst_ack_0,
          reqR => binary_582_inst_req_1,
          ackR => binary_582_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_588_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp22_583;
      tmp23_589 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111110010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_588_inst_req_0,
          ackL => binary_588_inst_ack_0,
          reqR => binary_588_inst_req_1,
          ackR => binary_588_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_597_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_593_wire;
      tmp24_598 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_597_inst_req_0,
          ackL => binary_597_inst_ack_0,
          reqR => binary_597_inst_req_1,
          ackR => binary_597_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_610_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_539;
      binary_610_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_610_inst_req_0,
          ackL => binary_610_inst_ack_0,
          reqR => binary_610_inst_req_1,
          ackR => binary_610_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_627_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_622;
      tmp27_628 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011110000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_627_inst_req_0,
          ackL => binary_627_inst_ack_0,
          reqR => binary_627_inst_req_1,
          ackR => binary_627_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_633_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp27_628;
      tmp28_634 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_633_inst_req_0,
          ackL => binary_633_inst_ack_0,
          reqR => binary_633_inst_req_1,
          ackR => binary_633_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_639_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_622;
      tmp34x_xi_640 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_639_inst_req_0,
          ackL => binary_639_inst_ack_0,
          reqR => binary_639_inst_req_1,
          ackR => binary_639_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_656_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_539;
      binary_656_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_656_inst_req_0,
          ackL => binary_656_inst_ack_0,
          reqR => binary_656_inst_req_1,
          ackR => binary_656_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_665_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_622;
      tmp29_666 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_665_inst_req_0,
          ackL => binary_665_inst_ack_0,
          reqR => binary_665_inst_req_1,
          ackR => binary_665_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_671_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp29_666;
      tmp30_672 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000111100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_671_inst_req_0,
          ackL => binary_671_inst_ack_0,
          reqR => binary_671_inst_req_1,
          ackR => binary_671_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_677_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_672;
      tmp31_678 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_677_inst_req_0,
          ackL => binary_677_inst_ack_0,
          reqR => binary_677_inst_req_1,
          ackR => binary_677_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_690_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_539;
      binary_690_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_690_inst_req_0,
          ackL => binary_690_inst_ack_0,
          reqR => binary_690_inst_req_1,
          ackR => binary_690_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_705_inst binary_991_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_701 & tmp23_589 & tmp23_589 & tmp33_701;
      tmp34_706 <= data_out(1 downto 1);
      tmp57_992 <= data_out(0 downto 0);
      reqL(1) <= binary_705_inst_req_0;
      reqL(0) <= binary_991_inst_req_0;
      binary_705_inst_ack_0 <= ackL(1);
      binary_991_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_705_inst_req_1;
      reqR(0) <= binary_991_inst_req_1;
      binary_705_inst_ack_1 <= ackR(1);
      binary_991_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_715_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp34_706 & tmp35_711;
      orx_xcondx_xi_716 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_715_inst_req_0,
          ackL => binary_715_inst_ack_0,
          reqR => binary_715_inst_req_1,
          ackR => binary_715_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_728_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_539;
      binary_728_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_728_inst_req_0,
          ackL => binary_728_inst_ack_0,
          reqR => binary_728_inst_req_1,
          ackR => binary_728_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_737_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_672;
      tmp36_738 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_737_inst_req_0,
          ackL => binary_737_inst_ack_0,
          reqR => binary_737_inst_req_1,
          ackR => binary_737_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_750_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_672;
      tmp5_751 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_750_inst_req_0,
          ackL => binary_750_inst_ack_0,
          reqR => binary_750_inst_req_1,
          ackR => binary_750_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_773_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_754;
      tmp_774 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_773_inst_req_0,
          ackL => binary_773_inst_ack_0,
          reqR => binary_773_inst_req_1,
          ackR => binary_773_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_778_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_751 & tmp_774;
      tmp17x_xix_xi_779 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_778_inst_req_0,
          ackL => binary_778_inst_ack_0,
          reqR => binary_778_inst_req_1,
          ackR => binary_778_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_784_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_754;
      tmpx_xix_xi_785 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_784_inst_req_0,
          ackL => binary_784_inst_ack_0,
          reqR => binary_784_inst_req_1,
          ackR => binary_784_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_790_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_785;
      tmp8_791 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_790_inst_req_0,
          ackL => binary_790_inst_ack_0,
          reqR => binary_790_inst_req_1,
          ackR => binary_790_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_812_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp39_808 & tmp37_761;
      tmp40_813 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_812_inst_req_0,
          ackL => binary_812_inst_ack_0,
          reqR => binary_812_inst_req_1,
          ackR => binary_812_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_820_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_816_wire;
      tmp41_821 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_820_inst_req_0,
          ackL => binary_820_inst_ack_0,
          reqR => binary_820_inst_req_1,
          ackR => binary_820_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_826_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_754;
      indvarx_xnextx_xi14x_xi_827 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_826_inst_req_0,
          ackL => binary_826_inst_ack_0,
          reqR => binary_826_inst_req_1,
          ackR => binary_826_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_839_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_785;
      xx_xsum20x_xi_840 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_839_inst_req_0,
          ackL => binary_839_inst_ack_0,
          reqR => binary_839_inst_req_1,
          ackR => binary_839_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_871_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xlcssax_xix_xi_860;
      tmp42_872 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_871_inst_req_0,
          ackL => binary_871_inst_ack_0,
          reqR => binary_871_inst_req_1,
          ackR => binary_871_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_891_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_887 & xx_xlcssa5x_xix_xi_847;
      tmp45_892 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_891_inst_req_0,
          ackL => binary_891_inst_ack_0,
          reqR => binary_891_inst_req_1,
          ackR => binary_891_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_906_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_895;
      tmp47_907 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_906_inst_req_0,
          ackL => binary_906_inst_ack_0,
          reqR => binary_906_inst_req_1,
          ackR => binary_906_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_912_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_895;
      tmp48_913 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_912_inst_req_0,
          ackL => binary_912_inst_ack_0,
          reqR => binary_912_inst_req_1,
          ackR => binary_912_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_917_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp47_907 & tmp48_913;
      tmp49_918 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_917_inst_req_0,
          ackL => binary_917_inst_ack_0,
          reqR => binary_917_inst_req_1,
          ackR => binary_917_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_923_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_918;
      tmp50_924 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_923_inst_req_0,
          ackL => binary_923_inst_ack_0,
          reqR => binary_923_inst_req_1,
          ackR => binary_923_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_928_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_924 & tmp49_918;
      tmp51_929 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_928_inst_req_0,
          ackL => binary_928_inst_ack_0,
          reqR => binary_928_inst_req_1,
          ackR => binary_928_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_938_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp52_933;
      tmp53_939 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1111111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_938_inst_req_0,
          ackL => binary_938_inst_ack_0,
          reqR => binary_938_inst_req_1,
          ackR => binary_938_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_951_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_539;
      binary_951_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_951_inst_req_0,
          ackL => binary_951_inst_ack_0,
          reqR => binary_951_inst_req_1,
          ackR => binary_951_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_971_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_672;
      xx_xsumx_xi_972 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_971_inst_req_0,
          ackL => binary_971_inst_ack_0,
          reqR => binary_971_inst_req_1,
          ackR => binary_971_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_1027_addr_0 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1027_root_address;
      ptr_deref_1027_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1027_addr_0_req_0,
          ackL => ptr_deref_1027_addr_0_ack_0,
          reqR => ptr_deref_1027_addr_0_req_1,
          ackR => ptr_deref_1027_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_1027_addr_1 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1027_root_address;
      ptr_deref_1027_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1027_addr_1_req_0,
          ackL => ptr_deref_1027_addr_1_ack_0,
          reqR => ptr_deref_1027_addr_1_req_1,
          ackR => ptr_deref_1027_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_1027_addr_2 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1027_root_address;
      ptr_deref_1027_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1027_addr_2_req_0,
          ackL => ptr_deref_1027_addr_2_ack_0,
          reqR => ptr_deref_1027_addr_2_req_1,
          ackR => ptr_deref_1027_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_1027_addr_3 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1027_root_address;
      ptr_deref_1027_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1027_addr_3_req_0,
          ackL => ptr_deref_1027_addr_3_ack_0,
          reqR => ptr_deref_1027_addr_3_req_1,
          ackR => ptr_deref_1027_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_1041_addr_0 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1041_root_address;
      ptr_deref_1041_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1041_addr_0_req_0,
          ackL => ptr_deref_1041_addr_0_ack_0,
          reqR => ptr_deref_1041_addr_0_req_1,
          ackR => ptr_deref_1041_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_1041_addr_1 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1041_root_address;
      ptr_deref_1041_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1041_addr_1_req_0,
          ackL => ptr_deref_1041_addr_1_ack_0,
          reqR => ptr_deref_1041_addr_1_req_1,
          ackR => ptr_deref_1041_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_1041_addr_2 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1041_root_address;
      ptr_deref_1041_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1041_addr_2_req_0,
          ackL => ptr_deref_1041_addr_2_ack_0,
          reqR => ptr_deref_1041_addr_2_req_1,
          ackR => ptr_deref_1041_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_1041_addr_3 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1041_root_address;
      ptr_deref_1041_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1041_addr_3_req_0,
          ackL => ptr_deref_1041_addr_3_ack_0,
          reqR => ptr_deref_1041_addr_3_req_1,
          ackR => ptr_deref_1041_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_1055_addr_0 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1055_root_address;
      ptr_deref_1055_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1055_addr_0_req_0,
          ackL => ptr_deref_1055_addr_0_ack_0,
          reqR => ptr_deref_1055_addr_0_req_1,
          ackR => ptr_deref_1055_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_1055_addr_1 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1055_root_address;
      ptr_deref_1055_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1055_addr_1_req_0,
          ackL => ptr_deref_1055_addr_1_ack_0,
          reqR => ptr_deref_1055_addr_1_req_1,
          ackR => ptr_deref_1055_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_1055_addr_2 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1055_root_address;
      ptr_deref_1055_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1055_addr_2_req_0,
          ackL => ptr_deref_1055_addr_2_ack_0,
          reqR => ptr_deref_1055_addr_2_req_1,
          ackR => ptr_deref_1055_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_1055_addr_3 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1055_root_address;
      ptr_deref_1055_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1055_addr_3_req_0,
          ackL => ptr_deref_1055_addr_3_ack_0,
          reqR => ptr_deref_1055_addr_3_req_1,
          ackR => ptr_deref_1055_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : ptr_deref_1071_addr_0 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1071_root_address;
      ptr_deref_1071_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1071_addr_0_req_0,
          ackL => ptr_deref_1071_addr_0_ack_0,
          reqR => ptr_deref_1071_addr_0_req_1,
          ackR => ptr_deref_1071_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : ptr_deref_1071_addr_1 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1071_root_address;
      ptr_deref_1071_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1071_addr_1_req_0,
          ackL => ptr_deref_1071_addr_1_ack_0,
          reqR => ptr_deref_1071_addr_1_req_1,
          ackR => ptr_deref_1071_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : ptr_deref_1071_addr_2 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1071_root_address;
      ptr_deref_1071_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1071_addr_2_req_0,
          ackL => ptr_deref_1071_addr_2_ack_0,
          reqR => ptr_deref_1071_addr_2_req_1,
          ackR => ptr_deref_1071_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : ptr_deref_1071_addr_3 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1071_root_address;
      ptr_deref_1071_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1071_addr_3_req_0,
          ackL => ptr_deref_1071_addr_3_ack_0,
          reqR => ptr_deref_1071_addr_3_req_1,
          ackR => ptr_deref_1071_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : ptr_deref_1085_addr_0 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1085_root_address;
      ptr_deref_1085_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1085_addr_0_req_0,
          ackL => ptr_deref_1085_addr_0_ack_0,
          reqR => ptr_deref_1085_addr_0_req_1,
          ackR => ptr_deref_1085_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : ptr_deref_1085_addr_1 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1085_root_address;
      ptr_deref_1085_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1085_addr_1_req_0,
          ackL => ptr_deref_1085_addr_1_ack_0,
          reqR => ptr_deref_1085_addr_1_req_1,
          ackR => ptr_deref_1085_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : ptr_deref_1085_addr_2 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1085_root_address;
      ptr_deref_1085_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1085_addr_2_req_0,
          ackL => ptr_deref_1085_addr_2_ack_0,
          reqR => ptr_deref_1085_addr_2_req_1,
          ackR => ptr_deref_1085_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : ptr_deref_1085_addr_3 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1085_root_address;
      ptr_deref_1085_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1085_addr_3_req_0,
          ackL => ptr_deref_1085_addr_3_ack_0,
          reqR => ptr_deref_1085_addr_3_req_1,
          ackR => ptr_deref_1085_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : ptr_deref_553_addr_0 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_0_req_0,
          ackL => ptr_deref_553_addr_0_ack_0,
          reqR => ptr_deref_553_addr_0_req_1,
          ackR => ptr_deref_553_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : ptr_deref_553_addr_1 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_1_req_0,
          ackL => ptr_deref_553_addr_1_ack_0,
          reqR => ptr_deref_553_addr_1_req_1,
          ackR => ptr_deref_553_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : ptr_deref_553_addr_2 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_2_req_0,
          ackL => ptr_deref_553_addr_2_ack_0,
          reqR => ptr_deref_553_addr_2_req_1,
          ackR => ptr_deref_553_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : ptr_deref_553_addr_3 
    SplitOperatorGroup75: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_553_root_address;
      ptr_deref_553_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_553_addr_3_req_0,
          ackL => ptr_deref_553_addr_3_ack_0,
          reqR => ptr_deref_553_addr_3_req_1,
          ackR => ptr_deref_553_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : ptr_deref_569_addr_0 
    SplitOperatorGroup76: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_0_req_0,
          ackL => ptr_deref_569_addr_0_ack_0,
          reqR => ptr_deref_569_addr_0_req_1,
          ackR => ptr_deref_569_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : ptr_deref_569_addr_1 
    SplitOperatorGroup77: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_1_req_0,
          ackL => ptr_deref_569_addr_1_ack_0,
          reqR => ptr_deref_569_addr_1_req_1,
          ackR => ptr_deref_569_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : ptr_deref_569_addr_2 
    SplitOperatorGroup78: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_2_req_0,
          ackL => ptr_deref_569_addr_2_ack_0,
          reqR => ptr_deref_569_addr_2_req_1,
          ackR => ptr_deref_569_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : ptr_deref_569_addr_3 
    SplitOperatorGroup79: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_569_root_address;
      ptr_deref_569_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_569_addr_3_req_0,
          ackL => ptr_deref_569_addr_3_ack_0,
          reqR => ptr_deref_569_addr_3_req_1,
          ackR => ptr_deref_569_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : ptr_deref_621_addr_0 
    SplitOperatorGroup80: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_621_root_address;
      ptr_deref_621_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_621_addr_0_req_0,
          ackL => ptr_deref_621_addr_0_ack_0,
          reqR => ptr_deref_621_addr_0_req_1,
          ackR => ptr_deref_621_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : ptr_deref_621_addr_1 
    SplitOperatorGroup81: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_621_root_address;
      ptr_deref_621_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_621_addr_1_req_0,
          ackL => ptr_deref_621_addr_1_ack_0,
          reqR => ptr_deref_621_addr_1_req_1,
          ackR => ptr_deref_621_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : ptr_deref_621_addr_2 
    SplitOperatorGroup82: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_621_root_address;
      ptr_deref_621_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_621_addr_2_req_0,
          ackL => ptr_deref_621_addr_2_ack_0,
          reqR => ptr_deref_621_addr_2_req_1,
          ackR => ptr_deref_621_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : ptr_deref_621_addr_3 
    SplitOperatorGroup83: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_621_root_address;
      ptr_deref_621_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_621_addr_3_req_0,
          ackL => ptr_deref_621_addr_3_ack_0,
          reqR => ptr_deref_621_addr_3_req_1,
          ackR => ptr_deref_621_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : ptr_deref_803_addr_0 
    SplitOperatorGroup84: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_803_root_address;
      ptr_deref_803_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_803_addr_0_req_0,
          ackL => ptr_deref_803_addr_0_ack_0,
          reqR => ptr_deref_803_addr_0_req_1,
          ackR => ptr_deref_803_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : ptr_deref_803_addr_1 
    SplitOperatorGroup85: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_803_root_address;
      ptr_deref_803_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_803_addr_1_req_0,
          ackL => ptr_deref_803_addr_1_ack_0,
          reqR => ptr_deref_803_addr_1_req_1,
          ackR => ptr_deref_803_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : ptr_deref_964_addr_0 
    SplitOperatorGroup86: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_964_root_address;
      ptr_deref_964_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_964_addr_0_req_0,
          ackL => ptr_deref_964_addr_0_ack_0,
          reqR => ptr_deref_964_addr_0_req_1,
          ackR => ptr_deref_964_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : ptr_deref_964_addr_1 
    SplitOperatorGroup87: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_964_root_address;
      ptr_deref_964_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_964_addr_1_req_0,
          ackL => ptr_deref_964_addr_1_ack_0,
          reqR => ptr_deref_964_addr_1_req_1,
          ackR => ptr_deref_964_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : ptr_deref_964_addr_2 
    SplitOperatorGroup88: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_964_root_address;
      ptr_deref_964_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_964_addr_2_req_0,
          ackL => ptr_deref_964_addr_2_ack_0,
          reqR => ptr_deref_964_addr_2_req_1,
          ackR => ptr_deref_964_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared split operator group (89) : ptr_deref_964_addr_3 
    SplitOperatorGroup89: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_964_root_address;
      ptr_deref_964_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_964_addr_3_req_0,
          ackL => ptr_deref_964_addr_3_ack_0,
          reqR => ptr_deref_964_addr_3_req_1,
          ackR => ptr_deref_964_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 89
    -- shared split operator group (90) : ptr_deref_985_addr_0 
    SplitOperatorGroup90: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_985_root_address;
      ptr_deref_985_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_985_addr_0_req_0,
          ackL => ptr_deref_985_addr_0_ack_0,
          reqR => ptr_deref_985_addr_0_req_1,
          ackR => ptr_deref_985_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 90
    -- shared split operator group (91) : ptr_deref_985_addr_1 
    SplitOperatorGroup91: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_985_root_address;
      ptr_deref_985_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_985_addr_1_req_0,
          ackL => ptr_deref_985_addr_1_ack_0,
          reqR => ptr_deref_985_addr_1_req_1,
          ackR => ptr_deref_985_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : ptr_deref_985_addr_2 
    SplitOperatorGroup92: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_985_root_address;
      ptr_deref_985_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_985_addr_2_req_0,
          ackL => ptr_deref_985_addr_2_ack_0,
          reqR => ptr_deref_985_addr_2_req_1,
          ackR => ptr_deref_985_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- shared split operator group (93) : ptr_deref_985_addr_3 
    SplitOperatorGroup93: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_985_root_address;
      ptr_deref_985_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_985_addr_3_req_0,
          ackL => ptr_deref_985_addr_3_ack_0,
          reqR => ptr_deref_985_addr_3_req_1,
          ackR => ptr_deref_985_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared load operator group (0) : ptr_deref_621_load_0 ptr_deref_621_load_3 ptr_deref_621_load_1 ptr_deref_553_load_0 ptr_deref_621_load_2 ptr_deref_569_load_0 ptr_deref_569_load_3 ptr_deref_553_load_3 ptr_deref_569_load_2 ptr_deref_553_load_2 ptr_deref_803_load_1 ptr_deref_803_load_0 ptr_deref_553_load_1 ptr_deref_882_load_0 ptr_deref_569_load_1 ptr_deref_1041_load_0 ptr_deref_1041_load_1 ptr_deref_1041_load_2 ptr_deref_1041_load_3 ptr_deref_1071_load_0 ptr_deref_1071_load_1 ptr_deref_1071_load_2 ptr_deref_1071_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(367 downto 0);
      signal data_out: std_logic_vector(183 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 22 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_621_load_0_req_0,
        ptr_deref_621_load_0_ack_0,
        ptr_deref_621_load_0_req_1,
        ptr_deref_621_load_0_ack_1,
        "ptr_deref_621_load_0",
        "memory_space_5" ,
        ptr_deref_621_data_0,
        ptr_deref_621_word_address_0,
        "ptr_deref_621_data_0",
        "ptr_deref_621_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_621_load_3_req_0,
        ptr_deref_621_load_3_ack_0,
        ptr_deref_621_load_3_req_1,
        ptr_deref_621_load_3_ack_1,
        "ptr_deref_621_load_3",
        "memory_space_5" ,
        ptr_deref_621_data_3,
        ptr_deref_621_word_address_3,
        "ptr_deref_621_data_3",
        "ptr_deref_621_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_621_load_1_req_0,
        ptr_deref_621_load_1_ack_0,
        ptr_deref_621_load_1_req_1,
        ptr_deref_621_load_1_ack_1,
        "ptr_deref_621_load_1",
        "memory_space_5" ,
        ptr_deref_621_data_1,
        ptr_deref_621_word_address_1,
        "ptr_deref_621_data_1",
        "ptr_deref_621_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_0_req_0,
        ptr_deref_553_load_0_ack_0,
        ptr_deref_553_load_0_req_1,
        ptr_deref_553_load_0_ack_1,
        "ptr_deref_553_load_0",
        "memory_space_5" ,
        ptr_deref_553_data_0,
        ptr_deref_553_word_address_0,
        "ptr_deref_553_data_0",
        "ptr_deref_553_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_621_load_2_req_0,
        ptr_deref_621_load_2_ack_0,
        ptr_deref_621_load_2_req_1,
        ptr_deref_621_load_2_ack_1,
        "ptr_deref_621_load_2",
        "memory_space_5" ,
        ptr_deref_621_data_2,
        ptr_deref_621_word_address_2,
        "ptr_deref_621_data_2",
        "ptr_deref_621_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_0_req_0,
        ptr_deref_569_load_0_ack_0,
        ptr_deref_569_load_0_req_1,
        ptr_deref_569_load_0_ack_1,
        "ptr_deref_569_load_0",
        "memory_space_5" ,
        ptr_deref_569_data_0,
        ptr_deref_569_word_address_0,
        "ptr_deref_569_data_0",
        "ptr_deref_569_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_3_req_0,
        ptr_deref_569_load_3_ack_0,
        ptr_deref_569_load_3_req_1,
        ptr_deref_569_load_3_ack_1,
        "ptr_deref_569_load_3",
        "memory_space_5" ,
        ptr_deref_569_data_3,
        ptr_deref_569_word_address_3,
        "ptr_deref_569_data_3",
        "ptr_deref_569_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_3_req_0,
        ptr_deref_553_load_3_ack_0,
        ptr_deref_553_load_3_req_1,
        ptr_deref_553_load_3_ack_1,
        "ptr_deref_553_load_3",
        "memory_space_5" ,
        ptr_deref_553_data_3,
        ptr_deref_553_word_address_3,
        "ptr_deref_553_data_3",
        "ptr_deref_553_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_2_req_0,
        ptr_deref_569_load_2_ack_0,
        ptr_deref_569_load_2_req_1,
        ptr_deref_569_load_2_ack_1,
        "ptr_deref_569_load_2",
        "memory_space_5" ,
        ptr_deref_569_data_2,
        ptr_deref_569_word_address_2,
        "ptr_deref_569_data_2",
        "ptr_deref_569_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_2_req_0,
        ptr_deref_553_load_2_ack_0,
        ptr_deref_553_load_2_req_1,
        ptr_deref_553_load_2_ack_1,
        "ptr_deref_553_load_2",
        "memory_space_5" ,
        ptr_deref_553_data_2,
        ptr_deref_553_word_address_2,
        "ptr_deref_553_data_2",
        "ptr_deref_553_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_803_load_1_req_0,
        ptr_deref_803_load_1_ack_0,
        ptr_deref_803_load_1_req_1,
        ptr_deref_803_load_1_ack_1,
        "ptr_deref_803_load_1",
        "memory_space_5" ,
        ptr_deref_803_data_1,
        ptr_deref_803_word_address_1,
        "ptr_deref_803_data_1",
        "ptr_deref_803_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_803_load_0_req_0,
        ptr_deref_803_load_0_ack_0,
        ptr_deref_803_load_0_req_1,
        ptr_deref_803_load_0_ack_1,
        "ptr_deref_803_load_0",
        "memory_space_5" ,
        ptr_deref_803_data_0,
        ptr_deref_803_word_address_0,
        "ptr_deref_803_data_0",
        "ptr_deref_803_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_553_load_1_req_0,
        ptr_deref_553_load_1_ack_0,
        ptr_deref_553_load_1_req_1,
        ptr_deref_553_load_1_ack_1,
        "ptr_deref_553_load_1",
        "memory_space_5" ,
        ptr_deref_553_data_1,
        ptr_deref_553_word_address_1,
        "ptr_deref_553_data_1",
        "ptr_deref_553_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_882_load_0_req_0,
        ptr_deref_882_load_0_ack_0,
        ptr_deref_882_load_0_req_1,
        ptr_deref_882_load_0_ack_1,
        "ptr_deref_882_load_0",
        "memory_space_5" ,
        ptr_deref_882_data_0,
        ptr_deref_882_word_address_0,
        "ptr_deref_882_data_0",
        "ptr_deref_882_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_569_load_1_req_0,
        ptr_deref_569_load_1_ack_0,
        ptr_deref_569_load_1_req_1,
        ptr_deref_569_load_1_ack_1,
        "ptr_deref_569_load_1",
        "memory_space_5" ,
        ptr_deref_569_data_1,
        ptr_deref_569_word_address_1,
        "ptr_deref_569_data_1",
        "ptr_deref_569_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1041_load_0_req_0,
        ptr_deref_1041_load_0_ack_0,
        ptr_deref_1041_load_0_req_1,
        ptr_deref_1041_load_0_ack_1,
        "ptr_deref_1041_load_0",
        "memory_space_5" ,
        ptr_deref_1041_data_0,
        ptr_deref_1041_word_address_0,
        "ptr_deref_1041_data_0",
        "ptr_deref_1041_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1041_load_1_req_0,
        ptr_deref_1041_load_1_ack_0,
        ptr_deref_1041_load_1_req_1,
        ptr_deref_1041_load_1_ack_1,
        "ptr_deref_1041_load_1",
        "memory_space_5" ,
        ptr_deref_1041_data_1,
        ptr_deref_1041_word_address_1,
        "ptr_deref_1041_data_1",
        "ptr_deref_1041_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1041_load_2_req_0,
        ptr_deref_1041_load_2_ack_0,
        ptr_deref_1041_load_2_req_1,
        ptr_deref_1041_load_2_ack_1,
        "ptr_deref_1041_load_2",
        "memory_space_5" ,
        ptr_deref_1041_data_2,
        ptr_deref_1041_word_address_2,
        "ptr_deref_1041_data_2",
        "ptr_deref_1041_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1041_load_3_req_0,
        ptr_deref_1041_load_3_ack_0,
        ptr_deref_1041_load_3_req_1,
        ptr_deref_1041_load_3_ack_1,
        "ptr_deref_1041_load_3",
        "memory_space_5" ,
        ptr_deref_1041_data_3,
        ptr_deref_1041_word_address_3,
        "ptr_deref_1041_data_3",
        "ptr_deref_1041_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1071_load_0_req_0,
        ptr_deref_1071_load_0_ack_0,
        ptr_deref_1071_load_0_req_1,
        ptr_deref_1071_load_0_ack_1,
        "ptr_deref_1071_load_0",
        "memory_space_5" ,
        ptr_deref_1071_data_0,
        ptr_deref_1071_word_address_0,
        "ptr_deref_1071_data_0",
        "ptr_deref_1071_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1071_load_1_req_0,
        ptr_deref_1071_load_1_ack_0,
        ptr_deref_1071_load_1_req_1,
        ptr_deref_1071_load_1_ack_1,
        "ptr_deref_1071_load_1",
        "memory_space_5" ,
        ptr_deref_1071_data_1,
        ptr_deref_1071_word_address_1,
        "ptr_deref_1071_data_1",
        "ptr_deref_1071_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1071_load_2_req_0,
        ptr_deref_1071_load_2_ack_0,
        ptr_deref_1071_load_2_req_1,
        ptr_deref_1071_load_2_ack_1,
        "ptr_deref_1071_load_2",
        "memory_space_5" ,
        ptr_deref_1071_data_2,
        ptr_deref_1071_word_address_2,
        "ptr_deref_1071_data_2",
        "ptr_deref_1071_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1071_load_3_req_0,
        ptr_deref_1071_load_3_ack_0,
        ptr_deref_1071_load_3_req_1,
        ptr_deref_1071_load_3_ack_1,
        "ptr_deref_1071_load_3",
        "memory_space_5" ,
        ptr_deref_1071_data_3,
        ptr_deref_1071_word_address_3,
        "ptr_deref_1071_data_3",
        "ptr_deref_1071_word_address_3" -- 
      );
      reqL(22) <= ptr_deref_621_load_0_req_0;
      reqL(21) <= ptr_deref_621_load_3_req_0;
      reqL(20) <= ptr_deref_621_load_1_req_0;
      reqL(19) <= ptr_deref_553_load_0_req_0;
      reqL(18) <= ptr_deref_621_load_2_req_0;
      reqL(17) <= ptr_deref_569_load_0_req_0;
      reqL(16) <= ptr_deref_569_load_3_req_0;
      reqL(15) <= ptr_deref_553_load_3_req_0;
      reqL(14) <= ptr_deref_569_load_2_req_0;
      reqL(13) <= ptr_deref_553_load_2_req_0;
      reqL(12) <= ptr_deref_803_load_1_req_0;
      reqL(11) <= ptr_deref_803_load_0_req_0;
      reqL(10) <= ptr_deref_553_load_1_req_0;
      reqL(9) <= ptr_deref_882_load_0_req_0;
      reqL(8) <= ptr_deref_569_load_1_req_0;
      reqL(7) <= ptr_deref_1041_load_0_req_0;
      reqL(6) <= ptr_deref_1041_load_1_req_0;
      reqL(5) <= ptr_deref_1041_load_2_req_0;
      reqL(4) <= ptr_deref_1041_load_3_req_0;
      reqL(3) <= ptr_deref_1071_load_0_req_0;
      reqL(2) <= ptr_deref_1071_load_1_req_0;
      reqL(1) <= ptr_deref_1071_load_2_req_0;
      reqL(0) <= ptr_deref_1071_load_3_req_0;
      ptr_deref_621_load_0_ack_0 <= ackL(22);
      ptr_deref_621_load_3_ack_0 <= ackL(21);
      ptr_deref_621_load_1_ack_0 <= ackL(20);
      ptr_deref_553_load_0_ack_0 <= ackL(19);
      ptr_deref_621_load_2_ack_0 <= ackL(18);
      ptr_deref_569_load_0_ack_0 <= ackL(17);
      ptr_deref_569_load_3_ack_0 <= ackL(16);
      ptr_deref_553_load_3_ack_0 <= ackL(15);
      ptr_deref_569_load_2_ack_0 <= ackL(14);
      ptr_deref_553_load_2_ack_0 <= ackL(13);
      ptr_deref_803_load_1_ack_0 <= ackL(12);
      ptr_deref_803_load_0_ack_0 <= ackL(11);
      ptr_deref_553_load_1_ack_0 <= ackL(10);
      ptr_deref_882_load_0_ack_0 <= ackL(9);
      ptr_deref_569_load_1_ack_0 <= ackL(8);
      ptr_deref_1041_load_0_ack_0 <= ackL(7);
      ptr_deref_1041_load_1_ack_0 <= ackL(6);
      ptr_deref_1041_load_2_ack_0 <= ackL(5);
      ptr_deref_1041_load_3_ack_0 <= ackL(4);
      ptr_deref_1071_load_0_ack_0 <= ackL(3);
      ptr_deref_1071_load_1_ack_0 <= ackL(2);
      ptr_deref_1071_load_2_ack_0 <= ackL(1);
      ptr_deref_1071_load_3_ack_0 <= ackL(0);
      reqR(22) <= ptr_deref_621_load_0_req_1;
      reqR(21) <= ptr_deref_621_load_3_req_1;
      reqR(20) <= ptr_deref_621_load_1_req_1;
      reqR(19) <= ptr_deref_553_load_0_req_1;
      reqR(18) <= ptr_deref_621_load_2_req_1;
      reqR(17) <= ptr_deref_569_load_0_req_1;
      reqR(16) <= ptr_deref_569_load_3_req_1;
      reqR(15) <= ptr_deref_553_load_3_req_1;
      reqR(14) <= ptr_deref_569_load_2_req_1;
      reqR(13) <= ptr_deref_553_load_2_req_1;
      reqR(12) <= ptr_deref_803_load_1_req_1;
      reqR(11) <= ptr_deref_803_load_0_req_1;
      reqR(10) <= ptr_deref_553_load_1_req_1;
      reqR(9) <= ptr_deref_882_load_0_req_1;
      reqR(8) <= ptr_deref_569_load_1_req_1;
      reqR(7) <= ptr_deref_1041_load_0_req_1;
      reqR(6) <= ptr_deref_1041_load_1_req_1;
      reqR(5) <= ptr_deref_1041_load_2_req_1;
      reqR(4) <= ptr_deref_1041_load_3_req_1;
      reqR(3) <= ptr_deref_1071_load_0_req_1;
      reqR(2) <= ptr_deref_1071_load_1_req_1;
      reqR(1) <= ptr_deref_1071_load_2_req_1;
      reqR(0) <= ptr_deref_1071_load_3_req_1;
      ptr_deref_621_load_0_ack_1 <= ackR(22);
      ptr_deref_621_load_3_ack_1 <= ackR(21);
      ptr_deref_621_load_1_ack_1 <= ackR(20);
      ptr_deref_553_load_0_ack_1 <= ackR(19);
      ptr_deref_621_load_2_ack_1 <= ackR(18);
      ptr_deref_569_load_0_ack_1 <= ackR(17);
      ptr_deref_569_load_3_ack_1 <= ackR(16);
      ptr_deref_553_load_3_ack_1 <= ackR(15);
      ptr_deref_569_load_2_ack_1 <= ackR(14);
      ptr_deref_553_load_2_ack_1 <= ackR(13);
      ptr_deref_803_load_1_ack_1 <= ackR(12);
      ptr_deref_803_load_0_ack_1 <= ackR(11);
      ptr_deref_553_load_1_ack_1 <= ackR(10);
      ptr_deref_882_load_0_ack_1 <= ackR(9);
      ptr_deref_569_load_1_ack_1 <= ackR(8);
      ptr_deref_1041_load_0_ack_1 <= ackR(7);
      ptr_deref_1041_load_1_ack_1 <= ackR(6);
      ptr_deref_1041_load_2_ack_1 <= ackR(5);
      ptr_deref_1041_load_3_ack_1 <= ackR(4);
      ptr_deref_1071_load_0_ack_1 <= ackR(3);
      ptr_deref_1071_load_1_ack_1 <= ackR(2);
      ptr_deref_1071_load_2_ack_1 <= ackR(1);
      ptr_deref_1071_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_621_word_address_0 & ptr_deref_621_word_address_3 & ptr_deref_621_word_address_1 & ptr_deref_553_word_address_0 & ptr_deref_621_word_address_2 & ptr_deref_569_word_address_0 & ptr_deref_569_word_address_3 & ptr_deref_553_word_address_3 & ptr_deref_569_word_address_2 & ptr_deref_553_word_address_2 & ptr_deref_803_word_address_1 & ptr_deref_803_word_address_0 & ptr_deref_553_word_address_1 & ptr_deref_882_word_address_0 & ptr_deref_569_word_address_1 & ptr_deref_1041_word_address_0 & ptr_deref_1041_word_address_1 & ptr_deref_1041_word_address_2 & ptr_deref_1041_word_address_3 & ptr_deref_1071_word_address_0 & ptr_deref_1071_word_address_1 & ptr_deref_1071_word_address_2 & ptr_deref_1071_word_address_3;
      ptr_deref_621_data_0 <= data_out(183 downto 176);
      ptr_deref_621_data_3 <= data_out(175 downto 168);
      ptr_deref_621_data_1 <= data_out(167 downto 160);
      ptr_deref_553_data_0 <= data_out(159 downto 152);
      ptr_deref_621_data_2 <= data_out(151 downto 144);
      ptr_deref_569_data_0 <= data_out(143 downto 136);
      ptr_deref_569_data_3 <= data_out(135 downto 128);
      ptr_deref_553_data_3 <= data_out(127 downto 120);
      ptr_deref_569_data_2 <= data_out(119 downto 112);
      ptr_deref_553_data_2 <= data_out(111 downto 104);
      ptr_deref_803_data_1 <= data_out(103 downto 96);
      ptr_deref_803_data_0 <= data_out(95 downto 88);
      ptr_deref_553_data_1 <= data_out(87 downto 80);
      ptr_deref_882_data_0 <= data_out(79 downto 72);
      ptr_deref_569_data_1 <= data_out(71 downto 64);
      ptr_deref_1041_data_0 <= data_out(63 downto 56);
      ptr_deref_1041_data_1 <= data_out(55 downto 48);
      ptr_deref_1041_data_2 <= data_out(47 downto 40);
      ptr_deref_1041_data_3 <= data_out(39 downto 32);
      ptr_deref_1071_data_0 <= data_out(31 downto 24);
      ptr_deref_1071_data_1 <= data_out(23 downto 16);
      ptr_deref_1071_data_2 <= data_out(15 downto 8);
      ptr_deref_1071_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 23,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 23,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_964_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_964_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_964_word_address_0) &  " data ptr_deref_964_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_964_data_0) severity note; --
        end if;
        if ptr_deref_964_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_964_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_964_word_address_3) &  " data ptr_deref_964_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_964_data_3) severity note; --
        end if;
        if ptr_deref_964_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_964_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_964_word_address_1) &  " data ptr_deref_964_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_964_data_1) severity note; --
        end if;
        if ptr_deref_964_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_964_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_964_word_address_2) &  " data ptr_deref_964_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_964_data_2) severity note; --
        end if;
        if ptr_deref_985_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_985_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_985_word_address_0) &  " data ptr_deref_985_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_985_data_0) severity note; --
        end if;
        if ptr_deref_985_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_985_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_985_word_address_1) &  " data ptr_deref_985_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_985_data_1) severity note; --
        end if;
        if ptr_deref_985_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_985_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_985_word_address_2) &  " data ptr_deref_985_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_985_data_2) severity note; --
        end if;
        if ptr_deref_985_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_985_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_985_word_address_3) &  " data ptr_deref_985_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_985_data_3) severity note; --
        end if;
        if ptr_deref_1027_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1027_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1027_word_address_0) &  " data ptr_deref_1027_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1027_data_0) severity note; --
        end if;
        if ptr_deref_1027_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1027_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1027_word_address_1) &  " data ptr_deref_1027_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1027_data_1) severity note; --
        end if;
        if ptr_deref_1027_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1027_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1027_word_address_2) &  " data ptr_deref_1027_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1027_data_2) severity note; --
        end if;
        if ptr_deref_1027_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1027_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1027_word_address_3) &  " data ptr_deref_1027_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1027_data_3) severity note; --
        end if;
        if ptr_deref_1055_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1055_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1055_word_address_0) &  " data ptr_deref_1055_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1055_data_0) severity note; --
        end if;
        if ptr_deref_1055_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1055_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1055_word_address_1) &  " data ptr_deref_1055_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1055_data_1) severity note; --
        end if;
        if ptr_deref_1055_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1055_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1055_word_address_2) &  " data ptr_deref_1055_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1055_data_2) severity note; --
        end if;
        if ptr_deref_1055_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1055_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1055_word_address_3) &  " data ptr_deref_1055_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1055_data_3) severity note; --
        end if;
        if ptr_deref_1085_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1085_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1085_word_address_0) &  " data ptr_deref_1085_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1085_data_0) severity note; --
        end if;
        if ptr_deref_1085_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1085_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1085_word_address_1) &  " data ptr_deref_1085_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1085_data_1) severity note; --
        end if;
        if ptr_deref_1085_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1085_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1085_word_address_2) &  " data ptr_deref_1085_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1085_data_2) severity note; --
        end if;
        if ptr_deref_1085_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1085_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1085_word_address_3) &  " data ptr_deref_1085_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1085_data_3) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_964_store_0 ptr_deref_964_store_3 ptr_deref_964_store_1 ptr_deref_964_store_2 ptr_deref_985_store_0 ptr_deref_985_store_1 ptr_deref_985_store_2 ptr_deref_985_store_3 ptr_deref_1027_store_0 ptr_deref_1027_store_1 ptr_deref_1027_store_2 ptr_deref_1027_store_3 ptr_deref_1055_store_0 ptr_deref_1055_store_1 ptr_deref_1055_store_2 ptr_deref_1055_store_3 ptr_deref_1085_store_0 ptr_deref_1085_store_1 ptr_deref_1085_store_2 ptr_deref_1085_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(319 downto 0);
      signal data_in: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 19 downto 0);
      -- 
    begin -- 
      reqL(19) <= ptr_deref_964_store_0_req_0;
      reqL(18) <= ptr_deref_964_store_3_req_0;
      reqL(17) <= ptr_deref_964_store_1_req_0;
      reqL(16) <= ptr_deref_964_store_2_req_0;
      reqL(15) <= ptr_deref_985_store_0_req_0;
      reqL(14) <= ptr_deref_985_store_1_req_0;
      reqL(13) <= ptr_deref_985_store_2_req_0;
      reqL(12) <= ptr_deref_985_store_3_req_0;
      reqL(11) <= ptr_deref_1027_store_0_req_0;
      reqL(10) <= ptr_deref_1027_store_1_req_0;
      reqL(9) <= ptr_deref_1027_store_2_req_0;
      reqL(8) <= ptr_deref_1027_store_3_req_0;
      reqL(7) <= ptr_deref_1055_store_0_req_0;
      reqL(6) <= ptr_deref_1055_store_1_req_0;
      reqL(5) <= ptr_deref_1055_store_2_req_0;
      reqL(4) <= ptr_deref_1055_store_3_req_0;
      reqL(3) <= ptr_deref_1085_store_0_req_0;
      reqL(2) <= ptr_deref_1085_store_1_req_0;
      reqL(1) <= ptr_deref_1085_store_2_req_0;
      reqL(0) <= ptr_deref_1085_store_3_req_0;
      ptr_deref_964_store_0_ack_0 <= ackL(19);
      ptr_deref_964_store_3_ack_0 <= ackL(18);
      ptr_deref_964_store_1_ack_0 <= ackL(17);
      ptr_deref_964_store_2_ack_0 <= ackL(16);
      ptr_deref_985_store_0_ack_0 <= ackL(15);
      ptr_deref_985_store_1_ack_0 <= ackL(14);
      ptr_deref_985_store_2_ack_0 <= ackL(13);
      ptr_deref_985_store_3_ack_0 <= ackL(12);
      ptr_deref_1027_store_0_ack_0 <= ackL(11);
      ptr_deref_1027_store_1_ack_0 <= ackL(10);
      ptr_deref_1027_store_2_ack_0 <= ackL(9);
      ptr_deref_1027_store_3_ack_0 <= ackL(8);
      ptr_deref_1055_store_0_ack_0 <= ackL(7);
      ptr_deref_1055_store_1_ack_0 <= ackL(6);
      ptr_deref_1055_store_2_ack_0 <= ackL(5);
      ptr_deref_1055_store_3_ack_0 <= ackL(4);
      ptr_deref_1085_store_0_ack_0 <= ackL(3);
      ptr_deref_1085_store_1_ack_0 <= ackL(2);
      ptr_deref_1085_store_2_ack_0 <= ackL(1);
      ptr_deref_1085_store_3_ack_0 <= ackL(0);
      reqR(19) <= ptr_deref_964_store_0_req_1;
      reqR(18) <= ptr_deref_964_store_3_req_1;
      reqR(17) <= ptr_deref_964_store_1_req_1;
      reqR(16) <= ptr_deref_964_store_2_req_1;
      reqR(15) <= ptr_deref_985_store_0_req_1;
      reqR(14) <= ptr_deref_985_store_1_req_1;
      reqR(13) <= ptr_deref_985_store_2_req_1;
      reqR(12) <= ptr_deref_985_store_3_req_1;
      reqR(11) <= ptr_deref_1027_store_0_req_1;
      reqR(10) <= ptr_deref_1027_store_1_req_1;
      reqR(9) <= ptr_deref_1027_store_2_req_1;
      reqR(8) <= ptr_deref_1027_store_3_req_1;
      reqR(7) <= ptr_deref_1055_store_0_req_1;
      reqR(6) <= ptr_deref_1055_store_1_req_1;
      reqR(5) <= ptr_deref_1055_store_2_req_1;
      reqR(4) <= ptr_deref_1055_store_3_req_1;
      reqR(3) <= ptr_deref_1085_store_0_req_1;
      reqR(2) <= ptr_deref_1085_store_1_req_1;
      reqR(1) <= ptr_deref_1085_store_2_req_1;
      reqR(0) <= ptr_deref_1085_store_3_req_1;
      ptr_deref_964_store_0_ack_1 <= ackR(19);
      ptr_deref_964_store_3_ack_1 <= ackR(18);
      ptr_deref_964_store_1_ack_1 <= ackR(17);
      ptr_deref_964_store_2_ack_1 <= ackR(16);
      ptr_deref_985_store_0_ack_1 <= ackR(15);
      ptr_deref_985_store_1_ack_1 <= ackR(14);
      ptr_deref_985_store_2_ack_1 <= ackR(13);
      ptr_deref_985_store_3_ack_1 <= ackR(12);
      ptr_deref_1027_store_0_ack_1 <= ackR(11);
      ptr_deref_1027_store_1_ack_1 <= ackR(10);
      ptr_deref_1027_store_2_ack_1 <= ackR(9);
      ptr_deref_1027_store_3_ack_1 <= ackR(8);
      ptr_deref_1055_store_0_ack_1 <= ackR(7);
      ptr_deref_1055_store_1_ack_1 <= ackR(6);
      ptr_deref_1055_store_2_ack_1 <= ackR(5);
      ptr_deref_1055_store_3_ack_1 <= ackR(4);
      ptr_deref_1085_store_0_ack_1 <= ackR(3);
      ptr_deref_1085_store_1_ack_1 <= ackR(2);
      ptr_deref_1085_store_2_ack_1 <= ackR(1);
      ptr_deref_1085_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_964_word_address_0 & ptr_deref_964_word_address_3 & ptr_deref_964_word_address_1 & ptr_deref_964_word_address_2 & ptr_deref_985_word_address_0 & ptr_deref_985_word_address_1 & ptr_deref_985_word_address_2 & ptr_deref_985_word_address_3 & ptr_deref_1027_word_address_0 & ptr_deref_1027_word_address_1 & ptr_deref_1027_word_address_2 & ptr_deref_1027_word_address_3 & ptr_deref_1055_word_address_0 & ptr_deref_1055_word_address_1 & ptr_deref_1055_word_address_2 & ptr_deref_1055_word_address_3 & ptr_deref_1085_word_address_0 & ptr_deref_1085_word_address_1 & ptr_deref_1085_word_address_2 & ptr_deref_1085_word_address_3;
      data_in <= ptr_deref_964_data_0 & ptr_deref_964_data_3 & ptr_deref_964_data_1 & ptr_deref_964_data_2 & ptr_deref_985_data_0 & ptr_deref_985_data_1 & ptr_deref_985_data_2 & ptr_deref_985_data_3 & ptr_deref_1027_data_0 & ptr_deref_1027_data_1 & ptr_deref_1027_data_2 & ptr_deref_1027_data_3 & ptr_deref_1055_data_0 & ptr_deref_1055_data_1 & ptr_deref_1055_data_2 & ptr_deref_1055_data_3 & ptr_deref_1085_data_0 & ptr_deref_1085_data_1 & ptr_deref_1085_data_2 & ptr_deref_1085_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 20,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 20,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_537_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_537_inst_ack_0 then -- 
            assert false report " ReadPipe chk_in0 to wire simple_obj_ref_537_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_537_inst_req_0;
      simple_obj_ref_537_inst_ack_0 <= ack(0);
      simple_obj_ref_537_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => chk_in0_pipe_read_req(0),
          oack => chk_in0_pipe_read_ack(0),
          odata => chk_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1105_inst_ack_0 then -- 
          assert false report " WritePipe rtt_in0 from wire type_cast_1107_wire value="  &  convert_slv_to_hex_string(type_cast_1107_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1105_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1105_inst_req_0;
      simple_obj_ref_1105_inst_ack_0 <= ack(0);
      data_in <= type_cast_1107_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => rtt_in0_pipe_write_req(0),
          oack => rtt_in0_pipe_write_ack(0),
          odata => rtt_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_687_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_690_wire value="  &  convert_slv_to_hex_string(binary_690_wire) severity note; --
        end if;
        if simple_obj_ref_653_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_656_wire value="  &  convert_slv_to_hex_string(binary_656_wire) severity note; --
        end if;
        if simple_obj_ref_725_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_728_wire value="  &  convert_slv_to_hex_string(binary_728_wire) severity note; --
        end if;
        if simple_obj_ref_948_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_951_wire value="  &  convert_slv_to_hex_string(binary_951_wire) severity note; --
        end if;
        if simple_obj_ref_607_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_610_wire value="  &  convert_slv_to_hex_string(binary_610_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_687_inst simple_obj_ref_653_inst simple_obj_ref_725_inst simple_obj_ref_948_inst simple_obj_ref_607_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal req, ack : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      req(4) <= simple_obj_ref_687_inst_req_0;
      req(3) <= simple_obj_ref_653_inst_req_0;
      req(2) <= simple_obj_ref_725_inst_req_0;
      req(1) <= simple_obj_ref_948_inst_req_0;
      req(0) <= simple_obj_ref_607_inst_req_0;
      simple_obj_ref_687_inst_ack_0 <= ack(4);
      simple_obj_ref_653_inst_ack_0 <= ack(3);
      simple_obj_ref_725_inst_ack_0 <= ack(2);
      simple_obj_ref_948_inst_ack_0 <= ack(1);
      simple_obj_ref_607_inst_ack_0 <= ack(0);
      data_in <= binary_690_wire & binary_656_wire & binary_728_wire & binary_951_wire & binary_610_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 5,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_697_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_697_call_req_0;
      call_stmt_697_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_697_call_req_1;
      call_stmt_697_call_ack_1 <= ackR(0);
      data_in <= tmp35x_xi_644;
      tmp32_697 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 16,
        owidth => 16,
        twidth => 2,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 16, twidth => 2, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_chk_1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_chk_1;
architecture Default of ahir_glue_chk_1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_chk_1_CP_4158_start: Boolean;
  -- links between control-path and data-path
  signal binary_1285_inst_ack_0 : boolean;
  signal type_cast_1173_inst_ack_0 : boolean;
  signal binary_1190_inst_ack_0 : boolean;
  signal ptr_deref_1201_load_2_req_0 : boolean;
  signal ptr_deref_1201_addr_0_ack_1 : boolean;
  signal binary_1163_inst_req_0 : boolean;
  signal ptr_deref_1201_addr_0_ack_0 : boolean;
  signal ptr_deref_1150_load_0_req_1 : boolean;
  signal ptr_deref_1201_addr_2_req_1 : boolean;
  signal binary_1213_inst_req_1 : boolean;
  signal ptr_deref_1201_addr_3_ack_1 : boolean;
  signal type_cast_1280_inst_req_0 : boolean;
  signal if_stmt_1179_branch_req_0 : boolean;
  signal binary_1295_inst_ack_0 : boolean;
  signal ptr_deref_1150_gather_scatter_ack_0 : boolean;
  signal binary_1285_inst_ack_1 : boolean;
  signal ptr_deref_1201_addr_3_req_0 : boolean;
  signal ptr_deref_1201_addr_1_ack_0 : boolean;
  signal binary_1207_inst_req_1 : boolean;
  signal ptr_deref_1150_load_2_ack_1 : boolean;
  signal ptr_deref_1201_addr_3_req_1 : boolean;
  signal ptr_deref_1201_addr_3_ack_0 : boolean;
  signal binary_1270_inst_req_1 : boolean;
  signal ptr_deref_1201_load_1_ack_0 : boolean;
  signal ptr_deref_1201_load_1_req_0 : boolean;
  signal binary_1290_inst_req_0 : boolean;
  signal phi_stmt_1334_req_1 : boolean;
  signal ptr_deref_1201_load_0_ack_0 : boolean;
  signal ptr_deref_1150_load_3_ack_1 : boolean;
  signal ptr_deref_1150_load_2_req_1 : boolean;
  signal binary_1257_inst_ack_1 : boolean;
  signal binary_1257_inst_req_1 : boolean;
  signal ptr_deref_1201_load_0_req_0 : boolean;
  signal binary_1257_inst_ack_0 : boolean;
  signal ptr_deref_1150_load_0_ack_1 : boolean;
  signal binary_1671_inst_ack_1 : boolean;
  signal binary_1257_inst_req_0 : boolean;
  signal type_cast_1158_inst_ack_0 : boolean;
  signal ptr_deref_1150_gather_scatter_req_0 : boolean;
  signal ptr_deref_1201_addr_2_ack_1 : boolean;
  signal binary_1207_inst_ack_1 : boolean;
  signal type_cast_1158_inst_req_0 : boolean;
  signal binary_1213_inst_ack_1 : boolean;
  signal if_stmt_1259_branch_ack_0 : boolean;
  signal ptr_deref_1201_addr_0_req_0 : boolean;
  signal ptr_deref_1150_load_3_req_1 : boolean;
  signal ptr_deref_1564_base_resize_ack_0 : boolean;
  signal if_stmt_1297_branch_ack_1 : boolean;
  signal if_stmt_1259_branch_req_0 : boolean;
  signal ptr_deref_1201_addr_0_req_1 : boolean;
  signal binary_1245_inst_ack_1 : boolean;
  signal binary_1207_inst_req_0 : boolean;
  signal ptr_deref_1201_root_address_inst_ack_0 : boolean;
  signal binary_1270_inst_req_0 : boolean;
  signal if_stmt_1179_branch_ack_1 : boolean;
  signal binary_1177_inst_req_0 : boolean;
  signal ptr_deref_1201_addr_1_req_1 : boolean;
  signal binary_1177_inst_ack_0 : boolean;
  signal binary_1213_inst_ack_0 : boolean;
  signal binary_1285_inst_req_0 : boolean;
  signal if_stmt_1179_branch_ack_0 : boolean;
  signal binary_1251_inst_req_0 : boolean;
  signal binary_1163_inst_ack_0 : boolean;
  signal ptr_deref_1201_addr_1_req_0 : boolean;
  signal ptr_deref_1201_load_2_ack_0 : boolean;
  signal binary_1169_inst_ack_1 : boolean;
  signal call_stmt_1277_call_req_1 : boolean;
  signal ptr_deref_1150_load_1_req_1 : boolean;
  signal binary_1295_inst_ack_1 : boolean;
  signal binary_1163_inst_req_1 : boolean;
  signal binary_1163_inst_ack_1 : boolean;
  signal binary_1251_inst_ack_0 : boolean;
  signal ptr_deref_1201_addr_1_ack_1 : boolean;
  signal ptr_deref_1201_load_3_ack_0 : boolean;
  signal binary_1270_inst_ack_0 : boolean;
  signal ptr_deref_1150_load_1_ack_1 : boolean;
  signal binary_1295_inst_req_1 : boolean;
  signal binary_1251_inst_req_1 : boolean;
  signal binary_1251_inst_ack_1 : boolean;
  signal binary_1207_inst_ack_0 : boolean;
  signal ptr_deref_1150_load_2_ack_0 : boolean;
  signal binary_1177_inst_req_1 : boolean;
  signal ptr_deref_1150_load_3_req_0 : boolean;
  signal ptr_deref_1150_load_3_ack_0 : boolean;
  signal call_stmt_1277_call_ack_1 : boolean;
  signal binary_1245_inst_req_0 : boolean;
  signal type_cast_1173_inst_req_0 : boolean;
  signal binary_1245_inst_ack_0 : boolean;
  signal ptr_deref_1201_base_resize_req_0 : boolean;
  signal binary_1177_inst_ack_1 : boolean;
  signal ptr_deref_1201_base_resize_ack_0 : boolean;
  signal binary_1245_inst_req_1 : boolean;
  signal ptr_deref_1201_root_address_inst_req_0 : boolean;
  signal ptr_deref_1564_root_address_inst_req_0 : boolean;
  signal ptr_deref_1201_addr_2_req_0 : boolean;
  signal binary_1190_inst_req_0 : boolean;
  signal ptr_deref_1201_addr_2_ack_0 : boolean;
  signal binary_1213_inst_req_0 : boolean;
  signal binary_1190_inst_req_1 : boolean;
  signal simple_obj_ref_1305_inst_ack_0 : boolean;
  signal if_stmt_1259_branch_ack_1 : boolean;
  signal ptr_deref_1150_load_2_req_0 : boolean;
  signal binary_1169_inst_req_1 : boolean;
  signal binary_1308_inst_ack_0 : boolean;
  signal type_cast_1436_inst_req_0 : boolean;
  signal type_cast_1340_inst_ack_0 : boolean;
  signal type_cast_1280_inst_ack_0 : boolean;
  signal simple_obj_ref_1233_inst_ack_0 : boolean;
  signal type_cast_1347_inst_req_0 : boolean;
  signal simple_obj_ref_1233_inst_req_0 : boolean;
  signal binary_1671_inst_ack_0 : boolean;
  signal ptr_deref_1201_load_3_req_0 : boolean;
  signal type_cast_1197_inst_ack_0 : boolean;
  signal type_cast_1197_inst_req_0 : boolean;
  signal call_stmt_1277_call_ack_0 : boolean;
  signal binary_1295_inst_req_0 : boolean;
  signal binary_1671_inst_req_0 : boolean;
  signal type_cast_1436_inst_ack_0 : boolean;
  signal ptr_deref_1150_load_1_ack_0 : boolean;
  signal ptr_deref_1150_load_1_req_0 : boolean;
  signal type_cast_1119_inst_req_0 : boolean;
  signal type_cast_1119_inst_ack_0 : boolean;
  signal ptr_deref_1201_load_0_ack_1 : boolean;
  signal array_obj_ref_1130_root_address_inst_req_0 : boolean;
  signal type_cast_1123_inst_req_0 : boolean;
  signal type_cast_1123_inst_ack_0 : boolean;
  signal array_obj_ref_1130_base_resize_req_0 : boolean;
  signal array_obj_ref_1130_base_resize_ack_0 : boolean;
  signal binary_1219_inst_ack_1 : boolean;
  signal ptr_deref_1201_gather_scatter_req_0 : boolean;
  signal ptr_deref_1134_root_address_inst_req_0 : boolean;
  signal ptr_deref_1201_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1130_root_address_inst_ack_0 : boolean;
  signal binary_1671_inst_req_1 : boolean;
  signal ptr_deref_1134_base_resize_ack_0 : boolean;
  signal if_stmt_1297_branch_ack_0 : boolean;
  signal binary_1236_inst_req_1 : boolean;
  signal binary_1236_inst_ack_0 : boolean;
  signal binary_1236_inst_req_0 : boolean;
  signal ptr_deref_1134_addr_0_req_0 : boolean;
  signal ptr_deref_1201_load_3_ack_1 : boolean;
  signal ptr_deref_1134_addr_0_ack_0 : boolean;
  signal array_obj_ref_1130_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1150_load_0_req_0 : boolean;
  signal simple_obj_ref_1118_inst_req_0 : boolean;
  signal simple_obj_ref_1118_inst_ack_0 : boolean;
  signal array_obj_ref_1130_final_reg_req_0 : boolean;
  signal binary_1169_inst_ack_0 : boolean;
  signal array_obj_ref_1130_final_reg_ack_0 : boolean;
  signal ptr_deref_1134_base_resize_req_0 : boolean;
  signal type_cast_1340_inst_req_0 : boolean;
  signal binary_1169_inst_req_0 : boolean;
  signal binary_1236_inst_ack_1 : boolean;
  signal ptr_deref_1134_root_address_inst_ack_0 : boolean;
  signal binary_1353_inst_req_0 : boolean;
  signal binary_1353_inst_ack_0 : boolean;
  signal phi_stmt_1334_req_0 : boolean;
  signal binary_1353_inst_req_1 : boolean;
  signal binary_1353_inst_ack_1 : boolean;
  signal if_stmt_1673_branch_ack_0 : boolean;
  signal binary_1317_inst_ack_0 : boolean;
  signal if_stmt_1673_branch_req_0 : boolean;
  signal simple_obj_ref_1305_inst_req_0 : boolean;
  signal if_stmt_1319_branch_ack_0 : boolean;
  signal binary_1219_inst_req_0 : boolean;
  signal binary_1317_inst_req_0 : boolean;
  signal binary_1290_inst_ack_0 : boolean;
  signal binary_1219_inst_ack_0 : boolean;
  signal binary_1270_inst_ack_1 : boolean;
  signal binary_1308_inst_ack_1 : boolean;
  signal if_stmt_1319_branch_ack_1 : boolean;
  signal binary_1330_inst_ack_1 : boolean;
  signal if_stmt_1297_branch_req_0 : boolean;
  signal binary_1308_inst_req_0 : boolean;
  signal binary_1285_inst_req_1 : boolean;
  signal binary_1308_inst_req_1 : boolean;
  signal binary_1317_inst_req_1 : boolean;
  signal binary_1317_inst_ack_1 : boolean;
  signal ptr_deref_1201_load_0_req_1 : boolean;
  signal phi_stmt_1341_req_0 : boolean;
  signal type_cast_1154_inst_req_0 : boolean;
  signal binary_1219_inst_req_1 : boolean;
  signal binary_1330_inst_req_0 : boolean;
  signal binary_1330_inst_ack_0 : boolean;
  signal binary_1330_inst_req_1 : boolean;
  signal if_stmt_1319_branch_req_0 : boolean;
  signal type_cast_1154_inst_ack_0 : boolean;
  signal array_obj_ref_1130_root_address_inst_req_1 : boolean;
  signal ptr_deref_1150_load_0_ack_0 : boolean;
  signal ptr_deref_1134_addr_0_req_1 : boolean;
  signal ptr_deref_1134_addr_0_ack_1 : boolean;
  signal ptr_deref_1134_addr_1_req_0 : boolean;
  signal ptr_deref_1201_load_3_req_1 : boolean;
  signal ptr_deref_1134_addr_1_ack_0 : boolean;
  signal simple_obj_ref_1187_inst_ack_0 : boolean;
  signal ptr_deref_1134_addr_1_req_1 : boolean;
  signal ptr_deref_1134_addr_1_ack_1 : boolean;
  signal ptr_deref_1564_addr_2_ack_1 : boolean;
  signal ptr_deref_1134_addr_2_req_0 : boolean;
  signal ptr_deref_1134_addr_2_ack_0 : boolean;
  signal simple_obj_ref_1187_inst_req_0 : boolean;
  signal ptr_deref_1134_addr_2_req_1 : boolean;
  signal ptr_deref_1134_addr_2_ack_1 : boolean;
  signal ptr_deref_1134_addr_3_req_0 : boolean;
  signal ptr_deref_1134_addr_3_ack_0 : boolean;
  signal if_stmt_1225_branch_ack_0 : boolean;
  signal ptr_deref_1134_addr_3_req_1 : boolean;
  signal ptr_deref_1134_addr_3_ack_1 : boolean;
  signal if_stmt_1673_branch_ack_1 : boolean;
  signal ptr_deref_1134_load_0_req_0 : boolean;
  signal ptr_deref_1134_load_0_ack_0 : boolean;
  signal if_stmt_1225_branch_ack_1 : boolean;
  signal ptr_deref_1134_load_1_req_0 : boolean;
  signal ptr_deref_1201_load_2_ack_1 : boolean;
  signal ptr_deref_1134_load_1_ack_0 : boolean;
  signal ptr_deref_1134_load_2_req_0 : boolean;
  signal ptr_deref_1201_load_2_req_1 : boolean;
  signal ptr_deref_1134_load_2_ack_0 : boolean;
  signal call_stmt_1277_call_req_0 : boolean;
  signal if_stmt_1225_branch_req_0 : boolean;
  signal ptr_deref_1134_load_3_req_0 : boolean;
  signal ptr_deref_1134_load_3_ack_0 : boolean;
  signal binary_1290_inst_ack_1 : boolean;
  signal ptr_deref_1134_load_0_req_1 : boolean;
  signal ptr_deref_1134_load_0_ack_1 : boolean;
  signal binary_1290_inst_req_1 : boolean;
  signal ptr_deref_1134_load_1_req_1 : boolean;
  signal ptr_deref_1134_load_1_ack_1 : boolean;
  signal ptr_deref_1134_load_2_req_1 : boolean;
  signal ptr_deref_1201_load_1_ack_1 : boolean;
  signal ptr_deref_1134_load_2_ack_1 : boolean;
  signal type_cast_1223_inst_ack_0 : boolean;
  signal ptr_deref_1134_load_3_req_1 : boolean;
  signal ptr_deref_1201_load_1_req_1 : boolean;
  signal type_cast_1223_inst_req_0 : boolean;
  signal ptr_deref_1134_load_3_ack_1 : boolean;
  signal ptr_deref_1134_gather_scatter_req_0 : boolean;
  signal ptr_deref_1134_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1267_inst_ack_0 : boolean;
  signal binary_1190_inst_ack_1 : boolean;
  signal ptr_deref_1564_addr_0_ack_1 : boolean;
  signal array_obj_ref_1139_base_resize_req_0 : boolean;
  signal array_obj_ref_1139_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1267_inst_req_0 : boolean;
  signal ptr_deref_1564_addr_0_req_1 : boolean;
  signal array_obj_ref_1139_root_address_inst_req_0 : boolean;
  signal ptr_deref_1564_addr_1_req_0 : boolean;
  signal ptr_deref_1564_addr_1_ack_0 : boolean;
  signal array_obj_ref_1139_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1139_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1139_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1564_addr_1_req_1 : boolean;
  signal ptr_deref_1564_store_1_ack_0 : boolean;
  signal ptr_deref_1564_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1564_addr_1_ack_1 : boolean;
  signal array_obj_ref_1139_final_reg_req_0 : boolean;
  signal ptr_deref_1564_addr_3_req_0 : boolean;
  signal array_obj_ref_1139_final_reg_ack_0 : boolean;
  signal ptr_deref_1564_gather_scatter_req_0 : boolean;
  signal ptr_deref_1564_addr_3_ack_0 : boolean;
  signal ptr_deref_1564_addr_3_req_1 : boolean;
  signal ptr_deref_1564_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1564_addr_3_ack_1 : boolean;
  signal ptr_deref_1564_addr_2_req_0 : boolean;
  signal ptr_deref_1564_store_1_req_0 : boolean;
  signal array_obj_ref_1146_base_resize_req_0 : boolean;
  signal ptr_deref_1564_addr_2_ack_0 : boolean;
  signal array_obj_ref_1146_base_resize_ack_0 : boolean;
  signal ptr_deref_1564_store_2_req_0 : boolean;
  signal ptr_deref_1564_store_2_ack_0 : boolean;
  signal ptr_deref_1564_store_3_ack_0 : boolean;
  signal array_obj_ref_1146_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1146_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1146_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1146_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1564_store_3_req_0 : boolean;
  signal ptr_deref_1564_addr_0_req_0 : boolean;
  signal array_obj_ref_1146_final_reg_req_0 : boolean;
  signal array_obj_ref_1146_final_reg_ack_0 : boolean;
  signal ptr_deref_1564_store_0_req_0 : boolean;
  signal ptr_deref_1564_store_0_ack_0 : boolean;
  signal ptr_deref_1564_base_resize_req_0 : boolean;
  signal ptr_deref_1564_addr_0_ack_0 : boolean;
  signal ptr_deref_1564_addr_2_req_1 : boolean;
  signal ptr_deref_1150_base_resize_req_0 : boolean;
  signal ptr_deref_1150_base_resize_ack_0 : boolean;
  signal ptr_deref_1150_root_address_inst_req_0 : boolean;
  signal ptr_deref_1150_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1150_addr_0_req_0 : boolean;
  signal ptr_deref_1150_addr_0_ack_0 : boolean;
  signal ptr_deref_1150_addr_0_req_1 : boolean;
  signal ptr_deref_1150_addr_0_ack_1 : boolean;
  signal ptr_deref_1150_addr_1_req_0 : boolean;
  signal ptr_deref_1150_addr_1_ack_0 : boolean;
  signal ptr_deref_1150_addr_1_req_1 : boolean;
  signal ptr_deref_1150_addr_1_ack_1 : boolean;
  signal ptr_deref_1150_addr_2_req_0 : boolean;
  signal ptr_deref_1150_addr_2_ack_0 : boolean;
  signal ptr_deref_1150_addr_2_req_1 : boolean;
  signal ptr_deref_1150_addr_2_ack_1 : boolean;
  signal ptr_deref_1150_addr_3_req_0 : boolean;
  signal ptr_deref_1150_addr_3_ack_0 : boolean;
  signal ptr_deref_1150_addr_3_req_1 : boolean;
  signal ptr_deref_1150_addr_3_ack_1 : boolean;
  signal binary_1358_inst_req_0 : boolean;
  signal binary_1358_inst_ack_0 : boolean;
  signal type_cast_1429_inst_req_0 : boolean;
  signal binary_1358_inst_req_1 : boolean;
  signal type_cast_1429_inst_ack_0 : boolean;
  signal binary_1358_inst_ack_1 : boolean;
  signal phi_stmt_1334_ack_0 : boolean;
  signal phi_stmt_1341_ack_0 : boolean;
  signal phi_stmt_1426_req_0 : boolean;
  signal binary_1364_inst_req_0 : boolean;
  signal binary_1364_inst_ack_0 : boolean;
  signal binary_1364_inst_req_1 : boolean;
  signal binary_1364_inst_ack_1 : boolean;
  signal phi_stmt_1426_ack_0 : boolean;
  signal phi_stmt_1433_ack_0 : boolean;
  signal phi_stmt_1439_ack_0 : boolean;
  signal binary_1370_inst_req_0 : boolean;
  signal binary_1370_inst_ack_0 : boolean;
  signal binary_1370_inst_req_1 : boolean;
  signal binary_1370_inst_ack_1 : boolean;
  signal array_obj_ref_1374_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1374_index_0_resize_ack_0 : boolean;
  signal type_cast_1682_inst_req_0 : boolean;
  signal array_obj_ref_1374_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1374_index_0_rename_ack_0 : boolean;
  signal type_cast_1682_inst_ack_0 : boolean;
  signal array_obj_ref_1374_offset_inst_req_0 : boolean;
  signal array_obj_ref_1374_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1374_base_resize_req_0 : boolean;
  signal array_obj_ref_1374_base_resize_ack_0 : boolean;
  signal array_obj_ref_1374_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1374_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1374_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1374_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1374_final_reg_req_0 : boolean;
  signal array_obj_ref_1374_final_reg_ack_0 : boolean;
  signal phi_stmt_1341_req_1 : boolean;
  signal type_cast_1378_inst_req_0 : boolean;
  signal type_cast_1378_inst_ack_0 : boolean;
  signal type_cast_1444_inst_req_0 : boolean;
  signal type_cast_1444_inst_ack_0 : boolean;
  signal phi_stmt_1439_req_1 : boolean;
  signal ptr_deref_1382_base_resize_req_0 : boolean;
  signal ptr_deref_1382_base_resize_ack_0 : boolean;
  signal ptr_deref_1382_root_address_inst_req_0 : boolean;
  signal ptr_deref_1382_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1382_addr_0_req_0 : boolean;
  signal type_cast_1686_inst_req_0 : boolean;
  signal ptr_deref_1382_addr_0_ack_0 : boolean;
  signal ptr_deref_1382_addr_0_req_1 : boolean;
  signal type_cast_1686_inst_ack_0 : boolean;
  signal ptr_deref_1382_addr_0_ack_1 : boolean;
  signal ptr_deref_1382_addr_1_req_0 : boolean;
  signal ptr_deref_1382_addr_1_ack_0 : boolean;
  signal ptr_deref_1382_addr_1_req_1 : boolean;
  signal ptr_deref_1382_addr_1_ack_1 : boolean;
  signal ptr_deref_1382_load_0_req_0 : boolean;
  signal ptr_deref_1382_load_0_ack_0 : boolean;
  signal ptr_deref_1382_load_1_req_0 : boolean;
  signal ptr_deref_1382_load_1_ack_0 : boolean;
  signal ptr_deref_1382_load_0_req_1 : boolean;
  signal ptr_deref_1382_load_0_ack_1 : boolean;
  signal ptr_deref_1382_load_1_req_1 : boolean;
  signal ptr_deref_1382_load_1_ack_1 : boolean;
  signal ptr_deref_1382_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_1684_inst_req_0 : boolean;
  signal ptr_deref_1382_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1684_inst_ack_0 : boolean;
  signal type_cast_1438_inst_req_0 : boolean;
  signal type_cast_1438_inst_ack_0 : boolean;
  signal type_cast_1386_inst_req_0 : boolean;
  signal type_cast_1386_inst_ack_0 : boolean;
  signal type_cast_1479_inst_req_0 : boolean;
  signal phi_stmt_1433_req_1 : boolean;
  signal type_cast_1479_inst_ack_0 : boolean;
  signal binary_1391_inst_req_0 : boolean;
  signal binary_1391_inst_ack_0 : boolean;
  signal binary_1391_inst_req_1 : boolean;
  signal phi_stmt_1474_req_1 : boolean;
  signal binary_1391_inst_ack_1 : boolean;
  signal type_cast_1395_inst_req_0 : boolean;
  signal type_cast_1395_inst_ack_0 : boolean;
  signal binary_1399_inst_req_0 : boolean;
  signal binary_1399_inst_ack_0 : boolean;
  signal binary_1399_inst_req_1 : boolean;
  signal binary_1399_inst_ack_1 : boolean;
  signal phi_stmt_1426_req_1 : boolean;
  signal binary_1405_inst_req_0 : boolean;
  signal binary_1405_inst_ack_0 : boolean;
  signal binary_1405_inst_req_1 : boolean;
  signal binary_1405_inst_ack_1 : boolean;
  signal phi_stmt_1433_req_0 : boolean;
  signal if_stmt_1407_branch_req_0 : boolean;
  signal if_stmt_1407_branch_ack_1 : boolean;
  signal if_stmt_1407_branch_ack_0 : boolean;
  signal type_cast_1477_inst_req_0 : boolean;
  signal binary_1418_inst_req_0 : boolean;
  signal type_cast_1477_inst_ack_0 : boolean;
  signal binary_1418_inst_ack_0 : boolean;
  signal binary_1418_inst_req_1 : boolean;
  signal binary_1418_inst_ack_1 : boolean;
  signal type_cast_1442_inst_req_0 : boolean;
  signal type_cast_1442_inst_ack_0 : boolean;
  signal array_obj_ref_1422_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1422_index_0_resize_ack_0 : boolean;
  signal phi_stmt_1474_req_0 : boolean;
  signal array_obj_ref_1422_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1422_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1422_offset_inst_req_0 : boolean;
  signal array_obj_ref_1422_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1422_base_resize_req_0 : boolean;
  signal array_obj_ref_1422_base_resize_ack_0 : boolean;
  signal phi_stmt_1439_req_0 : boolean;
  signal array_obj_ref_1422_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1422_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1422_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1422_root_address_inst_ack_1 : boolean;
  signal phi_stmt_1474_ack_0 : boolean;
  signal array_obj_ref_1422_final_reg_req_0 : boolean;
  signal array_obj_ref_1422_final_reg_ack_0 : boolean;
  signal binary_1450_inst_req_0 : boolean;
  signal binary_1450_inst_ack_0 : boolean;
  signal binary_1450_inst_req_1 : boolean;
  signal binary_1450_inst_ack_1 : boolean;
  signal if_stmt_1452_branch_req_0 : boolean;
  signal if_stmt_1452_branch_ack_1 : boolean;
  signal if_stmt_1452_branch_ack_0 : boolean;
  signal ptr_deref_1461_base_resize_req_0 : boolean;
  signal ptr_deref_1461_base_resize_ack_0 : boolean;
  signal ptr_deref_1461_root_address_inst_req_0 : boolean;
  signal ptr_deref_1461_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1461_addr_0_req_0 : boolean;
  signal ptr_deref_1461_addr_0_ack_0 : boolean;
  signal ptr_deref_1461_load_0_req_0 : boolean;
  signal ptr_deref_1461_load_0_ack_0 : boolean;
  signal ptr_deref_1461_load_0_req_1 : boolean;
  signal ptr_deref_1461_load_0_ack_1 : boolean;
  signal ptr_deref_1461_gather_scatter_req_0 : boolean;
  signal ptr_deref_1461_gather_scatter_ack_0 : boolean;
  signal type_cast_1465_inst_req_0 : boolean;
  signal type_cast_1465_inst_ack_0 : boolean;
  signal binary_1470_inst_req_0 : boolean;
  signal binary_1470_inst_ack_0 : boolean;
  signal binary_1470_inst_req_1 : boolean;
  signal binary_1470_inst_ack_1 : boolean;
  signal binary_1485_inst_req_0 : boolean;
  signal binary_1485_inst_ack_0 : boolean;
  signal binary_1485_inst_req_1 : boolean;
  signal binary_1485_inst_ack_1 : boolean;
  signal binary_1491_inst_req_0 : boolean;
  signal binary_1491_inst_ack_0 : boolean;
  signal binary_1491_inst_req_1 : boolean;
  signal binary_1491_inst_ack_1 : boolean;
  signal binary_1496_inst_req_0 : boolean;
  signal binary_1496_inst_ack_0 : boolean;
  signal binary_1496_inst_req_1 : boolean;
  signal binary_1496_inst_ack_1 : boolean;
  signal binary_1502_inst_req_0 : boolean;
  signal binary_1502_inst_ack_0 : boolean;
  signal binary_1502_inst_req_1 : boolean;
  signal binary_1502_inst_ack_1 : boolean;
  signal binary_1507_inst_req_0 : boolean;
  signal binary_1507_inst_ack_0 : boolean;
  signal binary_1507_inst_req_1 : boolean;
  signal binary_1507_inst_ack_1 : boolean;
  signal type_cast_1511_inst_req_0 : boolean;
  signal type_cast_1511_inst_ack_0 : boolean;
  signal binary_1517_inst_req_0 : boolean;
  signal binary_1517_inst_ack_0 : boolean;
  signal binary_1517_inst_req_1 : boolean;
  signal binary_1517_inst_ack_1 : boolean;
  signal if_stmt_1519_branch_req_0 : boolean;
  signal if_stmt_1519_branch_ack_1 : boolean;
  signal if_stmt_1519_branch_ack_0 : boolean;
  signal binary_1530_inst_req_0 : boolean;
  signal binary_1530_inst_ack_0 : boolean;
  signal binary_1530_inst_req_1 : boolean;
  signal binary_1530_inst_ack_1 : boolean;
  signal simple_obj_ref_1527_inst_req_0 : boolean;
  signal simple_obj_ref_1527_inst_ack_0 : boolean;
  signal array_obj_ref_1540_base_resize_req_0 : boolean;
  signal array_obj_ref_1540_base_resize_ack_0 : boolean;
  signal array_obj_ref_1540_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1540_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1540_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1540_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1540_final_reg_req_0 : boolean;
  signal array_obj_ref_1540_final_reg_ack_0 : boolean;
  signal ptr_deref_1543_base_resize_req_0 : boolean;
  signal ptr_deref_1543_base_resize_ack_0 : boolean;
  signal ptr_deref_1543_root_address_inst_req_0 : boolean;
  signal ptr_deref_1543_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1543_addr_0_req_0 : boolean;
  signal ptr_deref_1543_addr_0_ack_0 : boolean;
  signal ptr_deref_1543_addr_0_req_1 : boolean;
  signal ptr_deref_1543_addr_0_ack_1 : boolean;
  signal ptr_deref_1543_addr_1_req_0 : boolean;
  signal ptr_deref_1543_addr_1_ack_0 : boolean;
  signal ptr_deref_1543_addr_1_req_1 : boolean;
  signal ptr_deref_1543_addr_1_ack_1 : boolean;
  signal ptr_deref_1543_addr_2_req_0 : boolean;
  signal ptr_deref_1543_addr_2_ack_0 : boolean;
  signal ptr_deref_1543_addr_2_req_1 : boolean;
  signal ptr_deref_1543_addr_2_ack_1 : boolean;
  signal ptr_deref_1543_addr_3_req_0 : boolean;
  signal ptr_deref_1543_addr_3_ack_0 : boolean;
  signal ptr_deref_1543_addr_3_req_1 : boolean;
  signal ptr_deref_1543_addr_3_ack_1 : boolean;
  signal ptr_deref_1543_gather_scatter_req_0 : boolean;
  signal ptr_deref_1543_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1543_store_0_req_0 : boolean;
  signal ptr_deref_1543_store_0_ack_0 : boolean;
  signal ptr_deref_1543_store_1_req_0 : boolean;
  signal ptr_deref_1543_store_1_ack_0 : boolean;
  signal ptr_deref_1543_store_2_req_0 : boolean;
  signal ptr_deref_1543_store_2_ack_0 : boolean;
  signal ptr_deref_1543_store_3_req_0 : boolean;
  signal ptr_deref_1543_store_3_ack_0 : boolean;
  signal ptr_deref_1543_store_0_req_1 : boolean;
  signal ptr_deref_1543_store_0_ack_1 : boolean;
  signal ptr_deref_1543_store_1_req_1 : boolean;
  signal ptr_deref_1543_store_1_ack_1 : boolean;
  signal ptr_deref_1543_store_2_req_1 : boolean;
  signal ptr_deref_1543_store_2_ack_1 : boolean;
  signal ptr_deref_1543_store_3_req_1 : boolean;
  signal ptr_deref_1543_store_3_ack_1 : boolean;
  signal binary_1550_inst_req_0 : boolean;
  signal binary_1550_inst_ack_0 : boolean;
  signal binary_1550_inst_req_1 : boolean;
  signal binary_1550_inst_ack_1 : boolean;
  signal array_obj_ref_1554_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1554_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1554_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1554_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1554_offset_inst_req_0 : boolean;
  signal array_obj_ref_1554_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1554_base_resize_req_0 : boolean;
  signal array_obj_ref_1554_base_resize_ack_0 : boolean;
  signal array_obj_ref_1554_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1554_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1554_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1554_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1554_final_reg_req_0 : boolean;
  signal array_obj_ref_1554_final_reg_ack_0 : boolean;
  signal array_obj_ref_1561_base_resize_req_0 : boolean;
  signal array_obj_ref_1561_base_resize_ack_0 : boolean;
  signal array_obj_ref_1561_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1561_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1561_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1561_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1561_final_reg_req_0 : boolean;
  signal array_obj_ref_1561_final_reg_ack_0 : boolean;
  signal type_cast_1347_inst_ack_0 : boolean;
  signal ptr_deref_1564_store_0_req_1 : boolean;
  signal ptr_deref_1564_store_0_ack_1 : boolean;
  signal ptr_deref_1564_store_1_req_1 : boolean;
  signal ptr_deref_1564_store_1_ack_1 : boolean;
  signal ptr_deref_1564_store_2_req_1 : boolean;
  signal ptr_deref_1564_store_2_ack_1 : boolean;
  signal ptr_deref_1564_store_3_req_1 : boolean;
  signal ptr_deref_1564_store_3_ack_1 : boolean;
  signal binary_1570_inst_req_0 : boolean;
  signal binary_1570_inst_ack_0 : boolean;
  signal binary_1570_inst_req_1 : boolean;
  signal binary_1570_inst_ack_1 : boolean;
  signal if_stmt_1572_branch_req_0 : boolean;
  signal if_stmt_1572_branch_ack_1 : boolean;
  signal if_stmt_1572_branch_ack_0 : boolean;
  signal binary_1582_inst_req_0 : boolean;
  signal binary_1582_inst_ack_0 : boolean;
  signal binary_1582_inst_req_1 : boolean;
  signal binary_1582_inst_ack_1 : boolean;
  signal binary_1587_inst_req_0 : boolean;
  signal binary_1587_inst_ack_0 : boolean;
  signal binary_1587_inst_req_1 : boolean;
  signal binary_1587_inst_ack_1 : boolean;
  signal ternary_1593_inst_req_0 : boolean;
  signal ternary_1593_inst_ack_0 : boolean;
  signal binary_1599_inst_req_0 : boolean;
  signal binary_1599_inst_ack_0 : boolean;
  signal binary_1599_inst_req_1 : boolean;
  signal binary_1599_inst_ack_1 : boolean;
  signal array_obj_ref_1603_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1603_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1603_index_0_rename_req_0 : boolean;
  signal array_obj_ref_1603_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_1603_offset_inst_req_0 : boolean;
  signal array_obj_ref_1603_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1603_base_resize_req_0 : boolean;
  signal array_obj_ref_1603_base_resize_ack_0 : boolean;
  signal array_obj_ref_1603_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1603_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1603_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1603_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1603_final_reg_req_0 : boolean;
  signal array_obj_ref_1603_final_reg_ack_0 : boolean;
  signal ptr_deref_1606_base_resize_req_0 : boolean;
  signal ptr_deref_1606_base_resize_ack_0 : boolean;
  signal ptr_deref_1606_root_address_inst_req_0 : boolean;
  signal ptr_deref_1606_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1606_addr_0_req_0 : boolean;
  signal ptr_deref_1606_addr_0_ack_0 : boolean;
  signal ptr_deref_1606_addr_0_req_1 : boolean;
  signal ptr_deref_1606_addr_0_ack_1 : boolean;
  signal ptr_deref_1606_addr_1_req_0 : boolean;
  signal ptr_deref_1606_addr_1_ack_0 : boolean;
  signal ptr_deref_1606_addr_1_req_1 : boolean;
  signal ptr_deref_1606_addr_1_ack_1 : boolean;
  signal ptr_deref_1606_addr_2_req_0 : boolean;
  signal ptr_deref_1606_addr_2_ack_0 : boolean;
  signal ptr_deref_1606_addr_2_req_1 : boolean;
  signal ptr_deref_1606_addr_2_ack_1 : boolean;
  signal ptr_deref_1606_addr_3_req_0 : boolean;
  signal ptr_deref_1606_addr_3_ack_0 : boolean;
  signal ptr_deref_1606_addr_3_req_1 : boolean;
  signal ptr_deref_1606_addr_3_ack_1 : boolean;
  signal ptr_deref_1606_gather_scatter_req_0 : boolean;
  signal ptr_deref_1606_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1606_store_0_req_0 : boolean;
  signal ptr_deref_1606_store_0_ack_0 : boolean;
  signal ptr_deref_1606_store_1_req_0 : boolean;
  signal ptr_deref_1606_store_1_ack_0 : boolean;
  signal ptr_deref_1606_store_2_req_0 : boolean;
  signal ptr_deref_1606_store_2_ack_0 : boolean;
  signal ptr_deref_1606_store_3_req_0 : boolean;
  signal ptr_deref_1606_store_3_ack_0 : boolean;
  signal ptr_deref_1606_store_0_req_1 : boolean;
  signal ptr_deref_1606_store_0_ack_1 : boolean;
  signal ptr_deref_1606_store_1_req_1 : boolean;
  signal ptr_deref_1606_store_1_ack_1 : boolean;
  signal ptr_deref_1606_store_2_req_1 : boolean;
  signal ptr_deref_1606_store_2_ack_1 : boolean;
  signal ptr_deref_1606_store_3_req_1 : boolean;
  signal ptr_deref_1606_store_3_ack_1 : boolean;
  signal array_obj_ref_1612_base_resize_req_0 : boolean;
  signal array_obj_ref_1612_base_resize_ack_0 : boolean;
  signal array_obj_ref_1612_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1612_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1612_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1612_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1612_final_reg_req_0 : boolean;
  signal array_obj_ref_1612_final_reg_ack_0 : boolean;
  signal type_cast_1616_inst_req_0 : boolean;
  signal type_cast_1616_inst_ack_0 : boolean;
  signal ptr_deref_1620_base_resize_req_0 : boolean;
  signal ptr_deref_1620_base_resize_ack_0 : boolean;
  signal ptr_deref_1620_root_address_inst_req_0 : boolean;
  signal ptr_deref_1620_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1620_addr_0_req_0 : boolean;
  signal ptr_deref_1620_addr_0_ack_0 : boolean;
  signal ptr_deref_1620_addr_0_req_1 : boolean;
  signal ptr_deref_1620_addr_0_ack_1 : boolean;
  signal ptr_deref_1620_addr_1_req_0 : boolean;
  signal ptr_deref_1620_addr_1_ack_0 : boolean;
  signal ptr_deref_1620_addr_1_req_1 : boolean;
  signal ptr_deref_1620_addr_1_ack_1 : boolean;
  signal ptr_deref_1620_addr_2_req_0 : boolean;
  signal ptr_deref_1620_addr_2_ack_0 : boolean;
  signal ptr_deref_1620_addr_2_req_1 : boolean;
  signal ptr_deref_1620_addr_2_ack_1 : boolean;
  signal ptr_deref_1620_addr_3_req_0 : boolean;
  signal ptr_deref_1620_addr_3_ack_0 : boolean;
  signal ptr_deref_1620_addr_3_req_1 : boolean;
  signal ptr_deref_1620_addr_3_ack_1 : boolean;
  signal ptr_deref_1620_load_0_req_0 : boolean;
  signal ptr_deref_1620_load_0_ack_0 : boolean;
  signal ptr_deref_1620_load_1_req_0 : boolean;
  signal ptr_deref_1620_load_1_ack_0 : boolean;
  signal ptr_deref_1620_load_2_req_0 : boolean;
  signal ptr_deref_1620_load_2_ack_0 : boolean;
  signal ptr_deref_1620_load_3_req_0 : boolean;
  signal ptr_deref_1620_load_3_ack_0 : boolean;
  signal ptr_deref_1620_load_0_req_1 : boolean;
  signal ptr_deref_1620_load_0_ack_1 : boolean;
  signal ptr_deref_1620_load_1_req_1 : boolean;
  signal ptr_deref_1620_load_1_ack_1 : boolean;
  signal ptr_deref_1620_load_2_req_1 : boolean;
  signal ptr_deref_1620_load_2_ack_1 : boolean;
  signal ptr_deref_1620_load_3_req_1 : boolean;
  signal ptr_deref_1620_load_3_ack_1 : boolean;
  signal ptr_deref_1620_gather_scatter_req_0 : boolean;
  signal ptr_deref_1620_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1627_base_resize_req_0 : boolean;
  signal array_obj_ref_1627_base_resize_ack_0 : boolean;
  signal array_obj_ref_1627_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1627_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1627_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1627_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1627_final_reg_req_0 : boolean;
  signal array_obj_ref_1627_final_reg_ack_0 : boolean;
  signal type_cast_1631_inst_req_0 : boolean;
  signal type_cast_1631_inst_ack_0 : boolean;
  signal ptr_deref_1634_base_resize_req_0 : boolean;
  signal ptr_deref_1634_base_resize_ack_0 : boolean;
  signal ptr_deref_1634_root_address_inst_req_0 : boolean;
  signal ptr_deref_1634_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1634_addr_0_req_0 : boolean;
  signal ptr_deref_1634_addr_0_ack_0 : boolean;
  signal ptr_deref_1634_addr_0_req_1 : boolean;
  signal ptr_deref_1634_addr_0_ack_1 : boolean;
  signal ptr_deref_1634_addr_1_req_0 : boolean;
  signal ptr_deref_1634_addr_1_ack_0 : boolean;
  signal ptr_deref_1634_addr_1_req_1 : boolean;
  signal ptr_deref_1634_addr_1_ack_1 : boolean;
  signal ptr_deref_1634_addr_2_req_0 : boolean;
  signal ptr_deref_1634_addr_2_ack_0 : boolean;
  signal ptr_deref_1634_addr_2_req_1 : boolean;
  signal ptr_deref_1634_addr_2_ack_1 : boolean;
  signal ptr_deref_1634_addr_3_req_0 : boolean;
  signal ptr_deref_1634_addr_3_ack_0 : boolean;
  signal ptr_deref_1634_addr_3_req_1 : boolean;
  signal ptr_deref_1634_addr_3_ack_1 : boolean;
  signal ptr_deref_1634_gather_scatter_req_0 : boolean;
  signal ptr_deref_1634_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1634_store_0_req_0 : boolean;
  signal ptr_deref_1634_store_0_ack_0 : boolean;
  signal ptr_deref_1634_store_1_req_0 : boolean;
  signal ptr_deref_1634_store_1_ack_0 : boolean;
  signal ptr_deref_1634_store_2_req_0 : boolean;
  signal ptr_deref_1634_store_2_ack_0 : boolean;
  signal ptr_deref_1634_store_3_req_0 : boolean;
  signal ptr_deref_1634_store_3_ack_0 : boolean;
  signal ptr_deref_1634_store_0_req_1 : boolean;
  signal ptr_deref_1634_store_0_ack_1 : boolean;
  signal ptr_deref_1634_store_1_req_1 : boolean;
  signal ptr_deref_1634_store_1_ack_1 : boolean;
  signal ptr_deref_1634_store_2_req_1 : boolean;
  signal ptr_deref_1634_store_2_ack_1 : boolean;
  signal ptr_deref_1634_store_3_req_1 : boolean;
  signal ptr_deref_1634_store_3_ack_1 : boolean;
  signal array_obj_ref_1642_base_resize_req_0 : boolean;
  signal array_obj_ref_1642_base_resize_ack_0 : boolean;
  signal array_obj_ref_1642_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1642_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1642_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1642_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1642_final_reg_req_0 : boolean;
  signal array_obj_ref_1642_final_reg_ack_0 : boolean;
  signal type_cast_1646_inst_req_0 : boolean;
  signal type_cast_1646_inst_ack_0 : boolean;
  signal ptr_deref_1650_base_resize_req_0 : boolean;
  signal ptr_deref_1650_base_resize_ack_0 : boolean;
  signal ptr_deref_1650_root_address_inst_req_0 : boolean;
  signal ptr_deref_1650_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1650_addr_0_req_0 : boolean;
  signal ptr_deref_1650_addr_0_ack_0 : boolean;
  signal ptr_deref_1650_addr_0_req_1 : boolean;
  signal ptr_deref_1650_addr_0_ack_1 : boolean;
  signal ptr_deref_1650_addr_1_req_0 : boolean;
  signal ptr_deref_1650_addr_1_ack_0 : boolean;
  signal ptr_deref_1650_addr_1_req_1 : boolean;
  signal ptr_deref_1650_addr_1_ack_1 : boolean;
  signal ptr_deref_1650_addr_2_req_0 : boolean;
  signal ptr_deref_1650_addr_2_ack_0 : boolean;
  signal ptr_deref_1650_addr_2_req_1 : boolean;
  signal ptr_deref_1650_addr_2_ack_1 : boolean;
  signal ptr_deref_1650_addr_3_req_0 : boolean;
  signal ptr_deref_1650_addr_3_ack_0 : boolean;
  signal ptr_deref_1650_addr_3_req_1 : boolean;
  signal ptr_deref_1650_addr_3_ack_1 : boolean;
  signal ptr_deref_1650_load_0_req_0 : boolean;
  signal ptr_deref_1650_load_0_ack_0 : boolean;
  signal ptr_deref_1650_load_1_req_0 : boolean;
  signal ptr_deref_1650_load_1_ack_0 : boolean;
  signal ptr_deref_1650_load_2_req_0 : boolean;
  signal ptr_deref_1650_load_2_ack_0 : boolean;
  signal ptr_deref_1650_load_3_req_0 : boolean;
  signal ptr_deref_1650_load_3_ack_0 : boolean;
  signal ptr_deref_1650_load_0_req_1 : boolean;
  signal ptr_deref_1650_load_0_ack_1 : boolean;
  signal ptr_deref_1650_load_1_req_1 : boolean;
  signal ptr_deref_1650_load_1_ack_1 : boolean;
  signal ptr_deref_1650_load_2_req_1 : boolean;
  signal ptr_deref_1650_load_2_ack_1 : boolean;
  signal ptr_deref_1650_load_3_req_1 : boolean;
  signal ptr_deref_1650_load_3_ack_1 : boolean;
  signal ptr_deref_1650_gather_scatter_req_0 : boolean;
  signal ptr_deref_1650_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_1657_base_resize_req_0 : boolean;
  signal array_obj_ref_1657_base_resize_ack_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1657_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1657_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1657_final_reg_req_0 : boolean;
  signal array_obj_ref_1657_final_reg_ack_0 : boolean;
  signal type_cast_1661_inst_req_0 : boolean;
  signal type_cast_1661_inst_ack_0 : boolean;
  signal ptr_deref_1664_base_resize_req_0 : boolean;
  signal ptr_deref_1664_base_resize_ack_0 : boolean;
  signal ptr_deref_1664_root_address_inst_req_0 : boolean;
  signal ptr_deref_1664_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1664_addr_0_req_0 : boolean;
  signal ptr_deref_1664_addr_0_ack_0 : boolean;
  signal ptr_deref_1664_addr_0_req_1 : boolean;
  signal ptr_deref_1664_addr_0_ack_1 : boolean;
  signal ptr_deref_1664_addr_1_req_0 : boolean;
  signal ptr_deref_1664_addr_1_ack_0 : boolean;
  signal ptr_deref_1664_addr_1_req_1 : boolean;
  signal ptr_deref_1664_addr_1_ack_1 : boolean;
  signal ptr_deref_1664_addr_2_req_0 : boolean;
  signal ptr_deref_1664_addr_2_ack_0 : boolean;
  signal ptr_deref_1664_addr_2_req_1 : boolean;
  signal ptr_deref_1664_addr_2_ack_1 : boolean;
  signal ptr_deref_1664_addr_3_req_0 : boolean;
  signal ptr_deref_1664_addr_3_ack_0 : boolean;
  signal ptr_deref_1664_addr_3_req_1 : boolean;
  signal ptr_deref_1664_addr_3_ack_1 : boolean;
  signal ptr_deref_1664_gather_scatter_req_0 : boolean;
  signal ptr_deref_1664_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1664_store_0_req_0 : boolean;
  signal ptr_deref_1664_store_0_ack_0 : boolean;
  signal ptr_deref_1664_store_1_req_0 : boolean;
  signal ptr_deref_1664_store_1_ack_0 : boolean;
  signal ptr_deref_1664_store_2_req_0 : boolean;
  signal ptr_deref_1664_store_2_ack_0 : boolean;
  signal ptr_deref_1664_store_3_req_0 : boolean;
  signal ptr_deref_1664_store_3_ack_0 : boolean;
  signal ptr_deref_1664_store_0_req_1 : boolean;
  signal ptr_deref_1664_store_0_ack_1 : boolean;
  signal ptr_deref_1664_store_1_req_1 : boolean;
  signal ptr_deref_1664_store_1_ack_1 : boolean;
  signal ptr_deref_1664_store_2_req_1 : boolean;
  signal ptr_deref_1664_store_2_ack_1 : boolean;
  signal ptr_deref_1664_store_3_req_1 : boolean;
  signal ptr_deref_1664_store_3_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_chk_1_CP_4158: Block -- control-path 
    signal cp_elements: BooleanArray(979 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(979);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(979), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(141);
    cpelement_group_2 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(898));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(2),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(3) <= cp_elements(213);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(222) & cp_elements(900));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(249) & cp_elements(902));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(287) & cp_elements(904));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(7) <= OrReduce(cp_elements(308) & cp_elements(906));
    cp_elements(8) <= cp_elements(921);
    cp_elements(9) <= cp_elements(391);
    cp_elements(10) <= OrReduce(cp_elements(400) & cp_elements(923));
    cp_elements(11) <= cp_elements(956);
    cp_elements(12) <= OrReduce(cp_elements(430) & cp_elements(958));
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(489) & cp_elements(971));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(14) <= cp_elements(606);
    cp_elements(15) <= OrReduce(cp_elements(613) & cp_elements(973));
    cp_elements(16) <= cp_elements(779);
    cp_elements(17) <= cp_elements(876);
    cp_elements(18) <= OrReduce(cp_elements(975) & cp_elements(977));
    cp_elements(19) <= cp_elements(0);
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(21) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4290_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_1119_inst_req_0); -- 
    cp_elements(21) <= cp_elements(19);
    cp_elements(22) <= cp_elements(19);
    req_4285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => simple_obj_ref_1118_inst_req_0); -- 
    ack_4286_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1118_inst_ack_0, ack => cp_elements(23)); -- 
    ack_4291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1119_inst_ack_0, ack => cp_elements(24)); -- 
    cp_elements(25) <= cp_elements(24);
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(27));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4303_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => type_cast_1123_inst_req_0); -- 
    cp_elements(27) <= cp_elements(25);
    cp_elements(28) <= cp_elements(25);
    cp_elements(29) <= type_cast_1123_inst_ack_0;
    cp_elements(30) <= cp_elements(25);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_1130_final_reg_req_0); -- 
    cp_elements(32) <= cp_elements(29);
    base_resize_req_4315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => array_obj_ref_1130_base_resize_req_0); -- 
    base_resize_ack_4316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_base_resize_ack_0, ack => cp_elements(33)); -- 
    plus_base_rr_4321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => array_obj_ref_1130_root_address_inst_req_0); -- 
    plus_base_ra_4322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_root_address_inst_ack_0, ack => cp_elements(34)); -- 
    plus_base_cr_4323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_1130_root_address_inst_req_1); -- 
    plus_base_ca_4324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_root_address_inst_ack_1, ack => cp_elements(35)); -- 
    final_reg_ack_4329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1130_final_reg_ack_0, ack => cp_elements(36)); -- 
    base_resize_req_4342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_1134_base_resize_req_0); -- 
    base_resize_ack_4343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_base_resize_ack_0, ack => cp_elements(37)); -- 
    sum_rename_req_4347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_1134_root_address_inst_req_0); -- 
    cp_elements(38) <= ptr_deref_1134_root_address_inst_ack_0;
    cp_elements(39) <= cp_elements(38);
    rr_4355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => ptr_deref_1134_addr_0_req_0); -- 
    ra_4356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_0_ack_0, ack => cp_elements(40)); -- 
    cr_4357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_1134_addr_0_req_1); -- 
    ca_4358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_0_ack_1, ack => cp_elements(41)); -- 
    cp_elements(42) <= cp_elements(38);
    rr_4362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_1134_addr_1_req_0); -- 
    ra_4363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_1_ack_0, ack => cp_elements(43)); -- 
    cr_4364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_1134_addr_1_req_1); -- 
    ca_4365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_1_ack_1, ack => cp_elements(44)); -- 
    cp_elements(45) <= cp_elements(38);
    rr_4369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_1134_addr_2_req_0); -- 
    ra_4370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_2_ack_0, ack => cp_elements(46)); -- 
    cr_4371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_1134_addr_2_req_1); -- 
    ca_4372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_2_ack_1, ack => cp_elements(47)); -- 
    cp_elements(48) <= cp_elements(38);
    rr_4376_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_1134_addr_3_req_0); -- 
    ra_4377_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_3_ack_0, ack => cp_elements(49)); -- 
    cr_4378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_1134_addr_3_req_1); -- 
    ca_4379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_addr_3_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(41) & cp_elements(44) & cp_elements(47) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(52) <= cp_elements(51);
    rr_4389_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_1134_load_0_req_0); -- 
    ra_4390_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_0_ack_0, ack => cp_elements(53)); -- 
    cp_elements(54) <= cp_elements(51);
    rr_4394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_1134_load_1_req_0); -- 
    ra_4395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_1_ack_0, ack => cp_elements(55)); -- 
    cp_elements(56) <= cp_elements(51);
    rr_4399_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_1134_load_2_req_0); -- 
    ra_4400_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_2_ack_0, ack => cp_elements(57)); -- 
    cp_elements(58) <= cp_elements(51);
    rr_4404_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_1134_load_3_req_0); -- 
    ra_4405_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_3_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(55) & cp_elements(57) & cp_elements(59));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(61) <= cp_elements(60);
    cr_4415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_1134_load_0_req_1); -- 
    ca_4416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_0_ack_1, ack => cp_elements(62)); -- 
    cp_elements(63) <= cp_elements(60);
    cr_4420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_1134_load_1_req_1); -- 
    ca_4421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_1_ack_1, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(60);
    cr_4425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_1134_load_2_req_1); -- 
    ca_4426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_2_ack_1, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(60);
    cr_4430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_1134_load_3_req_1); -- 
    ca_4431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1134_load_3_ack_1, ack => cp_elements(68)); -- 
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(62) & cp_elements(64) & cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_4432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_1134_gather_scatter_req_0); -- 
    cp_elements(70) <= ptr_deref_1134_gather_scatter_ack_0;
    cp_elements(71) <= cp_elements(25);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_1139_final_reg_req_0); -- 
    cp_elements(73) <= cp_elements(70);
    base_resize_req_4444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_1139_base_resize_req_0); -- 
    base_resize_ack_4445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1139_base_resize_ack_0, ack => cp_elements(74)); -- 
    plus_base_rr_4450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_1139_root_address_inst_req_0); -- 
    plus_base_ra_4451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1139_root_address_inst_ack_0, ack => cp_elements(75)); -- 
    plus_base_cr_4452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_1139_root_address_inst_req_1); -- 
    plus_base_ca_4453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1139_root_address_inst_ack_1, ack => cp_elements(76)); -- 
    final_reg_ack_4458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1139_final_reg_ack_0, ack => cp_elements(77)); -- 
    cp_elements(78) <= cp_elements(25);
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(83));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => array_obj_ref_1146_final_reg_req_0); -- 
    cp_elements(80) <= cp_elements(29);
    base_resize_req_4469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => array_obj_ref_1146_base_resize_req_0); -- 
    base_resize_ack_4470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1146_base_resize_ack_0, ack => cp_elements(81)); -- 
    plus_base_rr_4475_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_1146_root_address_inst_req_0); -- 
    plus_base_ra_4476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1146_root_address_inst_ack_0, ack => cp_elements(82)); -- 
    plus_base_cr_4477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_1146_root_address_inst_req_1); -- 
    plus_base_ca_4478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1146_root_address_inst_ack_1, ack => cp_elements(83)); -- 
    final_reg_ack_4483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1146_final_reg_ack_0, ack => cp_elements(84)); -- 
    base_resize_req_4496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_1150_base_resize_req_0); -- 
    base_resize_ack_4497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_base_resize_ack_0, ack => cp_elements(85)); -- 
    sum_rename_req_4501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_1150_root_address_inst_req_0); -- 
    cp_elements(86) <= ptr_deref_1150_root_address_inst_ack_0;
    cp_elements(87) <= cp_elements(86);
    rr_4509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => ptr_deref_1150_addr_0_req_0); -- 
    ra_4510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_0_ack_0, ack => cp_elements(88)); -- 
    cr_4511_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_1150_addr_0_req_1); -- 
    ca_4512_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_0_ack_1, ack => cp_elements(89)); -- 
    cp_elements(90) <= cp_elements(86);
    rr_4516_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => ptr_deref_1150_addr_1_req_0); -- 
    ra_4517_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_1_ack_0, ack => cp_elements(91)); -- 
    cr_4518_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => ptr_deref_1150_addr_1_req_1); -- 
    ca_4519_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_1_ack_1, ack => cp_elements(92)); -- 
    cp_elements(93) <= cp_elements(86);
    rr_4523_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_1150_addr_2_req_0); -- 
    ra_4524_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_2_ack_0, ack => cp_elements(94)); -- 
    cr_4525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_1150_addr_2_req_1); -- 
    ca_4526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_2_ack_1, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(86);
    rr_4530_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_1150_addr_3_req_0); -- 
    ra_4531_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_3_ack_0, ack => cp_elements(97)); -- 
    cr_4532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_1150_addr_3_req_1); -- 
    ca_4533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_addr_3_ack_1, ack => cp_elements(98)); -- 
    cpelement_group_99 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(92) & cp_elements(95) & cp_elements(98));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(99),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(100) <= cp_elements(99);
    rr_4543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_1150_load_0_req_0); -- 
    ra_4544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_0_ack_0, ack => cp_elements(101)); -- 
    cp_elements(102) <= cp_elements(99);
    rr_4548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => ptr_deref_1150_load_1_req_0); -- 
    ra_4549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_1_ack_0, ack => cp_elements(103)); -- 
    cp_elements(104) <= cp_elements(99);
    rr_4553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_1150_load_2_req_0); -- 
    ra_4554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_2_ack_0, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(99);
    rr_4558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_1150_load_3_req_0); -- 
    ra_4559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_3_ack_0, ack => cp_elements(107)); -- 
    cpelement_group_108 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(101) & cp_elements(103) & cp_elements(105) & cp_elements(107));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(108),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(109) <= cp_elements(108);
    cr_4569_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_1150_load_0_req_1); -- 
    ca_4570_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_0_ack_1, ack => cp_elements(110)); -- 
    cp_elements(111) <= cp_elements(108);
    cr_4574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_1150_load_1_req_1); -- 
    ca_4575_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_1_ack_1, ack => cp_elements(112)); -- 
    cp_elements(113) <= cp_elements(108);
    cr_4579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_1150_load_2_req_1); -- 
    ca_4580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_2_ack_1, ack => cp_elements(114)); -- 
    cp_elements(115) <= cp_elements(108);
    cr_4584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_1150_load_3_req_1); -- 
    ca_4585_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_load_3_ack_1, ack => cp_elements(116)); -- 
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112) & cp_elements(114) & cp_elements(116));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_4586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_1150_gather_scatter_req_0); -- 
    merge_ack_4587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1150_gather_scatter_ack_0, ack => cp_elements(118)); -- 
    cpelement_group_119 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(120));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(119),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => type_cast_1154_inst_req_0); -- 
    cp_elements(120) <= cp_elements(25);
    ack_4597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1154_inst_ack_0, ack => cp_elements(121)); -- 
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(124));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => type_cast_1158_inst_req_0); -- 
    cp_elements(123) <= cp_elements(25);
    cp_elements(124) <= cp_elements(70);
    ack_4607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1158_inst_ack_0, ack => cp_elements(125)); -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(121) & cp_elements(125) & cp_elements(127));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => binary_1163_inst_req_0); -- 
    cp_elements(127) <= cp_elements(25);
    ra_4618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1163_inst_ack_0, ack => cp_elements(128)); -- 
    cr_4619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => binary_1163_inst_req_1); -- 
    ca_4620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1163_inst_ack_1, ack => cp_elements(129)); -- 
    cpelement_group_130 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(129) & cp_elements(131));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => binary_1169_inst_req_0); -- 
    cp_elements(131) <= cp_elements(25);
    ra_4630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1169_inst_ack_0, ack => cp_elements(132)); -- 
    cr_4631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => binary_1169_inst_req_1); -- 
    ca_4632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1169_inst_ack_1, ack => cp_elements(133)); -- 
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(135) & cp_elements(138));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => binary_1177_inst_req_0); -- 
    cp_elements(135) <= cp_elements(25);
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => type_cast_1173_inst_req_0); -- 
    cp_elements(137) <= cp_elements(25);
    ack_4644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1173_inst_ack_0, ack => cp_elements(138)); -- 
    ra_4649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1177_inst_ack_0, ack => cp_elements(139)); -- 
    cr_4650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => binary_1177_inst_req_1); -- 
    ca_4651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1177_inst_ack_1, ack => cp_elements(140)); -- 
    cpelement_group_141 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(77) & cp_elements(140));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(141),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(142) <= cp_elements(1);
    cp_elements(143) <= false;
    cp_elements(144) <= cp_elements(143);
    cp_elements(145) <= cp_elements(1);
    branch_req_4659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => if_stmt_1179_branch_req_0); -- 
    cp_elements(146) <= cp_elements(145);
    cp_elements(147) <= cp_elements(146);
    if_choice_transition_4664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1179_branch_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    else_choice_transition_4668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1179_branch_ack_0, ack => cp_elements(150)); -- 
    cpelement_group_151 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(152) & cp_elements(153));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(151),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => binary_1190_inst_req_0); -- 
    cp_elements(152) <= cp_elements(2);
    cp_elements(153) <= cp_elements(2);
    ra_4686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1190_inst_ack_0, ack => cp_elements(154)); -- 
    cr_4687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => binary_1190_inst_req_1); -- 
    ca_4688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1190_inst_ack_1, ack => cp_elements(155)); -- 
    pipe_wreq_4693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => simple_obj_ref_1187_inst_req_0); -- 
    pipe_wack_4694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1187_inst_ack_0, ack => cp_elements(156)); -- 
    cp_elements(157) <= cp_elements(150);
    cpelement_group_158 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(159) & cp_elements(160));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => type_cast_1197_inst_req_0); -- 
    cp_elements(159) <= cp_elements(157);
    cp_elements(160) <= cp_elements(157);
    ack_4707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1197_inst_ack_0, ack => cp_elements(161)); -- 
    base_resize_req_4720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => ptr_deref_1201_base_resize_req_0); -- 
    base_resize_ack_4721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_base_resize_ack_0, ack => cp_elements(162)); -- 
    sum_rename_req_4725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => ptr_deref_1201_root_address_inst_req_0); -- 
    cp_elements(163) <= ptr_deref_1201_root_address_inst_ack_0;
    cp_elements(164) <= cp_elements(163);
    rr_4733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => ptr_deref_1201_addr_0_req_0); -- 
    ra_4734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_0_ack_0, ack => cp_elements(165)); -- 
    cr_4735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => ptr_deref_1201_addr_0_req_1); -- 
    ca_4736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_0_ack_1, ack => cp_elements(166)); -- 
    cp_elements(167) <= cp_elements(163);
    rr_4740_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => ptr_deref_1201_addr_1_req_0); -- 
    ra_4741_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_1_ack_0, ack => cp_elements(168)); -- 
    cr_4742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => ptr_deref_1201_addr_1_req_1); -- 
    ca_4743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_1_ack_1, ack => cp_elements(169)); -- 
    cp_elements(170) <= cp_elements(163);
    rr_4747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => ptr_deref_1201_addr_2_req_0); -- 
    ra_4748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_2_ack_0, ack => cp_elements(171)); -- 
    cr_4749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => ptr_deref_1201_addr_2_req_1); -- 
    ca_4750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_2_ack_1, ack => cp_elements(172)); -- 
    cp_elements(173) <= cp_elements(163);
    rr_4754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => ptr_deref_1201_addr_3_req_0); -- 
    ra_4755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_3_ack_0, ack => cp_elements(174)); -- 
    cr_4756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(174), ack => ptr_deref_1201_addr_3_req_1); -- 
    ca_4757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_addr_3_ack_1, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(166) & cp_elements(169) & cp_elements(172) & cp_elements(175));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(177) <= cp_elements(176);
    rr_4767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => ptr_deref_1201_load_0_req_0); -- 
    ra_4768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_0_ack_0, ack => cp_elements(178)); -- 
    cp_elements(179) <= cp_elements(176);
    rr_4772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => ptr_deref_1201_load_1_req_0); -- 
    ra_4773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_1_ack_0, ack => cp_elements(180)); -- 
    cp_elements(181) <= cp_elements(176);
    rr_4777_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => ptr_deref_1201_load_2_req_0); -- 
    ra_4778_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_2_ack_0, ack => cp_elements(182)); -- 
    cp_elements(183) <= cp_elements(176);
    rr_4782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => ptr_deref_1201_load_3_req_0); -- 
    ra_4783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_3_ack_0, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(180) & cp_elements(182) & cp_elements(184));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(186) <= cp_elements(185);
    cr_4793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => ptr_deref_1201_load_0_req_1); -- 
    ca_4794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_0_ack_1, ack => cp_elements(187)); -- 
    cp_elements(188) <= cp_elements(185);
    cr_4798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_1201_load_1_req_1); -- 
    ca_4799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_1_ack_1, ack => cp_elements(189)); -- 
    cp_elements(190) <= cp_elements(185);
    cr_4803_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_1201_load_2_req_1); -- 
    ca_4804_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_2_ack_1, ack => cp_elements(191)); -- 
    cp_elements(192) <= cp_elements(185);
    cr_4808_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_1201_load_3_req_1); -- 
    ca_4809_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1201_load_3_ack_1, ack => cp_elements(193)); -- 
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(187) & cp_elements(189) & cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_4810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => ptr_deref_1201_gather_scatter_req_0); -- 
    cp_elements(195) <= ptr_deref_1201_gather_scatter_ack_0;
    cpelement_group_196 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(197) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(196),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => binary_1207_inst_req_0); -- 
    cp_elements(197) <= cp_elements(157);
    cp_elements(198) <= cp_elements(195);
    ra_4821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1207_inst_ack_0, ack => cp_elements(199)); -- 
    cr_4822_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => binary_1207_inst_req_1); -- 
    ca_4823_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1207_inst_ack_1, ack => cp_elements(200)); -- 
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(200) & cp_elements(202));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => binary_1213_inst_req_0); -- 
    cp_elements(202) <= cp_elements(157);
    ra_4833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1213_inst_ack_0, ack => cp_elements(203)); -- 
    cr_4834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => binary_1213_inst_req_1); -- 
    ca_4835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1213_inst_ack_1, ack => cp_elements(204)); -- 
    cpelement_group_205 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(206) & cp_elements(207));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(205),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4844_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => binary_1219_inst_req_0); -- 
    cp_elements(206) <= cp_elements(157);
    cp_elements(207) <= cp_elements(195);
    ra_4845_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1219_inst_ack_0, ack => cp_elements(208)); -- 
    cr_4846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => binary_1219_inst_req_1); -- 
    ca_4847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1219_inst_ack_1, ack => cp_elements(209)); -- 
    cpelement_group_210 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(209) & cp_elements(211));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(210),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_4856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => type_cast_1223_inst_req_0); -- 
    cp_elements(211) <= cp_elements(157);
    ack_4857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1223_inst_ack_0, ack => cp_elements(212)); -- 
    cpelement_group_213 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(204) & cp_elements(212));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(213),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(214) <= cp_elements(3);
    cp_elements(215) <= false;
    cp_elements(216) <= cp_elements(215);
    cp_elements(217) <= cp_elements(3);
    branch_req_4865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => if_stmt_1225_branch_req_0); -- 
    cp_elements(218) <= cp_elements(217);
    cp_elements(219) <= cp_elements(218);
    if_choice_transition_4870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1225_branch_ack_1, ack => cp_elements(220)); -- 
    cp_elements(221) <= cp_elements(218);
    else_choice_transition_4874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1225_branch_ack_0, ack => cp_elements(222)); -- 
    cpelement_group_223 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(224) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(223),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => binary_1236_inst_req_0); -- 
    cp_elements(224) <= cp_elements(4);
    cp_elements(225) <= cp_elements(4);
    ra_4892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1236_inst_ack_0, ack => cp_elements(226)); -- 
    cr_4893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => binary_1236_inst_req_1); -- 
    ca_4894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1236_inst_ack_1, ack => cp_elements(227)); -- 
    pipe_wreq_4899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => simple_obj_ref_1233_inst_req_0); -- 
    pipe_wack_4900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1233_inst_ack_0, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(220);
    cpelement_group_230 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(231) & cp_elements(232));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(230),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4912_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => binary_1245_inst_req_0); -- 
    cp_elements(231) <= cp_elements(229);
    cp_elements(232) <= cp_elements(229);
    ra_4913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1245_inst_ack_0, ack => cp_elements(233)); -- 
    cr_4914_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => binary_1245_inst_req_1); -- 
    ca_4915_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1245_inst_ack_1, ack => cp_elements(234)); -- 
    cpelement_group_235 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(234) & cp_elements(236));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(235),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => binary_1251_inst_req_0); -- 
    cp_elements(236) <= cp_elements(229);
    ra_4925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1251_inst_ack_0, ack => cp_elements(237)); -- 
    cr_4926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => binary_1251_inst_req_1); -- 
    ca_4927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1251_inst_ack_1, ack => cp_elements(238)); -- 
    cpelement_group_239 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(240));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(239),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => binary_1257_inst_req_0); -- 
    cp_elements(240) <= cp_elements(229);
    ra_4937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1257_inst_ack_0, ack => cp_elements(241)); -- 
    cr_4938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => binary_1257_inst_req_1); -- 
    ca_4939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1257_inst_ack_1, ack => cp_elements(242)); -- 
    cp_elements(243) <= cp_elements(242);
    cp_elements(244) <= false;
    cp_elements(245) <= cp_elements(244);
    cp_elements(246) <= cp_elements(242);
    branch_req_4947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => if_stmt_1259_branch_req_0); -- 
    cp_elements(247) <= cp_elements(246);
    cp_elements(248) <= cp_elements(247);
    if_choice_transition_4952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1259_branch_ack_1, ack => cp_elements(249)); -- 
    cp_elements(250) <= cp_elements(247);
    else_choice_transition_4956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1259_branch_ack_0, ack => cp_elements(251)); -- 
    crr_4992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => call_stmt_1277_call_req_0); -- 
    cpelement_group_252 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(253) & cp_elements(254));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(252),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_4973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => binary_1270_inst_req_0); -- 
    cp_elements(253) <= cp_elements(5);
    cp_elements(254) <= cp_elements(5);
    ra_4974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1270_inst_ack_0, ack => cp_elements(255)); -- 
    cr_4975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => binary_1270_inst_req_1); -- 
    ca_4976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1270_inst_ack_1, ack => cp_elements(256)); -- 
    pipe_wreq_4981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => simple_obj_ref_1267_inst_req_0); -- 
    pipe_wack_4982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1267_inst_ack_0, ack => cp_elements(257)); -- 
    cra_4993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1277_call_ack_0, ack => cp_elements(258)); -- 
    ccr_4997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => call_stmt_1277_call_req_1); -- 
    cca_4998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1277_call_ack_1, ack => cp_elements(259)); -- 
    cp_elements(260) <= cp_elements(259);
    cpelement_group_261 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(263));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(261),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5012_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => type_cast_1280_inst_req_0); -- 
    cp_elements(262) <= cp_elements(260);
    cp_elements(263) <= cp_elements(260);
    cp_elements(264) <= type_cast_1280_inst_ack_0;
    cpelement_group_265 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(266) & cp_elements(267) & cp_elements(268));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(265),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => binary_1285_inst_req_0); -- 
    cp_elements(266) <= cp_elements(260);
    cp_elements(267) <= cp_elements(264);
    cp_elements(268) <= cp_elements(260);
    ra_5024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1285_inst_ack_0, ack => cp_elements(269)); -- 
    cr_5025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => binary_1285_inst_req_1); -- 
    ca_5026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1285_inst_ack_1, ack => cp_elements(270)); -- 
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(272) & cp_elements(273) & cp_elements(274));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => binary_1290_inst_req_0); -- 
    cp_elements(272) <= cp_elements(260);
    cp_elements(273) <= cp_elements(264);
    cp_elements(274) <= cp_elements(260);
    ra_5037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1290_inst_ack_0, ack => cp_elements(275)); -- 
    cr_5038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => binary_1290_inst_req_1); -- 
    ca_5039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1290_inst_ack_1, ack => cp_elements(276)); -- 
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(270) & cp_elements(276) & cp_elements(278));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => binary_1295_inst_req_0); -- 
    cp_elements(278) <= cp_elements(260);
    ra_5050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1295_inst_ack_0, ack => cp_elements(279)); -- 
    cr_5051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => binary_1295_inst_req_1); -- 
    ca_5052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1295_inst_ack_1, ack => cp_elements(280)); -- 
    cp_elements(281) <= cp_elements(280);
    cp_elements(282) <= false;
    cp_elements(283) <= cp_elements(282);
    cp_elements(284) <= cp_elements(280);
    branch_req_5060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => if_stmt_1297_branch_req_0); -- 
    cp_elements(285) <= cp_elements(284);
    cp_elements(286) <= cp_elements(285);
    if_choice_transition_5065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1297_branch_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(285);
    else_choice_transition_5069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1297_branch_ack_0, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(292));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => binary_1308_inst_req_0); -- 
    cp_elements(291) <= cp_elements(6);
    cp_elements(292) <= cp_elements(6);
    ra_5087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1308_inst_ack_0, ack => cp_elements(293)); -- 
    cr_5088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => binary_1308_inst_req_1); -- 
    ca_5089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1308_inst_ack_1, ack => cp_elements(294)); -- 
    pipe_wreq_5094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => simple_obj_ref_1305_inst_req_0); -- 
    pipe_wack_5095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1305_inst_ack_0, ack => cp_elements(295)); -- 
    cp_elements(296) <= cp_elements(289);
    cpelement_group_297 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(298) & cp_elements(299));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(297),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => binary_1317_inst_req_0); -- 
    cp_elements(298) <= cp_elements(296);
    cp_elements(299) <= cp_elements(296);
    ra_5108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1317_inst_ack_0, ack => cp_elements(300)); -- 
    cr_5109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => binary_1317_inst_req_1); -- 
    ca_5110_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1317_inst_ack_1, ack => cp_elements(301)); -- 
    cp_elements(302) <= cp_elements(301);
    cp_elements(303) <= false;
    cp_elements(304) <= cp_elements(303);
    cp_elements(305) <= cp_elements(301);
    branch_req_5118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => if_stmt_1319_branch_req_0); -- 
    cp_elements(306) <= cp_elements(305);
    cp_elements(307) <= cp_elements(306);
    if_choice_transition_5123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1319_branch_ack_1, ack => cp_elements(308)); -- 
    cp_elements(309) <= cp_elements(306);
    else_choice_transition_5127_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1319_branch_ack_0, ack => cp_elements(310)); -- 
    cp_elements(311) <= cp_elements(7);
    cpelement_group_312 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(314));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(312),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(312), ack => binary_1330_inst_req_0); -- 
    cp_elements(313) <= cp_elements(311);
    cp_elements(314) <= cp_elements(311);
    ra_5142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1330_inst_ack_0, ack => cp_elements(315)); -- 
    cr_5143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => binary_1330_inst_req_1); -- 
    ca_5144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1330_inst_ack_1, ack => cp_elements(316)); -- 
    cp_elements(317) <= cp_elements(8);
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(319) & cp_elements(320));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => binary_1353_inst_req_0); -- 
    cp_elements(319) <= cp_elements(317);
    cp_elements(320) <= cp_elements(317);
    ra_5157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1353_inst_ack_0, ack => cp_elements(321)); -- 
    cr_5158_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => binary_1353_inst_req_1); -- 
    ca_5159_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1353_inst_ack_1, ack => cp_elements(322)); -- 
    cpelement_group_323 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(322) & cp_elements(324) & cp_elements(325));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(323),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => binary_1358_inst_req_0); -- 
    cp_elements(324) <= cp_elements(317);
    cp_elements(325) <= cp_elements(317);
    ra_5170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1358_inst_ack_0, ack => cp_elements(326)); -- 
    cr_5171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => binary_1358_inst_req_1); -- 
    ca_5172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1358_inst_ack_1, ack => cp_elements(327)); -- 
    cpelement_group_328 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(329) & cp_elements(330));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(328),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => binary_1364_inst_req_0); -- 
    cp_elements(329) <= cp_elements(317);
    cp_elements(330) <= cp_elements(317);
    ra_5182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1364_inst_ack_0, ack => cp_elements(331)); -- 
    cr_5183_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => binary_1364_inst_req_1); -- 
    ca_5184_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1364_inst_ack_1, ack => cp_elements(332)); -- 
    cpelement_group_333 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(332) & cp_elements(334));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(333),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => binary_1370_inst_req_0); -- 
    cp_elements(334) <= cp_elements(317);
    ra_5194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1370_inst_ack_0, ack => cp_elements(335)); -- 
    cr_5195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => binary_1370_inst_req_1); -- 
    ca_5196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1370_inst_ack_1, ack => cp_elements(336)); -- 
    index_resize_req_5211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => array_obj_ref_1374_index_0_resize_req_0); -- 
    cp_elements(337) <= cp_elements(317);
    cpelement_group_338 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(337) & cp_elements(346));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(338),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => array_obj_ref_1374_final_reg_req_0); -- 
    cp_elements(339) <= cp_elements(317);
    base_resize_req_5227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => array_obj_ref_1374_base_resize_req_0); -- 
    index_resize_ack_5212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_index_0_resize_ack_0, ack => cp_elements(340)); -- 
    scale_rename_req_5216_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => array_obj_ref_1374_index_0_rename_req_0); -- 
    scale_rename_ack_5217_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_index_0_rename_ack_0, ack => cp_elements(341)); -- 
    final_index_req_5221_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => array_obj_ref_1374_offset_inst_req_0); -- 
    final_index_ack_5222_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_offset_inst_ack_0, ack => cp_elements(342)); -- 
    base_resize_ack_5228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_base_resize_ack_0, ack => cp_elements(343)); -- 
    cpelement_group_344 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(342) & cp_elements(343));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_5233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(344), ack => array_obj_ref_1374_root_address_inst_req_0); -- 
    plus_base_ra_5234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_root_address_inst_ack_0, ack => cp_elements(345)); -- 
    plus_base_cr_5235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => array_obj_ref_1374_root_address_inst_req_1); -- 
    plus_base_ca_5236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_root_address_inst_ack_1, ack => cp_elements(346)); -- 
    final_reg_ack_5241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1374_final_reg_ack_0, ack => cp_elements(347)); -- 
    cpelement_group_348 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(348),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => type_cast_1378_inst_req_0); -- 
    cp_elements(349) <= cp_elements(317);
    ack_5251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1378_inst_ack_0, ack => cp_elements(350)); -- 
    base_resize_req_5264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => ptr_deref_1382_base_resize_req_0); -- 
    base_resize_ack_5265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_base_resize_ack_0, ack => cp_elements(351)); -- 
    sum_rename_req_5269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => ptr_deref_1382_root_address_inst_req_0); -- 
    cp_elements(352) <= ptr_deref_1382_root_address_inst_ack_0;
    cp_elements(353) <= cp_elements(352);
    rr_5277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => ptr_deref_1382_addr_0_req_0); -- 
    ra_5278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_addr_0_ack_0, ack => cp_elements(354)); -- 
    cr_5279_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(354), ack => ptr_deref_1382_addr_0_req_1); -- 
    ca_5280_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_addr_0_ack_1, ack => cp_elements(355)); -- 
    cp_elements(356) <= cp_elements(352);
    rr_5284_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => ptr_deref_1382_addr_1_req_0); -- 
    ra_5285_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_addr_1_ack_0, ack => cp_elements(357)); -- 
    cr_5286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => ptr_deref_1382_addr_1_req_1); -- 
    ca_5287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_addr_1_ack_1, ack => cp_elements(358)); -- 
    cpelement_group_359 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(355) & cp_elements(358));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(359),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(360) <= cp_elements(359);
    rr_5297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => ptr_deref_1382_load_0_req_0); -- 
    ra_5298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_0_ack_0, ack => cp_elements(361)); -- 
    cp_elements(362) <= cp_elements(359);
    rr_5302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => ptr_deref_1382_load_1_req_0); -- 
    ra_5303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_1_ack_0, ack => cp_elements(363)); -- 
    cpelement_group_364 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(363));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(364),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(365) <= cp_elements(364);
    cr_5313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(365), ack => ptr_deref_1382_load_0_req_1); -- 
    ca_5314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_0_ack_1, ack => cp_elements(366)); -- 
    cp_elements(367) <= cp_elements(364);
    cr_5318_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(367), ack => ptr_deref_1382_load_1_req_1); -- 
    ca_5319_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_load_1_ack_1, ack => cp_elements(368)); -- 
    cpelement_group_369 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(366) & cp_elements(368));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(369),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_5320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(369), ack => ptr_deref_1382_gather_scatter_req_0); -- 
    merge_ack_5321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1382_gather_scatter_ack_0, ack => cp_elements(370)); -- 
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(370) & cp_elements(372));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => type_cast_1386_inst_req_0); -- 
    cp_elements(372) <= cp_elements(317);
    ack_5331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1386_inst_ack_0, ack => cp_elements(373)); -- 
    cpelement_group_374 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(373) & cp_elements(375) & cp_elements(376));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(374),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(374), ack => binary_1391_inst_req_0); -- 
    cp_elements(375) <= cp_elements(317);
    cp_elements(376) <= cp_elements(317);
    ra_5342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1391_inst_ack_0, ack => cp_elements(377)); -- 
    cr_5343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(377), ack => binary_1391_inst_req_1); -- 
    ca_5344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1391_inst_ack_1, ack => cp_elements(378)); -- 
    cpelement_group_379 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(380) & cp_elements(383));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(379),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5360_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(379), ack => binary_1399_inst_req_0); -- 
    cp_elements(380) <= cp_elements(317);
    cpelement_group_381 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(327) & cp_elements(382));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(381),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => type_cast_1395_inst_req_0); -- 
    cp_elements(382) <= cp_elements(317);
    ack_5356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1395_inst_ack_0, ack => cp_elements(383)); -- 
    ra_5361_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1399_inst_ack_0, ack => cp_elements(384)); -- 
    cr_5362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => binary_1399_inst_req_1); -- 
    ca_5363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1399_inst_ack_1, ack => cp_elements(385)); -- 
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(387) & cp_elements(388));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => binary_1405_inst_req_0); -- 
    cp_elements(387) <= cp_elements(317);
    cp_elements(388) <= cp_elements(317);
    ra_5373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1405_inst_ack_0, ack => cp_elements(389)); -- 
    cr_5374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(389), ack => binary_1405_inst_req_1); -- 
    ca_5375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1405_inst_ack_1, ack => cp_elements(390)); -- 
    cpelement_group_391 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(378) & cp_elements(385) & cp_elements(390));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(391),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(392) <= cp_elements(9);
    cp_elements(393) <= false;
    cp_elements(394) <= cp_elements(393);
    cp_elements(395) <= cp_elements(9);
    branch_req_5383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(395), ack => if_stmt_1407_branch_req_0); -- 
    cp_elements(396) <= cp_elements(395);
    cp_elements(397) <= cp_elements(396);
    if_choice_transition_5388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1407_branch_ack_1, ack => cp_elements(398)); -- 
    cp_elements(399) <= cp_elements(396);
    else_choice_transition_5392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1407_branch_ack_0, ack => cp_elements(400)); -- 
    cp_elements(401) <= cp_elements(10);
    cpelement_group_402 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(403) & cp_elements(404));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(402),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => binary_1418_inst_req_0); -- 
    cp_elements(403) <= cp_elements(401);
    cp_elements(404) <= cp_elements(401);
    ra_5407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1418_inst_ack_0, ack => cp_elements(405)); -- 
    cr_5408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(405), ack => binary_1418_inst_req_1); -- 
    ca_5409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1418_inst_ack_1, ack => cp_elements(406)); -- 
    index_resize_req_5424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => array_obj_ref_1422_index_0_resize_req_0); -- 
    cp_elements(407) <= cp_elements(401);
    cpelement_group_408 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(407) & cp_elements(416));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(408),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5453_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(408), ack => array_obj_ref_1422_final_reg_req_0); -- 
    cp_elements(409) <= cp_elements(401);
    base_resize_req_5440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(409), ack => array_obj_ref_1422_base_resize_req_0); -- 
    index_resize_ack_5425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_index_0_resize_ack_0, ack => cp_elements(410)); -- 
    scale_rename_req_5429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(410), ack => array_obj_ref_1422_index_0_rename_req_0); -- 
    scale_rename_ack_5430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_index_0_rename_ack_0, ack => cp_elements(411)); -- 
    final_index_req_5434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => array_obj_ref_1422_offset_inst_req_0); -- 
    final_index_ack_5435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_offset_inst_ack_0, ack => cp_elements(412)); -- 
    base_resize_ack_5441_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_base_resize_ack_0, ack => cp_elements(413)); -- 
    cpelement_group_414 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(412) & cp_elements(413));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(414),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_5446_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => array_obj_ref_1422_root_address_inst_req_0); -- 
    plus_base_ra_5447_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_root_address_inst_ack_0, ack => cp_elements(415)); -- 
    plus_base_cr_5448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(415), ack => array_obj_ref_1422_root_address_inst_req_1); -- 
    plus_base_ca_5449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_root_address_inst_ack_1, ack => cp_elements(416)); -- 
    final_reg_ack_5454_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1422_final_reg_ack_0, ack => cp_elements(417)); -- 
    cp_elements(418) <= cp_elements(11);
    cpelement_group_419 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(420) & cp_elements(421));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(419),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(419), ack => binary_1450_inst_req_0); -- 
    cp_elements(420) <= cp_elements(418);
    cp_elements(421) <= cp_elements(418);
    ra_5467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1450_inst_ack_0, ack => cp_elements(422)); -- 
    cr_5468_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(422), ack => binary_1450_inst_req_1); -- 
    ca_5469_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1450_inst_ack_1, ack => cp_elements(423)); -- 
    cp_elements(424) <= cp_elements(423);
    cp_elements(425) <= false;
    cp_elements(426) <= cp_elements(425);
    cp_elements(427) <= cp_elements(423);
    branch_req_5477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(427), ack => if_stmt_1452_branch_req_0); -- 
    cp_elements(428) <= cp_elements(427);
    cp_elements(429) <= cp_elements(428);
    if_choice_transition_5482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1452_branch_ack_1, ack => cp_elements(430)); -- 
    cp_elements(431) <= cp_elements(428);
    cp_elements(432) <= if_stmt_1452_branch_ack_0;
    cp_elements(433) <= cp_elements(12);
    cp_elements(434) <= cp_elements(433);
    base_resize_req_5504_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(434), ack => ptr_deref_1461_base_resize_req_0); -- 
    base_resize_ack_5505_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_base_resize_ack_0, ack => cp_elements(435)); -- 
    sum_rename_req_5509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => ptr_deref_1461_root_address_inst_req_0); -- 
    sum_rename_ack_5510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_root_address_inst_ack_0, ack => cp_elements(436)); -- 
    root_rename_req_5514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => ptr_deref_1461_addr_0_req_0); -- 
    root_rename_ack_5515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_addr_0_ack_0, ack => cp_elements(437)); -- 
    rr_5525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(437), ack => ptr_deref_1461_load_0_req_0); -- 
    ra_5526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_load_0_ack_0, ack => cp_elements(438)); -- 
    cr_5536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => ptr_deref_1461_load_0_req_1); -- 
    ca_5537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_load_0_ack_1, ack => cp_elements(439)); -- 
    merge_req_5538_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(439), ack => ptr_deref_1461_gather_scatter_req_0); -- 
    merge_ack_5539_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1461_gather_scatter_ack_0, ack => cp_elements(440)); -- 
    cpelement_group_441 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(440) & cp_elements(442));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(441),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(441), ack => type_cast_1465_inst_req_0); -- 
    cp_elements(442) <= cp_elements(433);
    ack_5549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1465_inst_ack_0, ack => cp_elements(443)); -- 
    cpelement_group_444 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(443) & cp_elements(445) & cp_elements(446));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(444),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(444), ack => binary_1470_inst_req_0); -- 
    cp_elements(445) <= cp_elements(433);
    cp_elements(446) <= cp_elements(433);
    ra_5560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1470_inst_ack_0, ack => cp_elements(447)); -- 
    cr_5561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(447), ack => binary_1470_inst_req_1); -- 
    cp_elements(448) <= binary_1470_inst_ack_1;
    cp_elements(449) <= cp_elements(969);
    cpelement_group_450 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(451) & cp_elements(452));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(450),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(450), ack => binary_1485_inst_req_0); -- 
    cp_elements(451) <= cp_elements(449);
    cp_elements(452) <= cp_elements(449);
    ra_5575_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1485_inst_ack_0, ack => cp_elements(453)); -- 
    cr_5576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(453), ack => binary_1485_inst_req_1); -- 
    ca_5577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1485_inst_ack_1, ack => cp_elements(454)); -- 
    cpelement_group_455 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(456) & cp_elements(457));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(455),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => binary_1491_inst_req_0); -- 
    cp_elements(456) <= cp_elements(449);
    cp_elements(457) <= cp_elements(449);
    ra_5587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1491_inst_ack_0, ack => cp_elements(458)); -- 
    cr_5588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => binary_1491_inst_req_1); -- 
    ca_5589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1491_inst_ack_1, ack => cp_elements(459)); -- 
    cpelement_group_460 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(454) & cp_elements(459) & cp_elements(461));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(460),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => binary_1496_inst_req_0); -- 
    cp_elements(461) <= cp_elements(449);
    ra_5600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1496_inst_ack_0, ack => cp_elements(462)); -- 
    cr_5601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => binary_1496_inst_req_1); -- 
    cp_elements(463) <= binary_1496_inst_ack_1;
    cpelement_group_464 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(465) & cp_elements(466));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(464),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(464), ack => binary_1502_inst_req_0); -- 
    cp_elements(465) <= cp_elements(449);
    cp_elements(466) <= cp_elements(463);
    ra_5612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1502_inst_ack_0, ack => cp_elements(467)); -- 
    cr_5613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => binary_1502_inst_req_1); -- 
    ca_5614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1502_inst_ack_1, ack => cp_elements(468)); -- 
    cpelement_group_469 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(470) & cp_elements(471));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(469),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => binary_1507_inst_req_0); -- 
    cp_elements(470) <= cp_elements(449);
    cp_elements(471) <= cp_elements(463);
    ra_5625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_0, ack => cp_elements(472)); -- 
    cr_5626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(472), ack => binary_1507_inst_req_1); -- 
    ca_5627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1507_inst_ack_1, ack => cp_elements(473)); -- 
    cpelement_group_474 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(473) & cp_elements(475));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(474),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_5636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(474), ack => type_cast_1511_inst_req_0); -- 
    cp_elements(475) <= cp_elements(449);
    ack_5637_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1511_inst_ack_0, ack => cp_elements(476)); -- 
    cpelement_group_477 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(476) & cp_elements(478));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(477),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => binary_1517_inst_req_0); -- 
    cp_elements(478) <= cp_elements(449);
    ra_5647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1517_inst_ack_0, ack => cp_elements(479)); -- 
    cr_5648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(479), ack => binary_1517_inst_req_1); -- 
    ca_5649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1517_inst_ack_1, ack => cp_elements(480)); -- 
    cp_elements(481) <= cp_elements(480);
    cp_elements(482) <= false;
    cp_elements(483) <= cp_elements(482);
    cp_elements(484) <= cp_elements(480);
    branch_req_5657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => if_stmt_1519_branch_req_0); -- 
    cp_elements(485) <= cp_elements(484);
    cp_elements(486) <= cp_elements(485);
    if_choice_transition_5662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1519_branch_ack_1, ack => cp_elements(487)); -- 
    cp_elements(488) <= cp_elements(485);
    else_choice_transition_5666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1519_branch_ack_0, ack => cp_elements(489)); -- 
    cpelement_group_490 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(491) & cp_elements(492));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(490),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => binary_1530_inst_req_0); -- 
    cp_elements(491) <= cp_elements(13);
    cp_elements(492) <= cp_elements(13);
    ra_5684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1530_inst_ack_0, ack => cp_elements(493)); -- 
    cr_5685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(493), ack => binary_1530_inst_req_1); -- 
    ca_5686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1530_inst_ack_1, ack => cp_elements(494)); -- 
    pipe_wreq_5691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(494), ack => simple_obj_ref_1527_inst_req_0); -- 
    pipe_wack_5692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1527_inst_ack_0, ack => cp_elements(495)); -- 
    cp_elements(496) <= cp_elements(487);
    cp_elements(497) <= cp_elements(496);
    cpelement_group_498 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(497) & cp_elements(502));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(498),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(498), ack => array_obj_ref_1540_final_reg_req_0); -- 
    cp_elements(499) <= cp_elements(496);
    base_resize_req_5706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => array_obj_ref_1540_base_resize_req_0); -- 
    base_resize_ack_5707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1540_base_resize_ack_0, ack => cp_elements(500)); -- 
    plus_base_rr_5712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => array_obj_ref_1540_root_address_inst_req_0); -- 
    plus_base_ra_5713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1540_root_address_inst_ack_0, ack => cp_elements(501)); -- 
    plus_base_cr_5714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => array_obj_ref_1540_root_address_inst_req_1); -- 
    plus_base_ca_5715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1540_root_address_inst_ack_1, ack => cp_elements(502)); -- 
    final_reg_ack_5720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1540_final_reg_ack_0, ack => cp_elements(503)); -- 
    base_resize_req_5734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => ptr_deref_1543_base_resize_req_0); -- 
    cp_elements(504) <= cp_elements(496);
    cpelement_group_505 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(504) & cp_elements(520));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(505),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5775_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => ptr_deref_1543_gather_scatter_req_0); -- 
    base_resize_ack_5735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_base_resize_ack_0, ack => cp_elements(506)); -- 
    sum_rename_req_5739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_1543_root_address_inst_req_0); -- 
    cp_elements(507) <= ptr_deref_1543_root_address_inst_ack_0;
    cp_elements(508) <= cp_elements(507);
    rr_5747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(508), ack => ptr_deref_1543_addr_0_req_0); -- 
    ra_5748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_0_ack_0, ack => cp_elements(509)); -- 
    cr_5749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(509), ack => ptr_deref_1543_addr_0_req_1); -- 
    ca_5750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_0_ack_1, ack => cp_elements(510)); -- 
    cp_elements(511) <= cp_elements(507);
    rr_5754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(511), ack => ptr_deref_1543_addr_1_req_0); -- 
    ra_5755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_1_ack_0, ack => cp_elements(512)); -- 
    cr_5756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(512), ack => ptr_deref_1543_addr_1_req_1); -- 
    ca_5757_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_1_ack_1, ack => cp_elements(513)); -- 
    cp_elements(514) <= cp_elements(507);
    rr_5761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => ptr_deref_1543_addr_2_req_0); -- 
    ra_5762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_2_ack_0, ack => cp_elements(515)); -- 
    cr_5763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => ptr_deref_1543_addr_2_req_1); -- 
    ca_5764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_2_ack_1, ack => cp_elements(516)); -- 
    cp_elements(517) <= cp_elements(507);
    rr_5768_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => ptr_deref_1543_addr_3_req_0); -- 
    ra_5769_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_3_ack_0, ack => cp_elements(518)); -- 
    cr_5770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(518), ack => ptr_deref_1543_addr_3_req_1); -- 
    ca_5771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_addr_3_ack_1, ack => cp_elements(519)); -- 
    cpelement_group_520 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(510) & cp_elements(513) & cp_elements(516) & cp_elements(519));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(520),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(521) <= ptr_deref_1543_gather_scatter_ack_0;
    cp_elements(522) <= cp_elements(521);
    rr_5783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(522), ack => ptr_deref_1543_store_0_req_0); -- 
    ra_5784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_0_ack_0, ack => cp_elements(523)); -- 
    cp_elements(524) <= cp_elements(521);
    rr_5788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => ptr_deref_1543_store_1_req_0); -- 
    ra_5789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_1_ack_0, ack => cp_elements(525)); -- 
    cp_elements(526) <= cp_elements(521);
    rr_5793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(526), ack => ptr_deref_1543_store_2_req_0); -- 
    ra_5794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_2_ack_0, ack => cp_elements(527)); -- 
    cp_elements(528) <= cp_elements(521);
    rr_5798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => ptr_deref_1543_store_3_req_0); -- 
    ra_5799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_3_ack_0, ack => cp_elements(529)); -- 
    cpelement_group_530 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(523) & cp_elements(525) & cp_elements(527) & cp_elements(529));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(530),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(531) <= cp_elements(530);
    cp_elements(532) <= cp_elements(531);
    cr_5809_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(532), ack => ptr_deref_1543_store_0_req_1); -- 
    ca_5810_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_0_ack_1, ack => cp_elements(533)); -- 
    cp_elements(534) <= cp_elements(531);
    cr_5814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => ptr_deref_1543_store_1_req_1); -- 
    ca_5815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_1_ack_1, ack => cp_elements(535)); -- 
    cp_elements(536) <= cp_elements(531);
    cr_5819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(536), ack => ptr_deref_1543_store_2_req_1); -- 
    ca_5820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_2_ack_1, ack => cp_elements(537)); -- 
    cp_elements(538) <= cp_elements(531);
    cr_5824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(538), ack => ptr_deref_1543_store_3_req_1); -- 
    ca_5825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1543_store_3_ack_1, ack => cp_elements(539)); -- 
    cpelement_group_540 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(533) & cp_elements(535) & cp_elements(537) & cp_elements(539));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(540),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_541 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(542) & cp_elements(543));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(541),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_5834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => binary_1550_inst_req_0); -- 
    cp_elements(542) <= cp_elements(496);
    cp_elements(543) <= cp_elements(496);
    ra_5835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1550_inst_ack_0, ack => cp_elements(544)); -- 
    cr_5836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(544), ack => binary_1550_inst_req_1); -- 
    ca_5837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1550_inst_ack_1, ack => cp_elements(545)); -- 
    index_resize_req_5852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(545), ack => array_obj_ref_1554_index_0_resize_req_0); -- 
    cp_elements(546) <= cp_elements(496);
    cpelement_group_547 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(546) & cp_elements(555));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(547),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(547), ack => array_obj_ref_1554_final_reg_req_0); -- 
    cp_elements(548) <= cp_elements(496);
    base_resize_req_5868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => array_obj_ref_1554_base_resize_req_0); -- 
    index_resize_ack_5853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_index_0_resize_ack_0, ack => cp_elements(549)); -- 
    scale_rename_req_5857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(549), ack => array_obj_ref_1554_index_0_rename_req_0); -- 
    scale_rename_ack_5858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_index_0_rename_ack_0, ack => cp_elements(550)); -- 
    final_index_req_5862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => array_obj_ref_1554_offset_inst_req_0); -- 
    final_index_ack_5863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_offset_inst_ack_0, ack => cp_elements(551)); -- 
    base_resize_ack_5869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_base_resize_ack_0, ack => cp_elements(552)); -- 
    cpelement_group_553 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(551) & cp_elements(552));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(553),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_5874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(553), ack => array_obj_ref_1554_root_address_inst_req_0); -- 
    plus_base_ra_5875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_root_address_inst_ack_0, ack => cp_elements(554)); -- 
    plus_base_cr_5876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => array_obj_ref_1554_root_address_inst_req_1); -- 
    plus_base_ca_5877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_root_address_inst_ack_1, ack => cp_elements(555)); -- 
    final_reg_ack_5882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1554_final_reg_ack_0, ack => cp_elements(556)); -- 
    cp_elements(557) <= cp_elements(496);
    cpelement_group_558 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(557) & cp_elements(562));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(558),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_5906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(558), ack => array_obj_ref_1561_final_reg_req_0); -- 
    cp_elements(559) <= cp_elements(496);
    base_resize_req_5893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(559), ack => array_obj_ref_1561_base_resize_req_0); -- 
    base_resize_ack_5894_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1561_base_resize_ack_0, ack => cp_elements(560)); -- 
    plus_base_rr_5899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(560), ack => array_obj_ref_1561_root_address_inst_req_0); -- 
    plus_base_ra_5900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1561_root_address_inst_ack_0, ack => cp_elements(561)); -- 
    plus_base_cr_5901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(561), ack => array_obj_ref_1561_root_address_inst_req_1); -- 
    plus_base_ca_5902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1561_root_address_inst_ack_1, ack => cp_elements(562)); -- 
    cp_elements(563) <= array_obj_ref_1561_final_reg_ack_0;
    cpelement_group_564 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(530) & cp_elements(556) & cp_elements(563) & cp_elements(580));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(564),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_5962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => ptr_deref_1564_gather_scatter_req_0); -- 
    cp_elements(565) <= cp_elements(563);
    base_resize_req_5921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(565), ack => ptr_deref_1564_base_resize_req_0); -- 
    base_resize_ack_5922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_base_resize_ack_0, ack => cp_elements(566)); -- 
    sum_rename_req_5926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => ptr_deref_1564_root_address_inst_req_0); -- 
    cp_elements(567) <= ptr_deref_1564_root_address_inst_ack_0;
    cp_elements(568) <= cp_elements(567);
    rr_5934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_1564_addr_0_req_0); -- 
    ra_5935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_0_ack_0, ack => cp_elements(569)); -- 
    cr_5936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(569), ack => ptr_deref_1564_addr_0_req_1); -- 
    ca_5937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_0_ack_1, ack => cp_elements(570)); -- 
    cp_elements(571) <= cp_elements(567);
    rr_5941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => ptr_deref_1564_addr_1_req_0); -- 
    ra_5942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_1_ack_0, ack => cp_elements(572)); -- 
    cr_5943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(572), ack => ptr_deref_1564_addr_1_req_1); -- 
    ca_5944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_1_ack_1, ack => cp_elements(573)); -- 
    cp_elements(574) <= cp_elements(567);
    rr_5948_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => ptr_deref_1564_addr_2_req_0); -- 
    ra_5949_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_2_ack_0, ack => cp_elements(575)); -- 
    cr_5950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => ptr_deref_1564_addr_2_req_1); -- 
    ca_5951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_2_ack_1, ack => cp_elements(576)); -- 
    cp_elements(577) <= cp_elements(567);
    rr_5955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => ptr_deref_1564_addr_3_req_0); -- 
    ra_5956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_3_ack_0, ack => cp_elements(578)); -- 
    cr_5957_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => ptr_deref_1564_addr_3_req_1); -- 
    ca_5958_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_addr_3_ack_1, ack => cp_elements(579)); -- 
    cpelement_group_580 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(570) & cp_elements(573) & cp_elements(576) & cp_elements(579));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(580),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(581) <= ptr_deref_1564_gather_scatter_ack_0;
    cp_elements(582) <= cp_elements(581);
    rr_5970_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(582), ack => ptr_deref_1564_store_0_req_0); -- 
    ra_5971_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_0_ack_0, ack => cp_elements(583)); -- 
    cp_elements(584) <= cp_elements(581);
    rr_5975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => ptr_deref_1564_store_1_req_0); -- 
    ra_5976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_1_ack_0, ack => cp_elements(585)); -- 
    cp_elements(586) <= cp_elements(581);
    rr_5980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(586), ack => ptr_deref_1564_store_2_req_0); -- 
    ra_5981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_2_ack_0, ack => cp_elements(587)); -- 
    cp_elements(588) <= cp_elements(581);
    rr_5985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(588), ack => ptr_deref_1564_store_3_req_0); -- 
    ra_5986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_3_ack_0, ack => cp_elements(589)); -- 
    cpelement_group_590 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(583) & cp_elements(585) & cp_elements(587) & cp_elements(589));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(590),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(591) <= cp_elements(590);
    cr_5996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => ptr_deref_1564_store_0_req_1); -- 
    ca_5997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_0_ack_1, ack => cp_elements(592)); -- 
    cp_elements(593) <= cp_elements(590);
    cr_6001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_1564_store_1_req_1); -- 
    ca_6002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_1_ack_1, ack => cp_elements(594)); -- 
    cp_elements(595) <= cp_elements(590);
    cr_6006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => ptr_deref_1564_store_2_req_1); -- 
    ca_6007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_2_ack_1, ack => cp_elements(596)); -- 
    cp_elements(597) <= cp_elements(590);
    cr_6011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(597), ack => ptr_deref_1564_store_3_req_1); -- 
    ca_6012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1564_store_3_ack_1, ack => cp_elements(598)); -- 
    cpelement_group_599 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(592) & cp_elements(594) & cp_elements(596) & cp_elements(598));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(599),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_600 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(601) & cp_elements(602) & cp_elements(603));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(600),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => binary_1570_inst_req_0); -- 
    cp_elements(601) <= cp_elements(496);
    cp_elements(602) <= cp_elements(496);
    cp_elements(603) <= cp_elements(496);
    ra_6023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1570_inst_ack_0, ack => cp_elements(604)); -- 
    cr_6024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => binary_1570_inst_req_1); -- 
    ca_6025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1570_inst_ack_1, ack => cp_elements(605)); -- 
    cpelement_group_606 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(540) & cp_elements(599) & cp_elements(605));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(606),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(607) <= cp_elements(14);
    cp_elements(608) <= false;
    cp_elements(609) <= cp_elements(608);
    cp_elements(610) <= cp_elements(14);
    branch_req_6033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(610), ack => if_stmt_1572_branch_req_0); -- 
    cp_elements(611) <= cp_elements(610);
    cp_elements(612) <= cp_elements(611);
    if_choice_transition_6038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1572_branch_ack_1, ack => cp_elements(613)); -- 
    cp_elements(614) <= cp_elements(611);
    else_choice_transition_6042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1572_branch_ack_0, ack => cp_elements(615)); -- 
    cp_elements(616) <= cp_elements(15);
    cpelement_group_617 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(618) & cp_elements(619) & cp_elements(620));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(617),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(617), ack => binary_1582_inst_req_0); -- 
    cp_elements(618) <= cp_elements(616);
    cp_elements(619) <= cp_elements(616);
    cp_elements(620) <= cp_elements(616);
    ra_6058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1582_inst_ack_0, ack => cp_elements(621)); -- 
    cr_6059_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(621), ack => binary_1582_inst_req_1); -- 
    cp_elements(622) <= binary_1582_inst_ack_1;
    cpelement_group_623 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(624) & cp_elements(625) & cp_elements(626));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(623),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(623), ack => binary_1587_inst_req_0); -- 
    cp_elements(624) <= cp_elements(616);
    cp_elements(625) <= cp_elements(616);
    cp_elements(626) <= cp_elements(622);
    ra_6071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1587_inst_ack_0, ack => cp_elements(627)); -- 
    cr_6072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => binary_1587_inst_req_1); -- 
    ca_6073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1587_inst_ack_1, ack => cp_elements(628)); -- 
    cp_elements(629) <= cp_elements(616);
    cpelement_group_630 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(628) & cp_elements(629) & cp_elements(631) & cp_elements(632));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(630),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(630), ack => ternary_1593_inst_req_0); -- 
    cp_elements(631) <= cp_elements(616);
    cp_elements(632) <= cp_elements(622);
    ack_6085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ternary_1593_inst_ack_0, ack => cp_elements(633)); -- 
    cpelement_group_634 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(633) & cp_elements(635));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(634),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(634), ack => binary_1599_inst_req_0); -- 
    cp_elements(635) <= cp_elements(616);
    ra_6095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1599_inst_ack_0, ack => cp_elements(636)); -- 
    cr_6096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => binary_1599_inst_req_1); -- 
    ca_6097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1599_inst_ack_1, ack => cp_elements(637)); -- 
    index_resize_req_6112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(637), ack => array_obj_ref_1603_index_0_resize_req_0); -- 
    cp_elements(638) <= cp_elements(616);
    cpelement_group_639 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(638) & cp_elements(647));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(639),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => array_obj_ref_1603_final_reg_req_0); -- 
    cp_elements(640) <= cp_elements(616);
    base_resize_req_6128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => array_obj_ref_1603_base_resize_req_0); -- 
    index_resize_ack_6113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_index_0_resize_ack_0, ack => cp_elements(641)); -- 
    scale_rename_req_6117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(641), ack => array_obj_ref_1603_index_0_rename_req_0); -- 
    scale_rename_ack_6118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_index_0_rename_ack_0, ack => cp_elements(642)); -- 
    final_index_req_6122_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => array_obj_ref_1603_offset_inst_req_0); -- 
    final_index_ack_6123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_offset_inst_ack_0, ack => cp_elements(643)); -- 
    base_resize_ack_6129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_base_resize_ack_0, ack => cp_elements(644)); -- 
    cpelement_group_645 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(643) & cp_elements(644));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(645),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_6134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(645), ack => array_obj_ref_1603_root_address_inst_req_0); -- 
    plus_base_ra_6135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_root_address_inst_ack_0, ack => cp_elements(646)); -- 
    plus_base_cr_6136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(646), ack => array_obj_ref_1603_root_address_inst_req_1); -- 
    plus_base_ca_6137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_root_address_inst_ack_1, ack => cp_elements(647)); -- 
    final_reg_ack_6142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1603_final_reg_ack_0, ack => cp_elements(648)); -- 
    cpelement_group_649 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(648) & cp_elements(650) & cp_elements(666));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(649),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(649), ack => ptr_deref_1606_gather_scatter_req_0); -- 
    cp_elements(650) <= cp_elements(616);
    cp_elements(651) <= cp_elements(650);
    base_resize_req_6156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(651), ack => ptr_deref_1606_base_resize_req_0); -- 
    base_resize_ack_6157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_base_resize_ack_0, ack => cp_elements(652)); -- 
    sum_rename_req_6161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_1606_root_address_inst_req_0); -- 
    cp_elements(653) <= ptr_deref_1606_root_address_inst_ack_0;
    cp_elements(654) <= cp_elements(653);
    rr_6169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_1606_addr_0_req_0); -- 
    ra_6170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_0_ack_0, ack => cp_elements(655)); -- 
    cr_6171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(655), ack => ptr_deref_1606_addr_0_req_1); -- 
    ca_6172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_0_ack_1, ack => cp_elements(656)); -- 
    cp_elements(657) <= cp_elements(653);
    rr_6176_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(657), ack => ptr_deref_1606_addr_1_req_0); -- 
    ra_6177_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_1_ack_0, ack => cp_elements(658)); -- 
    cr_6178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => ptr_deref_1606_addr_1_req_1); -- 
    ca_6179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_1_ack_1, ack => cp_elements(659)); -- 
    cp_elements(660) <= cp_elements(653);
    rr_6183_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => ptr_deref_1606_addr_2_req_0); -- 
    ra_6184_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_2_ack_0, ack => cp_elements(661)); -- 
    cr_6185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(661), ack => ptr_deref_1606_addr_2_req_1); -- 
    ca_6186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_2_ack_1, ack => cp_elements(662)); -- 
    cp_elements(663) <= cp_elements(653);
    rr_6190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => ptr_deref_1606_addr_3_req_0); -- 
    ra_6191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_3_ack_0, ack => cp_elements(664)); -- 
    cr_6192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(664), ack => ptr_deref_1606_addr_3_req_1); -- 
    ca_6193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_addr_3_ack_1, ack => cp_elements(665)); -- 
    cpelement_group_666 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(656) & cp_elements(659) & cp_elements(662) & cp_elements(665));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(666),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(667) <= ptr_deref_1606_gather_scatter_ack_0;
    cp_elements(668) <= cp_elements(667);
    rr_6205_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => ptr_deref_1606_store_0_req_0); -- 
    ra_6206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_0_ack_0, ack => cp_elements(669)); -- 
    cp_elements(670) <= cp_elements(667);
    rr_6210_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(670), ack => ptr_deref_1606_store_1_req_0); -- 
    ra_6211_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_1_ack_0, ack => cp_elements(671)); -- 
    cp_elements(672) <= cp_elements(667);
    rr_6215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(672), ack => ptr_deref_1606_store_2_req_0); -- 
    ra_6216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_2_ack_0, ack => cp_elements(673)); -- 
    cp_elements(674) <= cp_elements(667);
    rr_6220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(674), ack => ptr_deref_1606_store_3_req_0); -- 
    ra_6221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_3_ack_0, ack => cp_elements(675)); -- 
    cpelement_group_676 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(669) & cp_elements(671) & cp_elements(673) & cp_elements(675));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(676),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(677) <= cp_elements(676);
    cp_elements(678) <= cp_elements(677);
    cr_6231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => ptr_deref_1606_store_0_req_1); -- 
    ca_6232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_0_ack_1, ack => cp_elements(679)); -- 
    cp_elements(680) <= cp_elements(677);
    cr_6236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => ptr_deref_1606_store_1_req_1); -- 
    ca_6237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_1_ack_1, ack => cp_elements(681)); -- 
    cp_elements(682) <= cp_elements(677);
    cr_6241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => ptr_deref_1606_store_2_req_1); -- 
    ca_6242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_2_ack_1, ack => cp_elements(683)); -- 
    cp_elements(684) <= cp_elements(677);
    cr_6246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_1606_store_3_req_1); -- 
    ca_6247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1606_store_3_ack_1, ack => cp_elements(685)); -- 
    cpelement_group_686 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(679) & cp_elements(681) & cp_elements(683) & cp_elements(685));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(686),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(687) <= cp_elements(616);
    cpelement_group_688 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(687) & cp_elements(692));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(688), ack => array_obj_ref_1612_final_reg_req_0); -- 
    cp_elements(689) <= cp_elements(616);
    base_resize_req_6258_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(689), ack => array_obj_ref_1612_base_resize_req_0); -- 
    base_resize_ack_6259_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_base_resize_ack_0, ack => cp_elements(690)); -- 
    plus_base_rr_6264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => array_obj_ref_1612_root_address_inst_req_0); -- 
    plus_base_ra_6265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_root_address_inst_ack_0, ack => cp_elements(691)); -- 
    plus_base_cr_6266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(691), ack => array_obj_ref_1612_root_address_inst_req_1); -- 
    plus_base_ca_6267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_root_address_inst_ack_1, ack => cp_elements(692)); -- 
    final_reg_ack_6272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1612_final_reg_ack_0, ack => cp_elements(693)); -- 
    cpelement_group_694 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(693) & cp_elements(695));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(694),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => type_cast_1616_inst_req_0); -- 
    cp_elements(695) <= cp_elements(616);
    cp_elements(696) <= type_cast_1616_inst_ack_0;
    cpelement_group_697 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(676) & cp_elements(696) & cp_elements(713));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(697),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(698) <= cp_elements(696);
    base_resize_req_6295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(698), ack => ptr_deref_1620_base_resize_req_0); -- 
    base_resize_ack_6296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_base_resize_ack_0, ack => cp_elements(699)); -- 
    sum_rename_req_6300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_1620_root_address_inst_req_0); -- 
    cp_elements(700) <= ptr_deref_1620_root_address_inst_ack_0;
    cp_elements(701) <= cp_elements(700);
    rr_6308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_1620_addr_0_req_0); -- 
    ra_6309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_0_ack_0, ack => cp_elements(702)); -- 
    cr_6310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => ptr_deref_1620_addr_0_req_1); -- 
    ca_6311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_0_ack_1, ack => cp_elements(703)); -- 
    cp_elements(704) <= cp_elements(700);
    rr_6315_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(704), ack => ptr_deref_1620_addr_1_req_0); -- 
    ra_6316_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_1_ack_0, ack => cp_elements(705)); -- 
    cr_6317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(705), ack => ptr_deref_1620_addr_1_req_1); -- 
    ca_6318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_1_ack_1, ack => cp_elements(706)); -- 
    cp_elements(707) <= cp_elements(700);
    rr_6322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(707), ack => ptr_deref_1620_addr_2_req_0); -- 
    ra_6323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_2_ack_0, ack => cp_elements(708)); -- 
    cr_6324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => ptr_deref_1620_addr_2_req_1); -- 
    ca_6325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_2_ack_1, ack => cp_elements(709)); -- 
    cp_elements(710) <= cp_elements(700);
    rr_6329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => ptr_deref_1620_addr_3_req_0); -- 
    ra_6330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_3_ack_0, ack => cp_elements(711)); -- 
    cr_6331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => ptr_deref_1620_addr_3_req_1); -- 
    ca_6332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_addr_3_ack_1, ack => cp_elements(712)); -- 
    cpelement_group_713 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(703) & cp_elements(706) & cp_elements(709) & cp_elements(712));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(713),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(714) <= cp_elements(697);
    rr_6342_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(714), ack => ptr_deref_1620_load_0_req_0); -- 
    ra_6343_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_0_ack_0, ack => cp_elements(715)); -- 
    cp_elements(716) <= cp_elements(697);
    rr_6347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(716), ack => ptr_deref_1620_load_1_req_0); -- 
    ra_6348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_1_ack_0, ack => cp_elements(717)); -- 
    cp_elements(718) <= cp_elements(697);
    rr_6352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(718), ack => ptr_deref_1620_load_2_req_0); -- 
    ra_6353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_2_ack_0, ack => cp_elements(719)); -- 
    cp_elements(720) <= cp_elements(697);
    rr_6357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => ptr_deref_1620_load_3_req_0); -- 
    ra_6358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_3_ack_0, ack => cp_elements(721)); -- 
    cpelement_group_722 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(715) & cp_elements(717) & cp_elements(719) & cp_elements(721));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(722),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(723) <= cp_elements(722);
    cr_6368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(723), ack => ptr_deref_1620_load_0_req_1); -- 
    ca_6369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_0_ack_1, ack => cp_elements(724)); -- 
    cp_elements(725) <= cp_elements(722);
    cr_6373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => ptr_deref_1620_load_1_req_1); -- 
    ca_6374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_1_ack_1, ack => cp_elements(726)); -- 
    cp_elements(727) <= cp_elements(722);
    cr_6378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => ptr_deref_1620_load_2_req_1); -- 
    ca_6379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_2_ack_1, ack => cp_elements(728)); -- 
    cp_elements(729) <= cp_elements(722);
    cr_6383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => ptr_deref_1620_load_3_req_1); -- 
    ca_6384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_load_3_ack_1, ack => cp_elements(730)); -- 
    cpelement_group_731 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(724) & cp_elements(726) & cp_elements(728) & cp_elements(730));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(731),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(731), ack => ptr_deref_1620_gather_scatter_req_0); -- 
    merge_ack_6386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1620_gather_scatter_ack_0, ack => cp_elements(732)); -- 
    cp_elements(733) <= cp_elements(616);
    cpelement_group_734 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(733) & cp_elements(738));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(734),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(734), ack => array_obj_ref_1627_final_reg_req_0); -- 
    cp_elements(735) <= cp_elements(616);
    base_resize_req_6397_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => array_obj_ref_1627_base_resize_req_0); -- 
    base_resize_ack_6398_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1627_base_resize_ack_0, ack => cp_elements(736)); -- 
    plus_base_rr_6403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => array_obj_ref_1627_root_address_inst_req_0); -- 
    plus_base_ra_6404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1627_root_address_inst_ack_0, ack => cp_elements(737)); -- 
    plus_base_cr_6405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => array_obj_ref_1627_root_address_inst_req_1); -- 
    plus_base_ca_6406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1627_root_address_inst_ack_1, ack => cp_elements(738)); -- 
    final_reg_ack_6411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1627_final_reg_ack_0, ack => cp_elements(739)); -- 
    cpelement_group_740 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(739) & cp_elements(741));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(740),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => type_cast_1631_inst_req_0); -- 
    cp_elements(741) <= cp_elements(616);
    cp_elements(742) <= type_cast_1631_inst_ack_0;
    cpelement_group_743 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(732) & cp_elements(742) & cp_elements(759));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(743),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(743), ack => ptr_deref_1634_gather_scatter_req_0); -- 
    cp_elements(744) <= cp_elements(742);
    base_resize_req_6435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => ptr_deref_1634_base_resize_req_0); -- 
    base_resize_ack_6436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_base_resize_ack_0, ack => cp_elements(745)); -- 
    sum_rename_req_6440_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => ptr_deref_1634_root_address_inst_req_0); -- 
    cp_elements(746) <= ptr_deref_1634_root_address_inst_ack_0;
    cp_elements(747) <= cp_elements(746);
    rr_6448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(747), ack => ptr_deref_1634_addr_0_req_0); -- 
    ra_6449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_0_ack_0, ack => cp_elements(748)); -- 
    cr_6450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(748), ack => ptr_deref_1634_addr_0_req_1); -- 
    ca_6451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_0_ack_1, ack => cp_elements(749)); -- 
    cp_elements(750) <= cp_elements(746);
    rr_6455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(750), ack => ptr_deref_1634_addr_1_req_0); -- 
    ra_6456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_1_ack_0, ack => cp_elements(751)); -- 
    cr_6457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(751), ack => ptr_deref_1634_addr_1_req_1); -- 
    ca_6458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_1_ack_1, ack => cp_elements(752)); -- 
    cp_elements(753) <= cp_elements(746);
    rr_6462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(753), ack => ptr_deref_1634_addr_2_req_0); -- 
    ra_6463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_2_ack_0, ack => cp_elements(754)); -- 
    cr_6464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(754), ack => ptr_deref_1634_addr_2_req_1); -- 
    ca_6465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_2_ack_1, ack => cp_elements(755)); -- 
    cp_elements(756) <= cp_elements(746);
    rr_6469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => ptr_deref_1634_addr_3_req_0); -- 
    ra_6470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_3_ack_0, ack => cp_elements(757)); -- 
    cr_6471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(757), ack => ptr_deref_1634_addr_3_req_1); -- 
    ca_6472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_addr_3_ack_1, ack => cp_elements(758)); -- 
    cpelement_group_759 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(749) & cp_elements(752) & cp_elements(755) & cp_elements(758));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(759),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(760) <= ptr_deref_1634_gather_scatter_ack_0;
    cp_elements(761) <= cp_elements(760);
    rr_6484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => ptr_deref_1634_store_0_req_0); -- 
    ra_6485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_0_ack_0, ack => cp_elements(762)); -- 
    cp_elements(763) <= cp_elements(760);
    rr_6489_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => ptr_deref_1634_store_1_req_0); -- 
    ra_6490_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_1_ack_0, ack => cp_elements(764)); -- 
    cp_elements(765) <= cp_elements(760);
    rr_6494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => ptr_deref_1634_store_2_req_0); -- 
    ra_6495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_2_ack_0, ack => cp_elements(766)); -- 
    cp_elements(767) <= cp_elements(760);
    rr_6499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => ptr_deref_1634_store_3_req_0); -- 
    ra_6500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_3_ack_0, ack => cp_elements(768)); -- 
    cpelement_group_769 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(762) & cp_elements(764) & cp_elements(766) & cp_elements(768));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(769),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(770) <= cp_elements(769);
    cr_6510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => ptr_deref_1634_store_0_req_1); -- 
    ca_6511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_0_ack_1, ack => cp_elements(771)); -- 
    cp_elements(772) <= cp_elements(769);
    cr_6515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => ptr_deref_1634_store_1_req_1); -- 
    ca_6516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_1_ack_1, ack => cp_elements(773)); -- 
    cp_elements(774) <= cp_elements(769);
    cr_6520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => ptr_deref_1634_store_2_req_1); -- 
    ca_6521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_2_ack_1, ack => cp_elements(775)); -- 
    cp_elements(776) <= cp_elements(769);
    cr_6525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => ptr_deref_1634_store_3_req_1); -- 
    ca_6526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1634_store_3_ack_1, ack => cp_elements(777)); -- 
    cpelement_group_778 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(771) & cp_elements(773) & cp_elements(775) & cp_elements(777));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(778),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_779 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(686) & cp_elements(778));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(779),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(780) <= cp_elements(615);
    cp_elements(781) <= cp_elements(780);
    cpelement_group_782 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(781) & cp_elements(786));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(782),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(782), ack => array_obj_ref_1642_final_reg_req_0); -- 
    cp_elements(783) <= cp_elements(780);
    base_resize_req_6540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => array_obj_ref_1642_base_resize_req_0); -- 
    base_resize_ack_6541_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1642_base_resize_ack_0, ack => cp_elements(784)); -- 
    plus_base_rr_6546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(784), ack => array_obj_ref_1642_root_address_inst_req_0); -- 
    plus_base_ra_6547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1642_root_address_inst_ack_0, ack => cp_elements(785)); -- 
    plus_base_cr_6548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => array_obj_ref_1642_root_address_inst_req_1); -- 
    plus_base_ca_6549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1642_root_address_inst_ack_1, ack => cp_elements(786)); -- 
    final_reg_ack_6554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1642_final_reg_ack_0, ack => cp_elements(787)); -- 
    cpelement_group_788 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(787) & cp_elements(789));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(788),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => type_cast_1646_inst_req_0); -- 
    cp_elements(789) <= cp_elements(780);
    ack_6564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1646_inst_ack_0, ack => cp_elements(790)); -- 
    base_resize_req_6577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => ptr_deref_1650_base_resize_req_0); -- 
    base_resize_ack_6578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_base_resize_ack_0, ack => cp_elements(791)); -- 
    sum_rename_req_6582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(791), ack => ptr_deref_1650_root_address_inst_req_0); -- 
    cp_elements(792) <= ptr_deref_1650_root_address_inst_ack_0;
    cp_elements(793) <= cp_elements(792);
    rr_6590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => ptr_deref_1650_addr_0_req_0); -- 
    ra_6591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_0_ack_0, ack => cp_elements(794)); -- 
    cr_6592_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => ptr_deref_1650_addr_0_req_1); -- 
    ca_6593_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_0_ack_1, ack => cp_elements(795)); -- 
    cp_elements(796) <= cp_elements(792);
    rr_6597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(796), ack => ptr_deref_1650_addr_1_req_0); -- 
    ra_6598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_1_ack_0, ack => cp_elements(797)); -- 
    cr_6599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => ptr_deref_1650_addr_1_req_1); -- 
    ca_6600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_1_ack_1, ack => cp_elements(798)); -- 
    cp_elements(799) <= cp_elements(792);
    rr_6604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => ptr_deref_1650_addr_2_req_0); -- 
    ra_6605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_2_ack_0, ack => cp_elements(800)); -- 
    cr_6606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => ptr_deref_1650_addr_2_req_1); -- 
    ca_6607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_2_ack_1, ack => cp_elements(801)); -- 
    cp_elements(802) <= cp_elements(792);
    rr_6611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(802), ack => ptr_deref_1650_addr_3_req_0); -- 
    ra_6612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_3_ack_0, ack => cp_elements(803)); -- 
    cr_6613_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => ptr_deref_1650_addr_3_req_1); -- 
    ca_6614_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_addr_3_ack_1, ack => cp_elements(804)); -- 
    cpelement_group_805 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(795) & cp_elements(798) & cp_elements(801) & cp_elements(804));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(805),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(806) <= cp_elements(805);
    rr_6624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_1650_load_0_req_0); -- 
    ra_6625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_0_ack_0, ack => cp_elements(807)); -- 
    cp_elements(808) <= cp_elements(805);
    rr_6629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => ptr_deref_1650_load_1_req_0); -- 
    ra_6630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_1_ack_0, ack => cp_elements(809)); -- 
    cp_elements(810) <= cp_elements(805);
    rr_6634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => ptr_deref_1650_load_2_req_0); -- 
    ra_6635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_2_ack_0, ack => cp_elements(811)); -- 
    cp_elements(812) <= cp_elements(805);
    rr_6639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => ptr_deref_1650_load_3_req_0); -- 
    ra_6640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_3_ack_0, ack => cp_elements(813)); -- 
    cpelement_group_814 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(807) & cp_elements(809) & cp_elements(811) & cp_elements(813));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(814),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(815) <= cp_elements(814);
    cr_6650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => ptr_deref_1650_load_0_req_1); -- 
    ca_6651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_0_ack_1, ack => cp_elements(816)); -- 
    cp_elements(817) <= cp_elements(814);
    cr_6655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(817), ack => ptr_deref_1650_load_1_req_1); -- 
    ca_6656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_1_ack_1, ack => cp_elements(818)); -- 
    cp_elements(819) <= cp_elements(814);
    cr_6660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(819), ack => ptr_deref_1650_load_2_req_1); -- 
    ca_6661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_2_ack_1, ack => cp_elements(820)); -- 
    cp_elements(821) <= cp_elements(814);
    cr_6665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(821), ack => ptr_deref_1650_load_3_req_1); -- 
    ca_6666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_load_3_ack_1, ack => cp_elements(822)); -- 
    cpelement_group_823 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(816) & cp_elements(818) & cp_elements(820) & cp_elements(822));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(823),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_6667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(823), ack => ptr_deref_1650_gather_scatter_req_0); -- 
    merge_ack_6668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1650_gather_scatter_ack_0, ack => cp_elements(824)); -- 
    cp_elements(825) <= cp_elements(780);
    cpelement_group_826 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(825) & cp_elements(830));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(826),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_6692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => array_obj_ref_1657_final_reg_req_0); -- 
    cp_elements(827) <= cp_elements(780);
    base_resize_req_6679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => array_obj_ref_1657_base_resize_req_0); -- 
    base_resize_ack_6680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_base_resize_ack_0, ack => cp_elements(828)); -- 
    plus_base_rr_6685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => array_obj_ref_1657_root_address_inst_req_0); -- 
    plus_base_ra_6686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_root_address_inst_ack_0, ack => cp_elements(829)); -- 
    plus_base_cr_6687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(829), ack => array_obj_ref_1657_root_address_inst_req_1); -- 
    plus_base_ca_6688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_root_address_inst_ack_1, ack => cp_elements(830)); -- 
    final_reg_ack_6693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1657_final_reg_ack_0, ack => cp_elements(831)); -- 
    cpelement_group_832 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(831) & cp_elements(833));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(832),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(832), ack => type_cast_1661_inst_req_0); -- 
    cp_elements(833) <= cp_elements(780);
    cp_elements(834) <= type_cast_1661_inst_ack_0;
    cpelement_group_835 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(824) & cp_elements(834) & cp_elements(851));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_6758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(835), ack => ptr_deref_1664_gather_scatter_req_0); -- 
    cp_elements(836) <= cp_elements(834);
    base_resize_req_6717_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(836), ack => ptr_deref_1664_base_resize_req_0); -- 
    base_resize_ack_6718_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_base_resize_ack_0, ack => cp_elements(837)); -- 
    sum_rename_req_6722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(837), ack => ptr_deref_1664_root_address_inst_req_0); -- 
    cp_elements(838) <= ptr_deref_1664_root_address_inst_ack_0;
    cp_elements(839) <= cp_elements(838);
    rr_6730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(839), ack => ptr_deref_1664_addr_0_req_0); -- 
    ra_6731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_0_ack_0, ack => cp_elements(840)); -- 
    cr_6732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => ptr_deref_1664_addr_0_req_1); -- 
    ca_6733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_0_ack_1, ack => cp_elements(841)); -- 
    cp_elements(842) <= cp_elements(838);
    rr_6737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(842), ack => ptr_deref_1664_addr_1_req_0); -- 
    ra_6738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_1_ack_0, ack => cp_elements(843)); -- 
    cr_6739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(843), ack => ptr_deref_1664_addr_1_req_1); -- 
    ca_6740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_1_ack_1, ack => cp_elements(844)); -- 
    cp_elements(845) <= cp_elements(838);
    rr_6744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => ptr_deref_1664_addr_2_req_0); -- 
    ra_6745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_2_ack_0, ack => cp_elements(846)); -- 
    cr_6746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(846), ack => ptr_deref_1664_addr_2_req_1); -- 
    ca_6747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_2_ack_1, ack => cp_elements(847)); -- 
    cp_elements(848) <= cp_elements(838);
    rr_6751_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => ptr_deref_1664_addr_3_req_0); -- 
    ra_6752_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_3_ack_0, ack => cp_elements(849)); -- 
    cr_6753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(849), ack => ptr_deref_1664_addr_3_req_1); -- 
    ca_6754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_addr_3_ack_1, ack => cp_elements(850)); -- 
    cpelement_group_851 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(841) & cp_elements(844) & cp_elements(847) & cp_elements(850));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(851),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(852) <= ptr_deref_1664_gather_scatter_ack_0;
    cp_elements(853) <= cp_elements(852);
    rr_6766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => ptr_deref_1664_store_0_req_0); -- 
    ra_6767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_0_ack_0, ack => cp_elements(854)); -- 
    cp_elements(855) <= cp_elements(852);
    rr_6771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(855), ack => ptr_deref_1664_store_1_req_0); -- 
    ra_6772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_1_ack_0, ack => cp_elements(856)); -- 
    cp_elements(857) <= cp_elements(852);
    rr_6776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => ptr_deref_1664_store_2_req_0); -- 
    ra_6777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_2_ack_0, ack => cp_elements(858)); -- 
    cp_elements(859) <= cp_elements(852);
    rr_6781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(859), ack => ptr_deref_1664_store_3_req_0); -- 
    ra_6782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_3_ack_0, ack => cp_elements(860)); -- 
    cpelement_group_861 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(854) & cp_elements(856) & cp_elements(858) & cp_elements(860));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(861),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(862) <= cp_elements(861);
    cr_6792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(862), ack => ptr_deref_1664_store_0_req_1); -- 
    ca_6793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_0_ack_1, ack => cp_elements(863)); -- 
    cp_elements(864) <= cp_elements(861);
    cr_6797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(864), ack => ptr_deref_1664_store_1_req_1); -- 
    ca_6798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_1_ack_1, ack => cp_elements(865)); -- 
    cp_elements(866) <= cp_elements(861);
    cr_6802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(866), ack => ptr_deref_1664_store_2_req_1); -- 
    ca_6803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_2_ack_1, ack => cp_elements(867)); -- 
    cp_elements(868) <= cp_elements(861);
    cr_6807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => ptr_deref_1664_store_3_req_1); -- 
    ca_6808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1664_store_3_ack_1, ack => cp_elements(869)); -- 
    cpelement_group_870 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(863) & cp_elements(865) & cp_elements(867) & cp_elements(869));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(870),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_871 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(872) & cp_elements(873));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(871),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_6817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => binary_1671_inst_req_0); -- 
    cp_elements(872) <= cp_elements(780);
    cp_elements(873) <= cp_elements(780);
    ra_6818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1671_inst_ack_0, ack => cp_elements(874)); -- 
    cr_6819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => binary_1671_inst_req_1); -- 
    ca_6820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1671_inst_ack_1, ack => cp_elements(875)); -- 
    cpelement_group_876 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(870) & cp_elements(875));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(876),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(877) <= cp_elements(17);
    cp_elements(878) <= false;
    cp_elements(879) <= cp_elements(878);
    cp_elements(880) <= cp_elements(17);
    branch_req_6828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(880), ack => if_stmt_1673_branch_req_0); -- 
    cp_elements(881) <= cp_elements(880);
    cp_elements(882) <= cp_elements(881);
    if_choice_transition_6833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1673_branch_ack_1, ack => cp_elements(883)); -- 
    cp_elements(884) <= cp_elements(881);
    else_choice_transition_6837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1673_branch_ack_0, ack => cp_elements(885)); -- 
    cp_elements(886) <= cp_elements(18);
    cpelement_group_887 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(888) & cp_elements(889));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(887),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(887), ack => type_cast_1682_inst_req_0); -- 
    cp_elements(888) <= cp_elements(886);
    cp_elements(889) <= cp_elements(886);
    ack_6852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1682_inst_ack_0, ack => cp_elements(890)); -- 
    cp_elements(891) <= cp_elements(890);
    cpelement_group_892 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(893) & cp_elements(894));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(892),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_6864_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(892), ack => type_cast_1686_inst_req_0); -- 
    cp_elements(893) <= cp_elements(891);
    cp_elements(894) <= cp_elements(891);
    ack_6865_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1686_inst_ack_0, ack => cp_elements(895)); -- 
    pipe_wreq_6870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(895), ack => simple_obj_ref_1684_inst_req_0); -- 
    pipe_wack_6871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1684_inst_ack_0, ack => cp_elements(896)); -- 
    cp_elements(897) <= false;
    cp_elements(898) <= cp_elements(897);
    cp_elements(899) <= false;
    cp_elements(900) <= cp_elements(899);
    cp_elements(901) <= false;
    cp_elements(902) <= cp_elements(901);
    cp_elements(903) <= false;
    cp_elements(904) <= cp_elements(903);
    cp_elements(905) <= false;
    cp_elements(906) <= cp_elements(905);
    cp_elements(907) <= cp_elements(398);
    cp_elements(908) <= cp_elements(907);
    req_6976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(908), ack => type_cast_1347_inst_req_0); -- 
    ack_6977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1347_inst_ack_0, ack => cp_elements(909)); -- 
    phi_stmt_1341_req_6978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(909), ack => phi_stmt_1341_req_1); -- 
    cp_elements(910) <= cp_elements(907);
    req_6988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(910), ack => type_cast_1340_inst_req_0); -- 
    ack_6989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1340_inst_ack_0, ack => cp_elements(911)); -- 
    phi_stmt_1334_req_6990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => phi_stmt_1334_req_1); -- 
    cpelement_group_912 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(909) & cp_elements(911));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(912),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(913) <= cp_elements(316);
    cp_elements(914) <= cp_elements(913);
    phi_stmt_1341_req_7005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(914), ack => phi_stmt_1341_req_0); -- 
    cp_elements(915) <= cp_elements(913);
    phi_stmt_1334_req_7017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(915), ack => phi_stmt_1334_req_0); -- 
    cpelement_group_916 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(914) & cp_elements(915));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(916),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(917) <= OrReduce(cp_elements(912) & cp_elements(916));
    cp_elements(918) <= cp_elements(917);
    phi_stmt_1334_ack_7022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1334_ack_0, ack => cp_elements(919)); -- 
    phi_stmt_1341_ack_7023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1341_ack_0, ack => cp_elements(920)); -- 
    cpelement_group_921 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(919) & cp_elements(920));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(921),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(922) <= false;
    cp_elements(923) <= cp_elements(922);
    cp_elements(924) <= cp_elements(310);
    cp_elements(925) <= cp_elements(924);
    cp_elements(926) <= cp_elements(925);
    cp_elements(927) <= cp_elements(925);
    req_7053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(927), ack => type_cast_1444_inst_req_0); -- 
    ack_7054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1444_inst_ack_0, ack => cp_elements(928)); -- 
    cpelement_group_929 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(926) & cp_elements(928));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(929),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1439_req_7055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => phi_stmt_1439_req_1); -- 
    cp_elements(930) <= cp_elements(924);
    cp_elements(931) <= cp_elements(930);
    cp_elements(932) <= cp_elements(930);
    req_7070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => type_cast_1438_inst_req_0); -- 
    ack_7071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1438_inst_ack_0, ack => cp_elements(933)); -- 
    cpelement_group_934 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(931) & cp_elements(933));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(934),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1433_req_7072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(934), ack => phi_stmt_1433_req_1); -- 
    cp_elements(935) <= cp_elements(924);
    phi_stmt_1426_req_7084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => phi_stmt_1426_req_1); -- 
    cpelement_group_936 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(929) & cp_elements(934) & cp_elements(935));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(936),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(937) <= cp_elements(417);
    cp_elements(938) <= cp_elements(937);
    cp_elements(939) <= cp_elements(938);
    req_7097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(939), ack => type_cast_1442_inst_req_0); -- 
    ack_7098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1442_inst_ack_0, ack => cp_elements(940)); -- 
    cp_elements(941) <= cp_elements(938);
    cpelement_group_942 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(940) & cp_elements(941));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(942),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1439_req_7104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(942), ack => phi_stmt_1439_req_0); -- 
    cp_elements(943) <= cp_elements(937);
    cp_elements(944) <= cp_elements(943);
    req_7114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => type_cast_1436_inst_req_0); -- 
    ack_7115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1436_inst_ack_0, ack => cp_elements(945)); -- 
    cp_elements(946) <= cp_elements(943);
    cpelement_group_947 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(945) & cp_elements(946));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(947),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1433_req_7121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(947), ack => phi_stmt_1433_req_0); -- 
    cp_elements(948) <= cp_elements(937);
    req_7131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(948), ack => type_cast_1429_inst_req_0); -- 
    ack_7132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1429_inst_ack_0, ack => cp_elements(949)); -- 
    phi_stmt_1426_req_7133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => phi_stmt_1426_req_0); -- 
    cpelement_group_950 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(942) & cp_elements(947) & cp_elements(949));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(950),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(951) <= OrReduce(cp_elements(936) & cp_elements(950));
    cp_elements(952) <= cp_elements(951);
    phi_stmt_1426_ack_7138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1426_ack_0, ack => cp_elements(953)); -- 
    phi_stmt_1433_ack_7139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1433_ack_0, ack => cp_elements(954)); -- 
    phi_stmt_1439_ack_7140_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1439_ack_0, ack => cp_elements(955)); -- 
    cpelement_group_956 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(953) & cp_elements(954) & cp_elements(955));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(956),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(957) <= false;
    cp_elements(958) <= cp_elements(957);
    cp_elements(959) <= cp_elements(432);
    cp_elements(960) <= cp_elements(432);
    req_7170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(960), ack => type_cast_1479_inst_req_0); -- 
    ack_7171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1479_inst_ack_0, ack => cp_elements(961)); -- 
    cpelement_group_962 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(959) & cp_elements(961));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(962),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1474_req_7172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(962), ack => phi_stmt_1474_req_1); -- 
    cp_elements(963) <= cp_elements(448);
    req_7185_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(963), ack => type_cast_1477_inst_req_0); -- 
    ack_7186_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1477_inst_ack_0, ack => cp_elements(964)); -- 
    cp_elements(965) <= cp_elements(448);
    cpelement_group_966 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(964) & cp_elements(965));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(966),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1474_req_7192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(966), ack => phi_stmt_1474_req_0); -- 
    cp_elements(967) <= OrReduce(cp_elements(962) & cp_elements(966));
    cp_elements(968) <= cp_elements(967);
    phi_stmt_1474_ack_7197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1474_ack_0, ack => cp_elements(969)); -- 
    cp_elements(970) <= false;
    cp_elements(971) <= cp_elements(970);
    cp_elements(972) <= false;
    cp_elements(973) <= cp_elements(972);
    cp_elements(974) <= false;
    cp_elements(975) <= cp_elements(974);
    cp_elements(976) <= OrReduce(cp_elements(16) & cp_elements(885));
    cp_elements(977) <= cp_elements(976);
    cp_elements(978) <= OrReduce(cp_elements(156) & cp_elements(228) & cp_elements(257) & cp_elements(295) & cp_elements(495) & cp_elements(883) & cp_elements(896));
    cp_elements(979) <= cp_elements(978);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_1130_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1130_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1130_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1139_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1139_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1139_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1146_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1146_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1146_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1374_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1374_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1374_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1374_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1422_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1422_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1422_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1422_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1540_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1540_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1540_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1554_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1554_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1554_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1554_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1561_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1561_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1561_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1603_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1603_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_1603_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1603_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1612_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1612_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1612_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1627_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1627_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1627_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1642_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1642_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1642_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1657_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1657_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1657_root_address : std_logic_vector(15 downto 0);
    signal binary_1190_wire : std_logic_vector(31 downto 0);
    signal binary_1236_wire : std_logic_vector(31 downto 0);
    signal binary_1270_wire : std_logic_vector(31 downto 0);
    signal binary_1308_wire : std_logic_vector(31 downto 0);
    signal binary_1530_wire : std_logic_vector(31 downto 0);
    signal elt5x_xi11_1617 : std_logic_vector(31 downto 0);
    signal elt5x_xi_1647 : std_logic_vector(31 downto 0);
    signal expr_1189_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1235_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1269_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1307_wire_constant : std_logic_vector(31 downto 0);
    signal expr_1529_wire_constant : std_logic_vector(31 downto 0);
    signal indvarx_xi12x_xi_1334 : std_logic_vector(31 downto 0);
    signal indvarx_xnextx_xi14x_xi_1406 : std_logic_vector(31 downto 0);
    signal orx_xcondx_xi_1296 : std_logic_vector(0 downto 0);
    signal ptr_deref_1134_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1134_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1134_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1134_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1134_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1134_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1150_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1150_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1150_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1150_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1150_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1201_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1201_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1201_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1201_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1201_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1382_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1382_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1382_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1461_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1461_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1461_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1461_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1461_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1543_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1543_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1543_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1543_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1543_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1543_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1564_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1564_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1564_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1564_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1564_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1564_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1606_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1606_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1606_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1606_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1606_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1606_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1620_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1620_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1620_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1620_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1620_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1634_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1634_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1634_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1634_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1634_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1634_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1650_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1650_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1650_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1650_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1650_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1664_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1664_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1664_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1664_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1664_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1664_word_offset_3 : std_logic_vector(15 downto 0);
    signal scevgep12x_xix_xi_1379 : std_logic_vector(31 downto 0);
    signal scevgep14x_xix_xi_1423 : std_logic_vector(31 downto 0);
    signal scevgep_1375 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1118_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1373_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1373_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1421_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1421_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1553_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1553_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1602_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_1602_scaled : std_logic_vector(15 downto 0);
    signal tmp13_1120 : std_logic_vector(31 downto 0);
    signal tmp14_1124 : std_logic_vector(31 downto 0);
    signal tmp15_1131 : std_logic_vector(31 downto 0);
    signal tmp16_1135 : std_logic_vector(31 downto 0);
    signal tmp17_1140 : std_logic_vector(31 downto 0);
    signal tmp17x_xix_xi_1359 : std_logic_vector(31 downto 0);
    signal tmp18_1147 : std_logic_vector(31 downto 0);
    signal tmp19_1151 : std_logic_vector(31 downto 0);
    signal tmp20_1155 : std_logic_vector(31 downto 0);
    signal tmp21_1159 : std_logic_vector(31 downto 0);
    signal tmp22_1164 : std_logic_vector(31 downto 0);
    signal tmp23_1170 : std_logic_vector(31 downto 0);
    signal tmp24_1178 : std_logic_vector(0 downto 0);
    signal tmp25_1198 : std_logic_vector(31 downto 0);
    signal tmp26_1202 : std_logic_vector(31 downto 0);
    signal tmp27_1208 : std_logic_vector(31 downto 0);
    signal tmp28_1214 : std_logic_vector(0 downto 0);
    signal tmp29_1246 : std_logic_vector(31 downto 0);
    signal tmp30_1252 : std_logic_vector(31 downto 0);
    signal tmp31_1258 : std_logic_vector(0 downto 0);
    signal tmp32_1277 : std_logic_vector(15 downto 0);
    signal tmp33_1281 : std_logic_vector(31 downto 0);
    signal tmp34_1286 : std_logic_vector(0 downto 0);
    signal tmp34x_xi_1220 : std_logic_vector(31 downto 0);
    signal tmp35_1291 : std_logic_vector(0 downto 0);
    signal tmp35x_xi_1224 : std_logic_vector(15 downto 0);
    signal tmp36_1318 : std_logic_vector(0 downto 0);
    signal tmp37_1341 : std_logic_vector(31 downto 0);
    signal tmp38_1383 : std_logic_vector(15 downto 0);
    signal tmp39_1387 : std_logic_vector(31 downto 0);
    signal tmp40_1392 : std_logic_vector(31 downto 0);
    signal tmp41_1400 : std_logic_vector(0 downto 0);
    signal tmp42_1451 : std_logic_vector(0 downto 0);
    signal tmp43_1462 : std_logic_vector(7 downto 0);
    signal tmp44_1466 : std_logic_vector(31 downto 0);
    signal tmp45_1471 : std_logic_vector(31 downto 0);
    signal tmp46_1474 : std_logic_vector(31 downto 0);
    signal tmp47_1486 : std_logic_vector(31 downto 0);
    signal tmp48_1492 : std_logic_vector(31 downto 0);
    signal tmp49_1497 : std_logic_vector(31 downto 0);
    signal tmp50_1503 : std_logic_vector(31 downto 0);
    signal tmp51_1508 : std_logic_vector(31 downto 0);
    signal tmp52_1512 : std_logic_vector(15 downto 0);
    signal tmp53_1518 : std_logic_vector(0 downto 0);
    signal tmp54_1541 : std_logic_vector(31 downto 0);
    signal tmp55_1555 : std_logic_vector(31 downto 0);
    signal tmp56_1562 : std_logic_vector(31 downto 0);
    signal tmp57_1571 : std_logic_vector(0 downto 0);
    signal tmp58_1583 : std_logic_vector(31 downto 0);
    signal tmp59_1588 : std_logic_vector(0 downto 0);
    signal tmp5_1331 : std_logic_vector(31 downto 0);
    signal tmp60_1594 : std_logic_vector(31 downto 0);
    signal tmp61_1600 : std_logic_vector(31 downto 0);
    signal tmp62_1604 : std_logic_vector(31 downto 0);
    signal tmp63_1613 : std_logic_vector(31 downto 0);
    signal tmp64_1628 : std_logic_vector(31 downto 0);
    signal tmp65_1632 : std_logic_vector(31 downto 0);
    signal tmp66_1643 : std_logic_vector(31 downto 0);
    signal tmp67_1658 : std_logic_vector(31 downto 0);
    signal tmp68_1662 : std_logic_vector(31 downto 0);
    signal tmp69_1672 : std_logic_vector(0 downto 0);
    signal tmp70_1683 : std_logic_vector(31 downto 0);
    signal tmp8_1371 : std_logic_vector(31 downto 0);
    signal tmp_1354 : std_logic_vector(31 downto 0);
    signal tmpx_xix_xi_1365 : std_logic_vector(31 downto 0);
    signal type_cast_1168_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1173_wire : std_logic_vector(31 downto 0);
    signal type_cast_1176_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1206_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1212_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1218_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1244_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1250_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1256_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1316_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1329_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1338_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1340_wire : std_logic_vector(31 downto 0);
    signal type_cast_1345_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1347_wire : std_logic_vector(31 downto 0);
    signal type_cast_1352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1363_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1369_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1395_wire : std_logic_vector(31 downto 0);
    signal type_cast_1398_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1404_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1417_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1429_wire : std_logic_vector(31 downto 0);
    signal type_cast_1432_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1436_wire : std_logic_vector(31 downto 0);
    signal type_cast_1438_wire : std_logic_vector(31 downto 0);
    signal type_cast_1442_wire : std_logic_vector(31 downto 0);
    signal type_cast_1444_wire : std_logic_vector(31 downto 0);
    signal type_cast_1449_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1477_wire : std_logic_vector(31 downto 0);
    signal type_cast_1479_wire : std_logic_vector(31 downto 0);
    signal type_cast_1484_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1490_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1501_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1516_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_1549_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1597_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1670_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1686_wire : std_logic_vector(31 downto 0);
    signal val6x_xi12_1621 : std_logic_vector(31 downto 0);
    signal val6x_xi_1651 : std_logic_vector(31 downto 0);
    signal xx_xinx_xlcssax_xix_xi_1433 : std_logic_vector(31 downto 0);
    signal xx_xlcssa5x_xix_xi_1426 : std_logic_vector(31 downto 0);
    signal xx_xlcssax_xix_xi_1439 : std_logic_vector(31 downto 0);
    signal xx_xsum20x_xi_1419 : std_logic_vector(31 downto 0);
    signal xx_xsumx_xi_1551 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1130_final_offset <= "0000000000001100";
    array_obj_ref_1139_final_offset <= "0000000000001110";
    array_obj_ref_1146_final_offset <= "0000000000010000";
    array_obj_ref_1374_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1422_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1540_final_offset <= "0000000001010000";
    array_obj_ref_1554_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1561_final_offset <= "0000000001010100";
    array_obj_ref_1603_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_1612_final_offset <= "0000000000011110";
    array_obj_ref_1627_final_offset <= "0000000000011100";
    array_obj_ref_1642_final_offset <= "0000000000011110";
    array_obj_ref_1657_final_offset <= "0000000000011100";
    expr_1189_wire_constant <= "11111111111111111111100000000000";
    expr_1235_wire_constant <= "11111111111111111111100000000000";
    expr_1269_wire_constant <= "11111111111111111111100000000000";
    expr_1307_wire_constant <= "11111111111111111111100000000000";
    expr_1529_wire_constant <= "11111111111111111111100000000000";
    ptr_deref_1134_word_offset_0 <= "0000000000000000";
    ptr_deref_1134_word_offset_1 <= "0000000000000001";
    ptr_deref_1134_word_offset_2 <= "0000000000000010";
    ptr_deref_1134_word_offset_3 <= "0000000000000011";
    ptr_deref_1150_word_offset_0 <= "0000000000000000";
    ptr_deref_1150_word_offset_1 <= "0000000000000001";
    ptr_deref_1150_word_offset_2 <= "0000000000000010";
    ptr_deref_1150_word_offset_3 <= "0000000000000011";
    ptr_deref_1201_word_offset_0 <= "0000000000000000";
    ptr_deref_1201_word_offset_1 <= "0000000000000001";
    ptr_deref_1201_word_offset_2 <= "0000000000000010";
    ptr_deref_1201_word_offset_3 <= "0000000000000011";
    ptr_deref_1382_word_offset_0 <= "0000000000000000";
    ptr_deref_1382_word_offset_1 <= "0000000000000001";
    ptr_deref_1461_word_offset_0 <= "0000000000000000";
    ptr_deref_1543_word_offset_0 <= "0000000000000000";
    ptr_deref_1543_word_offset_1 <= "0000000000000001";
    ptr_deref_1543_word_offset_2 <= "0000000000000010";
    ptr_deref_1543_word_offset_3 <= "0000000000000011";
    ptr_deref_1564_word_offset_0 <= "0000000000000000";
    ptr_deref_1564_word_offset_1 <= "0000000000000001";
    ptr_deref_1564_word_offset_2 <= "0000000000000010";
    ptr_deref_1564_word_offset_3 <= "0000000000000011";
    ptr_deref_1606_word_offset_0 <= "0000000000000000";
    ptr_deref_1606_word_offset_1 <= "0000000000000001";
    ptr_deref_1606_word_offset_2 <= "0000000000000010";
    ptr_deref_1606_word_offset_3 <= "0000000000000011";
    ptr_deref_1620_word_offset_0 <= "0000000000000000";
    ptr_deref_1620_word_offset_1 <= "0000000000000001";
    ptr_deref_1620_word_offset_2 <= "0000000000000010";
    ptr_deref_1620_word_offset_3 <= "0000000000000011";
    ptr_deref_1634_word_offset_0 <= "0000000000000000";
    ptr_deref_1634_word_offset_1 <= "0000000000000001";
    ptr_deref_1634_word_offset_2 <= "0000000000000010";
    ptr_deref_1634_word_offset_3 <= "0000000000000011";
    ptr_deref_1650_word_offset_0 <= "0000000000000000";
    ptr_deref_1650_word_offset_1 <= "0000000000000001";
    ptr_deref_1650_word_offset_2 <= "0000000000000010";
    ptr_deref_1650_word_offset_3 <= "0000000000000011";
    ptr_deref_1664_word_offset_0 <= "0000000000000000";
    ptr_deref_1664_word_offset_1 <= "0000000000000001";
    ptr_deref_1664_word_offset_2 <= "0000000000000010";
    ptr_deref_1664_word_offset_3 <= "0000000000000011";
    type_cast_1168_wire_constant <= "11111111111111111111111111110010";
    type_cast_1176_wire_constant <= "00000000000000000000000000010100";
    type_cast_1206_wire_constant <= "00000000000000000000000011110000";
    type_cast_1212_wire_constant <= "00000000000000000000000001000000";
    type_cast_1218_wire_constant <= "00000000000000000000000000010000";
    type_cast_1244_wire_constant <= "00000000000000000000000000000010";
    type_cast_1250_wire_constant <= "00000000000000000000000000111100";
    type_cast_1256_wire_constant <= "00000000000000000000000000010100";
    type_cast_1316_wire_constant <= "00000000000000000000000000000001";
    type_cast_1329_wire_constant <= "11111111111111111111111111111110";
    type_cast_1338_wire_constant <= "00000000000000000000000000000000";
    type_cast_1345_wire_constant <= "00000000000000000000000000000000";
    type_cast_1352_wire_constant <= "11111111111111111111111111111110";
    type_cast_1363_wire_constant <= "00000000000000000000000000000001";
    type_cast_1369_wire_constant <= "00000000000000000000000000001110";
    type_cast_1398_wire_constant <= "00000000000000000000000000000001";
    type_cast_1404_wire_constant <= "00000000000000000000000000000001";
    type_cast_1417_wire_constant <= "00000000000000000000000000010000";
    type_cast_1432_wire_constant <= "00000000000000000000000000000000";
    type_cast_1449_wire_constant <= "00000000000000000000000000000001";
    type_cast_1484_wire_constant <= "00000000000000001111111111111111";
    type_cast_1490_wire_constant <= "00000000000000000000000000010000";
    type_cast_1501_wire_constant <= "00000000000000000000000000010000";
    type_cast_1516_wire_constant <= "1111111111111111";
    type_cast_1549_wire_constant <= "00000000000000000000000000001110";
    type_cast_1597_wire_constant <= "00000000000000000000000000000000";
    type_cast_1670_wire_constant <= "11111111111111111111111111111111";
    phi_stmt_1334: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1338_wire_constant & type_cast_1340_wire;
      req <= phi_stmt_1334_req_0 & phi_stmt_1334_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1334_ack_0,
          idata => idata,
          odata => indvarx_xi12x_xi_1334,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1334
    phi_stmt_1341: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1345_wire_constant & type_cast_1347_wire;
      req <= phi_stmt_1341_req_0 & phi_stmt_1341_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1341_ack_0,
          idata => idata,
          odata => tmp37_1341,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1341
    phi_stmt_1426: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1429_wire & type_cast_1432_wire_constant;
      req <= phi_stmt_1426_req_0 & phi_stmt_1426_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1426_ack_0,
          idata => idata,
          odata => xx_xlcssa5x_xix_xi_1426,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1426
    phi_stmt_1433: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1436_wire & type_cast_1438_wire;
      req <= phi_stmt_1433_req_0 & phi_stmt_1433_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1433_ack_0,
          idata => idata,
          odata => xx_xinx_xlcssax_xix_xi_1433,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1433
    phi_stmt_1439: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1442_wire & type_cast_1444_wire;
      req <= phi_stmt_1439_req_0 & phi_stmt_1439_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1439_ack_0,
          idata => idata,
          odata => xx_xlcssax_xix_xi_1439,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1439
    phi_stmt_1474: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1477_wire & type_cast_1479_wire;
      req <= phi_stmt_1474_req_0 & phi_stmt_1474_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1474_ack_0,
          idata => idata,
          odata => tmp46_1474,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1474
    ternary_1593_inst: SelectBase generic map(data_width => 32) -- 
      port map( x => tmp22_1164, y => tmp58_1583, sel => tmp59_1588, z => tmp60_1594, req => ternary_1593_inst_req_0, ack => ternary_1593_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1130_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1130_resized_base_address, req => array_obj_ref_1130_base_resize_req_0, ack => array_obj_ref_1130_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1130_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1130_root_address, dout => tmp15_1131, req => array_obj_ref_1130_final_reg_req_0, ack => array_obj_ref_1130_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1139_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1139_resized_base_address, req => array_obj_ref_1139_base_resize_req_0, ack => array_obj_ref_1139_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1139_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1139_root_address, dout => tmp17_1140, req => array_obj_ref_1139_final_reg_req_0, ack => array_obj_ref_1139_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1146_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1146_resized_base_address, req => array_obj_ref_1146_base_resize_req_0, ack => array_obj_ref_1146_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1146_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1146_root_address, dout => tmp18_1147, req => array_obj_ref_1146_final_reg_req_0, ack => array_obj_ref_1146_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1374_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1374_resized_base_address, req => array_obj_ref_1374_base_resize_req_0, ack => array_obj_ref_1374_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1374_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1374_root_address, dout => scevgep_1375, req => array_obj_ref_1374_final_reg_req_0, ack => array_obj_ref_1374_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1374_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_1371, dout => simple_obj_ref_1373_resized, req => array_obj_ref_1374_index_0_resize_req_0, ack => array_obj_ref_1374_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1374_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1373_scaled, dout => array_obj_ref_1374_final_offset, req => array_obj_ref_1374_offset_inst_req_0, ack => array_obj_ref_1374_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1422_resized_base_address, req => array_obj_ref_1422_base_resize_req_0, ack => array_obj_ref_1422_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1422_root_address, dout => scevgep14x_xix_xi_1423, req => array_obj_ref_1422_final_reg_req_0, ack => array_obj_ref_1422_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsum20x_xi_1419, dout => simple_obj_ref_1421_resized, req => array_obj_ref_1422_index_0_resize_req_0, ack => array_obj_ref_1422_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1422_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1421_scaled, dout => array_obj_ref_1422_final_offset, req => array_obj_ref_1422_offset_inst_req_0, ack => array_obj_ref_1422_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1540_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1540_resized_base_address, req => array_obj_ref_1540_base_resize_req_0, ack => array_obj_ref_1540_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1540_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1540_root_address, dout => tmp54_1541, req => array_obj_ref_1540_final_reg_req_0, ack => array_obj_ref_1540_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1554_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1554_resized_base_address, req => array_obj_ref_1554_base_resize_req_0, ack => array_obj_ref_1554_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1554_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1554_root_address, dout => tmp55_1555, req => array_obj_ref_1554_final_reg_req_0, ack => array_obj_ref_1554_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1554_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xsumx_xi_1551, dout => simple_obj_ref_1553_resized, req => array_obj_ref_1554_index_0_resize_req_0, ack => array_obj_ref_1554_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1554_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1553_scaled, dout => array_obj_ref_1554_final_offset, req => array_obj_ref_1554_offset_inst_req_0, ack => array_obj_ref_1554_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1561_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1561_resized_base_address, req => array_obj_ref_1561_base_resize_req_0, ack => array_obj_ref_1561_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1561_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1561_root_address, dout => tmp56_1562, req => array_obj_ref_1561_final_reg_req_0, ack => array_obj_ref_1561_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1603_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp19_1151, dout => array_obj_ref_1603_resized_base_address, req => array_obj_ref_1603_base_resize_req_0, ack => array_obj_ref_1603_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1603_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1603_root_address, dout => tmp62_1604, req => array_obj_ref_1603_final_reg_req_0, ack => array_obj_ref_1603_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1603_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp61_1600, dout => simple_obj_ref_1602_resized, req => array_obj_ref_1603_index_0_resize_req_0, ack => array_obj_ref_1603_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1603_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_1602_scaled, dout => array_obj_ref_1603_final_offset, req => array_obj_ref_1603_offset_inst_req_0, ack => array_obj_ref_1603_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1612_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1612_resized_base_address, req => array_obj_ref_1612_base_resize_req_0, ack => array_obj_ref_1612_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1612_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1612_root_address, dout => tmp63_1613, req => array_obj_ref_1612_final_reg_req_0, ack => array_obj_ref_1612_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1627_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1627_resized_base_address, req => array_obj_ref_1627_base_resize_req_0, ack => array_obj_ref_1627_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1627_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1627_root_address, dout => tmp64_1628, req => array_obj_ref_1627_final_reg_req_0, ack => array_obj_ref_1627_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1642_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1135, dout => array_obj_ref_1642_resized_base_address, req => array_obj_ref_1642_base_resize_req_0, ack => array_obj_ref_1642_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1642_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1642_root_address, dout => tmp66_1643, req => array_obj_ref_1642_final_reg_req_0, ack => array_obj_ref_1642_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1657_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_1124, dout => array_obj_ref_1657_resized_base_address, req => array_obj_ref_1657_base_resize_req_0, ack => array_obj_ref_1657_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1657_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1657_root_address, dout => tmp67_1658, req => array_obj_ref_1657_final_reg_req_0, ack => array_obj_ref_1657_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1134_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp15_1131, dout => ptr_deref_1134_resized_base_address, req => ptr_deref_1134_base_resize_req_0, ack => ptr_deref_1134_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1150_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_1147, dout => ptr_deref_1150_resized_base_address, req => ptr_deref_1150_base_resize_req_0, ack => ptr_deref_1150_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1201_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp25_1198, dout => ptr_deref_1201_resized_base_address, req => ptr_deref_1201_base_resize_req_0, ack => ptr_deref_1201_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1382_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => scevgep12x_xix_xi_1379, dout => ptr_deref_1382_resized_base_address, req => ptr_deref_1382_base_resize_req_0, ack => ptr_deref_1382_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1461_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => xx_xinx_xlcssax_xix_xi_1433, dout => ptr_deref_1461_resized_base_address, req => ptr_deref_1461_base_resize_req_0, ack => ptr_deref_1461_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1543_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp54_1541, dout => ptr_deref_1543_resized_base_address, req => ptr_deref_1543_base_resize_req_0, ack => ptr_deref_1543_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1564_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp56_1562, dout => ptr_deref_1564_resized_base_address, req => ptr_deref_1564_base_resize_req_0, ack => ptr_deref_1564_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1606_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_1147, dout => ptr_deref_1606_resized_base_address, req => ptr_deref_1606_base_resize_req_0, ack => ptr_deref_1606_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1620_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi11_1617, dout => ptr_deref_1620_resized_base_address, req => ptr_deref_1620_base_resize_req_0, ack => ptr_deref_1620_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1634_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp65_1632, dout => ptr_deref_1634_resized_base_address, req => ptr_deref_1634_base_resize_req_0, ack => ptr_deref_1634_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1650_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => elt5x_xi_1647, dout => ptr_deref_1650_resized_base_address, req => ptr_deref_1650_base_resize_req_0, ack => ptr_deref_1650_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1664_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp68_1662, dout => ptr_deref_1664_resized_base_address, req => ptr_deref_1664_base_resize_req_0, ack => ptr_deref_1664_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1119_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1118_wire, dout => tmp13_1120, req => type_cast_1119_inst_req_0, ack => type_cast_1119_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1123_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_1120, dout => tmp14_1124, req => type_cast_1123_inst_req_0, ack => type_cast_1123_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1154_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp19_1151, dout => tmp20_1155, req => type_cast_1154_inst_req_0, ack => type_cast_1154_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1158_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp16_1135, dout => tmp21_1159, req => type_cast_1158_inst_req_0, ack => type_cast_1158_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1173_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp23_1170, dout => type_cast_1173_wire, req => type_cast_1173_inst_req_0, ack => type_cast_1173_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1197_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_1140, dout => tmp25_1198, req => type_cast_1197_inst_req_0, ack => type_cast_1197_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1223_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp34x_xi_1220, dout => tmp35x_xi_1224, req => type_cast_1223_inst_req_0, ack => type_cast_1223_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1280_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp32_1277, dout => tmp33_1281, req => type_cast_1280_inst_req_0, ack => type_cast_1280_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1340_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => indvarx_xnextx_xi14x_xi_1406, dout => type_cast_1340_wire, req => type_cast_1340_inst_req_0, ack => type_cast_1340_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1347_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_1392, dout => type_cast_1347_wire, req => type_cast_1347_inst_req_0, ack => type_cast_1347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1378_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => scevgep_1375, dout => scevgep12x_xix_xi_1379, req => type_cast_1378_inst_req_0, ack => type_cast_1378_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1386_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp38_1383, dout => tmp39_1387, req => type_cast_1386_inst_req_0, ack => type_cast_1386_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1395_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_1359, dout => type_cast_1395_wire, req => type_cast_1395_inst_req_0, ack => type_cast_1395_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1429_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_1392, dout => type_cast_1429_wire, req => type_cast_1429_inst_req_0, ack => type_cast_1429_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1436_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => scevgep14x_xix_xi_1423, dout => type_cast_1436_wire, req => type_cast_1436_inst_req_0, ack => type_cast_1436_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1438_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17_1140, dout => type_cast_1438_wire, req => type_cast_1438_inst_req_0, ack => type_cast_1438_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1442_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp17x_xix_xi_1359, dout => type_cast_1442_wire, req => type_cast_1442_inst_req_0, ack => type_cast_1442_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1444_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp30_1252, dout => type_cast_1444_wire, req => type_cast_1444_inst_req_0, ack => type_cast_1444_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1465_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 32, flow_through => false ) 
      port map( din => tmp43_1462, dout => tmp44_1466, req => type_cast_1465_inst_req_0, ack => type_cast_1465_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1477_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp45_1471, dout => type_cast_1477_wire, req => type_cast_1477_inst_req_0, ack => type_cast_1477_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1479_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => xx_xlcssa5x_xix_xi_1426, dout => type_cast_1479_wire, req => type_cast_1479_inst_req_0, ack => type_cast_1479_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1511_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp51_1508, dout => tmp52_1512, req => type_cast_1511_inst_req_0, ack => type_cast_1511_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1616_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp63_1613, dout => elt5x_xi11_1617, req => type_cast_1616_inst_req_0, ack => type_cast_1616_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1631_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp64_1628, dout => tmp65_1632, req => type_cast_1631_inst_req_0, ack => type_cast_1631_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1646_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp66_1643, dout => elt5x_xi_1647, req => type_cast_1646_inst_req_0, ack => type_cast_1646_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1661_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp67_1658, dout => tmp68_1662, req => type_cast_1661_inst_req_0, ack => type_cast_1661_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1682_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp14_1124, dout => tmp70_1683, req => type_cast_1682_inst_req_0, ack => type_cast_1682_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1686_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp70_1683, dout => type_cast_1686_wire, req => type_cast_1686_inst_req_0, ack => type_cast_1686_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1374_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1374_index_0_rename_ack_0 <= array_obj_ref_1374_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1373_resized;
      simple_obj_ref_1373_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_1422_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1422_index_0_rename_ack_0 <= array_obj_ref_1422_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1421_resized;
      simple_obj_ref_1421_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_1554_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1554_index_0_rename_ack_0 <= array_obj_ref_1554_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1553_resized;
      simple_obj_ref_1553_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_1603_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_1603_index_0_rename_ack_0 <= array_obj_ref_1603_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_1602_resized;
      simple_obj_ref_1602_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1134_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1134_gather_scatter_ack_0 <= ptr_deref_1134_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1134_data_3 & ptr_deref_1134_data_2 & ptr_deref_1134_data_1 & ptr_deref_1134_data_0;
      tmp16_1135 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1134_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1134_root_address_inst_ack_0 <= ptr_deref_1134_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1134_resized_base_address;
      ptr_deref_1134_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1150_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1150_gather_scatter_ack_0 <= ptr_deref_1150_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1150_data_3 & ptr_deref_1150_data_2 & ptr_deref_1150_data_1 & ptr_deref_1150_data_0;
      tmp19_1151 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1150_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1150_root_address_inst_ack_0 <= ptr_deref_1150_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1150_resized_base_address;
      ptr_deref_1150_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1201_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1201_gather_scatter_ack_0 <= ptr_deref_1201_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1201_data_3 & ptr_deref_1201_data_2 & ptr_deref_1201_data_1 & ptr_deref_1201_data_0;
      tmp26_1202 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1201_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1201_root_address_inst_ack_0 <= ptr_deref_1201_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1201_resized_base_address;
      ptr_deref_1201_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1382_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1382_gather_scatter_ack_0 <= ptr_deref_1382_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1382_data_1 & ptr_deref_1382_data_0;
      tmp38_1383 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1382_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1382_root_address_inst_ack_0 <= ptr_deref_1382_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1382_resized_base_address;
      ptr_deref_1382_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1461_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1461_addr_0_ack_0 <= ptr_deref_1461_addr_0_req_0;
      aggregated_sig <= ptr_deref_1461_root_address;
      ptr_deref_1461_word_address_0 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1461_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1461_gather_scatter_ack_0 <= ptr_deref_1461_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1461_data_0;
      tmp43_1462 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1461_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1461_root_address_inst_ack_0 <= ptr_deref_1461_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1461_resized_base_address;
      ptr_deref_1461_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1543_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1543_gather_scatter_ack_0 <= ptr_deref_1543_gather_scatter_req_0;
      aggregated_sig <= tmp17_1140;
      ptr_deref_1543_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1543_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1543_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1543_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1543_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1543_root_address_inst_ack_0 <= ptr_deref_1543_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1543_resized_base_address;
      ptr_deref_1543_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1564_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1564_gather_scatter_ack_0 <= ptr_deref_1564_gather_scatter_req_0;
      aggregated_sig <= tmp55_1555;
      ptr_deref_1564_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1564_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1564_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1564_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1564_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1564_root_address_inst_ack_0 <= ptr_deref_1564_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1564_resized_base_address;
      ptr_deref_1564_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1606_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1606_gather_scatter_ack_0 <= ptr_deref_1606_gather_scatter_req_0;
      aggregated_sig <= tmp62_1604;
      ptr_deref_1606_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1606_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1606_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1606_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1606_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1606_root_address_inst_ack_0 <= ptr_deref_1606_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1606_resized_base_address;
      ptr_deref_1606_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1620_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1620_gather_scatter_ack_0 <= ptr_deref_1620_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1620_data_3 & ptr_deref_1620_data_2 & ptr_deref_1620_data_1 & ptr_deref_1620_data_0;
      val6x_xi12_1621 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1620_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1620_root_address_inst_ack_0 <= ptr_deref_1620_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1620_resized_base_address;
      ptr_deref_1620_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1634_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1634_gather_scatter_ack_0 <= ptr_deref_1634_gather_scatter_req_0;
      aggregated_sig <= val6x_xi12_1621;
      ptr_deref_1634_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1634_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1634_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1634_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1634_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1634_root_address_inst_ack_0 <= ptr_deref_1634_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1634_resized_base_address;
      ptr_deref_1634_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1650_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1650_gather_scatter_ack_0 <= ptr_deref_1650_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1650_data_3 & ptr_deref_1650_data_2 & ptr_deref_1650_data_1 & ptr_deref_1650_data_0;
      val6x_xi_1651 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1650_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1650_root_address_inst_ack_0 <= ptr_deref_1650_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1650_resized_base_address;
      ptr_deref_1650_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1664_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1664_gather_scatter_ack_0 <= ptr_deref_1664_gather_scatter_req_0;
      aggregated_sig <= val6x_xi_1651;
      ptr_deref_1664_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1664_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1664_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1664_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1664_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1664_root_address_inst_ack_0 <= ptr_deref_1664_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1664_resized_base_address;
      ptr_deref_1664_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_1179_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp24_1178;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1179_branch_req_0,
          ack0 => if_stmt_1179_branch_ack_0,
          ack1 => if_stmt_1179_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1225_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp28_1214;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1225_branch_req_0,
          ack0 => if_stmt_1225_branch_ack_0,
          ack1 => if_stmt_1225_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1259_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp31_1258;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1259_branch_req_0,
          ack0 => if_stmt_1259_branch_ack_0,
          ack1 => if_stmt_1259_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1297_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= orx_xcondx_xi_1296;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1297_branch_req_0,
          ack0 => if_stmt_1297_branch_ack_0,
          ack1 => if_stmt_1297_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1319_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp36_1318;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1319_branch_req_0,
          ack0 => if_stmt_1319_branch_ack_0,
          ack1 => if_stmt_1319_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1407_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp41_1400;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1407_branch_req_0,
          ack0 => if_stmt_1407_branch_ack_0,
          ack1 => if_stmt_1407_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1452_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp42_1451;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1452_branch_req_0,
          ack0 => if_stmt_1452_branch_ack_0,
          ack1 => if_stmt_1452_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1519_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp53_1518;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1519_branch_req_0,
          ack0 => if_stmt_1519_branch_ack_0,
          ack1 => if_stmt_1519_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1572_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp57_1571;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1572_branch_req_0,
          ack0 => if_stmt_1572_branch_ack_0,
          ack1 => if_stmt_1572_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1673_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp69_1672;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1673_branch_req_0,
          ack0 => if_stmt_1673_branch_ack_0,
          ack1 => if_stmt_1673_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1130_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1130_resized_base_address;
      array_obj_ref_1130_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1130_root_address_inst_req_0,
          ackL => array_obj_ref_1130_root_address_inst_ack_0,
          reqR => array_obj_ref_1130_root_address_inst_req_1,
          ackR => array_obj_ref_1130_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1139_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1139_resized_base_address;
      array_obj_ref_1139_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1139_root_address_inst_req_0,
          ackL => array_obj_ref_1139_root_address_inst_ack_0,
          reqR => array_obj_ref_1139_root_address_inst_req_1,
          ackR => array_obj_ref_1139_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1146_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1146_resized_base_address;
      array_obj_ref_1146_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1146_root_address_inst_req_0,
          ackL => array_obj_ref_1146_root_address_inst_ack_0,
          reqR => array_obj_ref_1146_root_address_inst_req_1,
          ackR => array_obj_ref_1146_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1374_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1374_final_offset & array_obj_ref_1374_resized_base_address;
      array_obj_ref_1374_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1374_root_address_inst_req_0,
          ackL => array_obj_ref_1374_root_address_inst_ack_0,
          reqR => array_obj_ref_1374_root_address_inst_req_1,
          ackR => array_obj_ref_1374_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1422_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1422_final_offset & array_obj_ref_1422_resized_base_address;
      array_obj_ref_1422_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1422_root_address_inst_req_0,
          ackL => array_obj_ref_1422_root_address_inst_ack_0,
          reqR => array_obj_ref_1422_root_address_inst_req_1,
          ackR => array_obj_ref_1422_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1540_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1540_resized_base_address;
      array_obj_ref_1540_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1540_root_address_inst_req_0,
          ackL => array_obj_ref_1540_root_address_inst_ack_0,
          reqR => array_obj_ref_1540_root_address_inst_req_1,
          ackR => array_obj_ref_1540_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1554_root_address_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1554_final_offset & array_obj_ref_1554_resized_base_address;
      array_obj_ref_1554_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1554_root_address_inst_req_0,
          ackL => array_obj_ref_1554_root_address_inst_ack_0,
          reqR => array_obj_ref_1554_root_address_inst_req_1,
          ackR => array_obj_ref_1554_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1561_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1561_resized_base_address;
      array_obj_ref_1561_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001010100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1561_root_address_inst_req_0,
          ackL => array_obj_ref_1561_root_address_inst_ack_0,
          reqR => array_obj_ref_1561_root_address_inst_req_1,
          ackR => array_obj_ref_1561_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1603_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1603_final_offset & array_obj_ref_1603_resized_base_address;
      array_obj_ref_1603_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1603_root_address_inst_req_0,
          ackL => array_obj_ref_1603_root_address_inst_ack_0,
          reqR => array_obj_ref_1603_root_address_inst_req_1,
          ackR => array_obj_ref_1603_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1612_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1612_resized_base_address;
      array_obj_ref_1612_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1612_root_address_inst_req_0,
          ackL => array_obj_ref_1612_root_address_inst_ack_0,
          reqR => array_obj_ref_1612_root_address_inst_req_1,
          ackR => array_obj_ref_1612_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1627_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1627_resized_base_address;
      array_obj_ref_1627_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1627_root_address_inst_req_0,
          ackL => array_obj_ref_1627_root_address_inst_ack_0,
          reqR => array_obj_ref_1627_root_address_inst_req_1,
          ackR => array_obj_ref_1627_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_1642_root_address_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1642_resized_base_address;
      array_obj_ref_1642_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1642_root_address_inst_req_0,
          ackL => array_obj_ref_1642_root_address_inst_ack_0,
          reqR => array_obj_ref_1642_root_address_inst_req_1,
          ackR => array_obj_ref_1642_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_1657_root_address_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1657_resized_base_address;
      array_obj_ref_1657_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1657_root_address_inst_req_0,
          ackL => array_obj_ref_1657_root_address_inst_ack_0,
          reqR => array_obj_ref_1657_root_address_inst_req_1,
          ackR => array_obj_ref_1657_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_1163_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_1155 & tmp21_1159;
      tmp22_1164 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1163_inst_req_0,
          ackL => binary_1163_inst_ack_0,
          reqR => binary_1163_inst_req_1,
          ackR => binary_1163_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_1169_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp22_1164;
      tmp23_1170 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111110010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1169_inst_req_0,
          ackL => binary_1169_inst_ack_0,
          reqR => binary_1169_inst_req_1,
          ackR => binary_1169_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1177_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1173_wire;
      tmp24_1178 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1177_inst_req_0,
          ackL => binary_1177_inst_ack_0,
          reqR => binary_1177_inst_req_1,
          ackR => binary_1177_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1190_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1120;
      binary_1190_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_1190_inst_req_0,
          ackL => binary_1190_inst_ack_0,
          reqR => binary_1190_inst_req_1,
          ackR => binary_1190_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1207_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_1202;
      tmp27_1208 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000011110000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1207_inst_req_0,
          ackL => binary_1207_inst_ack_0,
          reqR => binary_1207_inst_req_1,
          ackR => binary_1207_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1213_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp27_1208;
      tmp28_1214 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1213_inst_req_0,
          ackL => binary_1213_inst_ack_0,
          reqR => binary_1213_inst_req_1,
          ackR => binary_1213_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1219_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_1202;
      tmp34x_xi_1220 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1219_inst_req_0,
          ackL => binary_1219_inst_ack_0,
          reqR => binary_1219_inst_req_1,
          ackR => binary_1219_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1236_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1120;
      binary_1236_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_1236_inst_req_0,
          ackL => binary_1236_inst_ack_0,
          reqR => binary_1236_inst_req_1,
          ackR => binary_1236_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1245_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp26_1202;
      tmp29_1246 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1245_inst_req_0,
          ackL => binary_1245_inst_ack_0,
          reqR => binary_1245_inst_req_1,
          ackR => binary_1245_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1251_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp29_1246;
      tmp30_1252 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000111100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1251_inst_req_0,
          ackL => binary_1251_inst_ack_0,
          reqR => binary_1251_inst_req_1,
          ackR => binary_1251_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1257_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_1252;
      tmp31_1258 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1257_inst_req_0,
          ackL => binary_1257_inst_ack_0,
          reqR => binary_1257_inst_req_1,
          ackR => binary_1257_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1270_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1120;
      binary_1270_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_1270_inst_req_0,
          ackL => binary_1270_inst_ack_0,
          reqR => binary_1270_inst_req_1,
          ackR => binary_1270_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1285_inst binary_1570_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_1281 & tmp23_1170 & tmp23_1170 & tmp33_1281;
      tmp34_1286 <= data_out(1 downto 1);
      tmp57_1571 <= data_out(0 downto 0);
      reqL(1) <= binary_1285_inst_req_0;
      reqL(0) <= binary_1570_inst_req_0;
      binary_1285_inst_ack_0 <= ackL(1);
      binary_1570_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1285_inst_req_1;
      reqR(0) <= binary_1570_inst_req_1;
      binary_1285_inst_ack_1 <= ackR(1);
      binary_1570_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1290_inst binary_1587_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp33_1281 & tmp30_1252 & tmp22_1164 & tmp58_1583;
      tmp35_1291 <= data_out(1 downto 1);
      tmp59_1588 <= data_out(0 downto 0);
      reqL(1) <= binary_1290_inst_req_0;
      reqL(0) <= binary_1587_inst_req_0;
      binary_1290_inst_ack_0 <= ackL(1);
      binary_1587_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1290_inst_req_1;
      reqR(0) <= binary_1587_inst_req_1;
      binary_1290_inst_ack_1 <= ackR(1);
      binary_1587_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_1295_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp34_1286 & tmp35_1291;
      orx_xcondx_xi_1296 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1295_inst_req_0,
          ackL => binary_1295_inst_ack_0,
          reqR => binary_1295_inst_req_1,
          ackR => binary_1295_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_1308_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1120;
      binary_1308_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_1308_inst_req_0,
          ackL => binary_1308_inst_ack_0,
          reqR => binary_1308_inst_req_1,
          ackR => binary_1308_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_1317_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_1252;
      tmp36_1318 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1317_inst_req_0,
          ackL => binary_1317_inst_ack_0,
          reqR => binary_1317_inst_req_1,
          ackR => binary_1317_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_1330_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_1252;
      tmp5_1331 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1330_inst_req_0,
          ackL => binary_1330_inst_ack_0,
          reqR => binary_1330_inst_req_1,
          ackR => binary_1330_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_1353_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_1334;
      tmp_1354 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1353_inst_req_0,
          ackL => binary_1353_inst_ack_0,
          reqR => binary_1353_inst_req_1,
          ackR => binary_1353_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_1358_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp5_1331 & tmp_1354;
      tmp17x_xix_xi_1359 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1358_inst_req_0,
          ackL => binary_1358_inst_ack_0,
          reqR => binary_1358_inst_req_1,
          ackR => binary_1358_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_1364_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_1334;
      tmpx_xix_xi_1365 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1364_inst_req_0,
          ackL => binary_1364_inst_ack_0,
          reqR => binary_1364_inst_req_1,
          ackR => binary_1364_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_1370_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_1365;
      tmp8_1371 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1370_inst_req_0,
          ackL => binary_1370_inst_ack_0,
          reqR => binary_1370_inst_req_1,
          ackR => binary_1370_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_1391_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp39_1387 & tmp37_1341;
      tmp40_1392 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1391_inst_req_0,
          ackL => binary_1391_inst_ack_0,
          reqR => binary_1391_inst_req_1,
          ackR => binary_1391_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_1399_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1395_wire;
      tmp41_1400 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1399_inst_req_0,
          ackL => binary_1399_inst_ack_0,
          reqR => binary_1399_inst_req_1,
          ackR => binary_1399_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_1405_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xi12x_xi_1334;
      indvarx_xnextx_xi14x_xi_1406 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1405_inst_req_0,
          ackL => binary_1405_inst_ack_0,
          reqR => binary_1405_inst_req_1,
          ackR => binary_1405_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_1418_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmpx_xix_xi_1365;
      xx_xsum20x_xi_1419 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1418_inst_req_0,
          ackL => binary_1418_inst_ack_0,
          reqR => binary_1418_inst_req_1,
          ackR => binary_1418_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_1450_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xlcssax_xix_xi_1439;
      tmp42_1451 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1450_inst_req_0,
          ackL => binary_1450_inst_ack_0,
          reqR => binary_1450_inst_req_1,
          ackR => binary_1450_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_1470_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp44_1466 & xx_xlcssa5x_xix_xi_1426;
      tmp45_1471 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1470_inst_req_0,
          ackL => binary_1470_inst_ack_0,
          reqR => binary_1470_inst_req_1,
          ackR => binary_1470_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_1485_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_1474;
      tmp47_1486 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000001111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1485_inst_req_0,
          ackL => binary_1485_inst_ack_0,
          reqR => binary_1485_inst_req_1,
          ackR => binary_1485_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : binary_1491_inst 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp46_1474;
      tmp48_1492 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1491_inst_req_0,
          ackL => binary_1491_inst_ack_0,
          reqR => binary_1491_inst_req_1,
          ackR => binary_1491_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : binary_1496_inst 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp47_1486 & tmp48_1492;
      tmp49_1497 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1496_inst_req_0,
          ackL => binary_1496_inst_ack_0,
          reqR => binary_1496_inst_req_1,
          ackR => binary_1496_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : binary_1502_inst 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp49_1497;
      tmp50_1503 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1502_inst_req_0,
          ackL => binary_1502_inst_ack_0,
          reqR => binary_1502_inst_req_1,
          ackR => binary_1502_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : binary_1507_inst 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp50_1503 & tmp49_1497;
      tmp51_1508 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1507_inst_req_0,
          ackL => binary_1507_inst_ack_0,
          reqR => binary_1507_inst_req_1,
          ackR => binary_1507_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : binary_1517_inst 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp52_1512;
      tmp53_1518 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "1111111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1517_inst_req_0,
          ackL => binary_1517_inst_ack_0,
          reqR => binary_1517_inst_req_1,
          ackR => binary_1517_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : binary_1530_inst 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp13_1120;
      binary_1530_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_1530_inst_req_0,
          ackL => binary_1530_inst_ack_0,
          reqR => binary_1530_inst_req_1,
          ackR => binary_1530_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : binary_1550_inst 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp30_1252;
      xx_xsumx_xi_1551 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1550_inst_req_0,
          ackL => binary_1550_inst_ack_0,
          reqR => binary_1550_inst_req_1,
          ackR => binary_1550_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : binary_1582_inst 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp23_1170 & tmp33_1281;
      tmp58_1583 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1582_inst_req_0,
          ackL => binary_1582_inst_ack_0,
          reqR => binary_1582_inst_req_1,
          ackR => binary_1582_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : binary_1599_inst 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1597_wire_constant & tmp60_1594;
      tmp61_1600 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1599_inst_req_0,
          ackL => binary_1599_inst_ack_0,
          reqR => binary_1599_inst_req_1,
          ackR => binary_1599_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : binary_1671_inst 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp14_1124;
      tmp69_1672 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1671_inst_req_0,
          ackL => binary_1671_inst_ack_0,
          reqR => binary_1671_inst_req_1,
          ackR => binary_1671_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_1134_addr_0 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1134_root_address;
      ptr_deref_1134_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1134_addr_0_req_0,
          ackL => ptr_deref_1134_addr_0_ack_0,
          reqR => ptr_deref_1134_addr_0_req_1,
          ackR => ptr_deref_1134_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_1134_addr_1 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1134_root_address;
      ptr_deref_1134_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1134_addr_1_req_0,
          ackL => ptr_deref_1134_addr_1_ack_0,
          reqR => ptr_deref_1134_addr_1_req_1,
          ackR => ptr_deref_1134_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_1134_addr_2 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1134_root_address;
      ptr_deref_1134_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1134_addr_2_req_0,
          ackL => ptr_deref_1134_addr_2_ack_0,
          reqR => ptr_deref_1134_addr_2_req_1,
          ackR => ptr_deref_1134_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_1134_addr_3 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1134_root_address;
      ptr_deref_1134_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1134_addr_3_req_0,
          ackL => ptr_deref_1134_addr_3_ack_0,
          reqR => ptr_deref_1134_addr_3_req_1,
          ackR => ptr_deref_1134_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_1150_addr_0 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1150_root_address;
      ptr_deref_1150_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1150_addr_0_req_0,
          ackL => ptr_deref_1150_addr_0_ack_0,
          reqR => ptr_deref_1150_addr_0_req_1,
          ackR => ptr_deref_1150_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_1150_addr_1 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1150_root_address;
      ptr_deref_1150_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1150_addr_1_req_0,
          ackL => ptr_deref_1150_addr_1_ack_0,
          reqR => ptr_deref_1150_addr_1_req_1,
          ackR => ptr_deref_1150_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_1150_addr_2 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1150_root_address;
      ptr_deref_1150_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1150_addr_2_req_0,
          ackL => ptr_deref_1150_addr_2_ack_0,
          reqR => ptr_deref_1150_addr_2_req_1,
          ackR => ptr_deref_1150_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_1150_addr_3 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1150_root_address;
      ptr_deref_1150_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1150_addr_3_req_0,
          ackL => ptr_deref_1150_addr_3_ack_0,
          reqR => ptr_deref_1150_addr_3_req_1,
          ackR => ptr_deref_1150_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_1201_addr_0 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1201_root_address;
      ptr_deref_1201_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1201_addr_0_req_0,
          ackL => ptr_deref_1201_addr_0_ack_0,
          reqR => ptr_deref_1201_addr_0_req_1,
          ackR => ptr_deref_1201_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_1201_addr_1 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1201_root_address;
      ptr_deref_1201_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1201_addr_1_req_0,
          ackL => ptr_deref_1201_addr_1_ack_0,
          reqR => ptr_deref_1201_addr_1_req_1,
          ackR => ptr_deref_1201_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_1201_addr_2 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1201_root_address;
      ptr_deref_1201_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1201_addr_2_req_0,
          ackL => ptr_deref_1201_addr_2_ack_0,
          reqR => ptr_deref_1201_addr_2_req_1,
          ackR => ptr_deref_1201_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_1201_addr_3 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1201_root_address;
      ptr_deref_1201_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1201_addr_3_req_0,
          ackL => ptr_deref_1201_addr_3_ack_0,
          reqR => ptr_deref_1201_addr_3_req_1,
          ackR => ptr_deref_1201_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : ptr_deref_1382_addr_0 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1382_root_address;
      ptr_deref_1382_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1382_addr_0_req_0,
          ackL => ptr_deref_1382_addr_0_ack_0,
          reqR => ptr_deref_1382_addr_0_req_1,
          ackR => ptr_deref_1382_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : ptr_deref_1382_addr_1 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1382_root_address;
      ptr_deref_1382_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1382_addr_1_req_0,
          ackL => ptr_deref_1382_addr_1_ack_0,
          reqR => ptr_deref_1382_addr_1_req_1,
          ackR => ptr_deref_1382_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : ptr_deref_1543_addr_0 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1543_root_address;
      ptr_deref_1543_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1543_addr_0_req_0,
          ackL => ptr_deref_1543_addr_0_ack_0,
          reqR => ptr_deref_1543_addr_0_req_1,
          ackR => ptr_deref_1543_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : ptr_deref_1543_addr_1 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1543_root_address;
      ptr_deref_1543_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1543_addr_1_req_0,
          ackL => ptr_deref_1543_addr_1_ack_0,
          reqR => ptr_deref_1543_addr_1_req_1,
          ackR => ptr_deref_1543_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : ptr_deref_1543_addr_2 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1543_root_address;
      ptr_deref_1543_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1543_addr_2_req_0,
          ackL => ptr_deref_1543_addr_2_ack_0,
          reqR => ptr_deref_1543_addr_2_req_1,
          ackR => ptr_deref_1543_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : ptr_deref_1543_addr_3 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1543_root_address;
      ptr_deref_1543_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1543_addr_3_req_0,
          ackL => ptr_deref_1543_addr_3_ack_0,
          reqR => ptr_deref_1543_addr_3_req_1,
          ackR => ptr_deref_1543_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : ptr_deref_1564_addr_0 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1564_root_address;
      ptr_deref_1564_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1564_addr_0_req_0,
          ackL => ptr_deref_1564_addr_0_ack_0,
          reqR => ptr_deref_1564_addr_0_req_1,
          ackR => ptr_deref_1564_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : ptr_deref_1564_addr_1 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1564_root_address;
      ptr_deref_1564_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1564_addr_1_req_0,
          ackL => ptr_deref_1564_addr_1_ack_0,
          reqR => ptr_deref_1564_addr_1_req_1,
          ackR => ptr_deref_1564_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : ptr_deref_1564_addr_2 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1564_root_address;
      ptr_deref_1564_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1564_addr_2_req_0,
          ackL => ptr_deref_1564_addr_2_ack_0,
          reqR => ptr_deref_1564_addr_2_req_1,
          ackR => ptr_deref_1564_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : ptr_deref_1564_addr_3 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1564_root_address;
      ptr_deref_1564_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1564_addr_3_req_0,
          ackL => ptr_deref_1564_addr_3_ack_0,
          reqR => ptr_deref_1564_addr_3_req_1,
          ackR => ptr_deref_1564_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : ptr_deref_1606_addr_0 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1606_root_address;
      ptr_deref_1606_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1606_addr_0_req_0,
          ackL => ptr_deref_1606_addr_0_ack_0,
          reqR => ptr_deref_1606_addr_0_req_1,
          ackR => ptr_deref_1606_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : ptr_deref_1606_addr_1 
    SplitOperatorGroup75: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1606_root_address;
      ptr_deref_1606_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1606_addr_1_req_0,
          ackL => ptr_deref_1606_addr_1_ack_0,
          reqR => ptr_deref_1606_addr_1_req_1,
          ackR => ptr_deref_1606_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : ptr_deref_1606_addr_2 
    SplitOperatorGroup76: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1606_root_address;
      ptr_deref_1606_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1606_addr_2_req_0,
          ackL => ptr_deref_1606_addr_2_ack_0,
          reqR => ptr_deref_1606_addr_2_req_1,
          ackR => ptr_deref_1606_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : ptr_deref_1606_addr_3 
    SplitOperatorGroup77: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1606_root_address;
      ptr_deref_1606_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1606_addr_3_req_0,
          ackL => ptr_deref_1606_addr_3_ack_0,
          reqR => ptr_deref_1606_addr_3_req_1,
          ackR => ptr_deref_1606_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared split operator group (78) : ptr_deref_1620_addr_0 
    SplitOperatorGroup78: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1620_root_address;
      ptr_deref_1620_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1620_addr_0_req_0,
          ackL => ptr_deref_1620_addr_0_ack_0,
          reqR => ptr_deref_1620_addr_0_req_1,
          ackR => ptr_deref_1620_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 78
    -- shared split operator group (79) : ptr_deref_1620_addr_1 
    SplitOperatorGroup79: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1620_root_address;
      ptr_deref_1620_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1620_addr_1_req_0,
          ackL => ptr_deref_1620_addr_1_ack_0,
          reqR => ptr_deref_1620_addr_1_req_1,
          ackR => ptr_deref_1620_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 79
    -- shared split operator group (80) : ptr_deref_1620_addr_2 
    SplitOperatorGroup80: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1620_root_address;
      ptr_deref_1620_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1620_addr_2_req_0,
          ackL => ptr_deref_1620_addr_2_ack_0,
          reqR => ptr_deref_1620_addr_2_req_1,
          ackR => ptr_deref_1620_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 80
    -- shared split operator group (81) : ptr_deref_1620_addr_3 
    SplitOperatorGroup81: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1620_root_address;
      ptr_deref_1620_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1620_addr_3_req_0,
          ackL => ptr_deref_1620_addr_3_ack_0,
          reqR => ptr_deref_1620_addr_3_req_1,
          ackR => ptr_deref_1620_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 81
    -- shared split operator group (82) : ptr_deref_1634_addr_0 
    SplitOperatorGroup82: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1634_root_address;
      ptr_deref_1634_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1634_addr_0_req_0,
          ackL => ptr_deref_1634_addr_0_ack_0,
          reqR => ptr_deref_1634_addr_0_req_1,
          ackR => ptr_deref_1634_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 82
    -- shared split operator group (83) : ptr_deref_1634_addr_1 
    SplitOperatorGroup83: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1634_root_address;
      ptr_deref_1634_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1634_addr_1_req_0,
          ackL => ptr_deref_1634_addr_1_ack_0,
          reqR => ptr_deref_1634_addr_1_req_1,
          ackR => ptr_deref_1634_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 83
    -- shared split operator group (84) : ptr_deref_1634_addr_2 
    SplitOperatorGroup84: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1634_root_address;
      ptr_deref_1634_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1634_addr_2_req_0,
          ackL => ptr_deref_1634_addr_2_ack_0,
          reqR => ptr_deref_1634_addr_2_req_1,
          ackR => ptr_deref_1634_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 84
    -- shared split operator group (85) : ptr_deref_1634_addr_3 
    SplitOperatorGroup85: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1634_root_address;
      ptr_deref_1634_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1634_addr_3_req_0,
          ackL => ptr_deref_1634_addr_3_ack_0,
          reqR => ptr_deref_1634_addr_3_req_1,
          ackR => ptr_deref_1634_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 85
    -- shared split operator group (86) : ptr_deref_1650_addr_0 
    SplitOperatorGroup86: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1650_root_address;
      ptr_deref_1650_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1650_addr_0_req_0,
          ackL => ptr_deref_1650_addr_0_ack_0,
          reqR => ptr_deref_1650_addr_0_req_1,
          ackR => ptr_deref_1650_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 86
    -- shared split operator group (87) : ptr_deref_1650_addr_1 
    SplitOperatorGroup87: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1650_root_address;
      ptr_deref_1650_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1650_addr_1_req_0,
          ackL => ptr_deref_1650_addr_1_ack_0,
          reqR => ptr_deref_1650_addr_1_req_1,
          ackR => ptr_deref_1650_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 87
    -- shared split operator group (88) : ptr_deref_1650_addr_2 
    SplitOperatorGroup88: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1650_root_address;
      ptr_deref_1650_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1650_addr_2_req_0,
          ackL => ptr_deref_1650_addr_2_ack_0,
          reqR => ptr_deref_1650_addr_2_req_1,
          ackR => ptr_deref_1650_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 88
    -- shared split operator group (89) : ptr_deref_1650_addr_3 
    SplitOperatorGroup89: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1650_root_address;
      ptr_deref_1650_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1650_addr_3_req_0,
          ackL => ptr_deref_1650_addr_3_ack_0,
          reqR => ptr_deref_1650_addr_3_req_1,
          ackR => ptr_deref_1650_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 89
    -- shared split operator group (90) : ptr_deref_1664_addr_0 
    SplitOperatorGroup90: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1664_root_address;
      ptr_deref_1664_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1664_addr_0_req_0,
          ackL => ptr_deref_1664_addr_0_ack_0,
          reqR => ptr_deref_1664_addr_0_req_1,
          ackR => ptr_deref_1664_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 90
    -- shared split operator group (91) : ptr_deref_1664_addr_1 
    SplitOperatorGroup91: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1664_root_address;
      ptr_deref_1664_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1664_addr_1_req_0,
          ackL => ptr_deref_1664_addr_1_ack_0,
          reqR => ptr_deref_1664_addr_1_req_1,
          ackR => ptr_deref_1664_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 91
    -- shared split operator group (92) : ptr_deref_1664_addr_2 
    SplitOperatorGroup92: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1664_root_address;
      ptr_deref_1664_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1664_addr_2_req_0,
          ackL => ptr_deref_1664_addr_2_ack_0,
          reqR => ptr_deref_1664_addr_2_req_1,
          ackR => ptr_deref_1664_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 92
    -- shared split operator group (93) : ptr_deref_1664_addr_3 
    SplitOperatorGroup93: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1664_root_address;
      ptr_deref_1664_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1664_addr_3_req_0,
          ackL => ptr_deref_1664_addr_3_ack_0,
          reqR => ptr_deref_1664_addr_3_req_1,
          ackR => ptr_deref_1664_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 93
    -- shared load operator group (0) : ptr_deref_1150_load_3 ptr_deref_1150_load_2 ptr_deref_1134_load_2 ptr_deref_1150_load_1 ptr_deref_1150_load_0 ptr_deref_1201_load_2 ptr_deref_1134_load_1 ptr_deref_1134_load_0 ptr_deref_1134_load_3 ptr_deref_1201_load_3 ptr_deref_1461_load_0 ptr_deref_1620_load_0 ptr_deref_1382_load_1 ptr_deref_1382_load_0 ptr_deref_1201_load_1 ptr_deref_1201_load_0 ptr_deref_1620_load_1 ptr_deref_1620_load_2 ptr_deref_1620_load_3 ptr_deref_1650_load_0 ptr_deref_1650_load_1 ptr_deref_1650_load_2 ptr_deref_1650_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(367 downto 0);
      signal data_out: std_logic_vector(183 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 22 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1150_load_3_req_0,
        ptr_deref_1150_load_3_ack_0,
        ptr_deref_1150_load_3_req_1,
        ptr_deref_1150_load_3_ack_1,
        "ptr_deref_1150_load_3",
        "memory_space_5" ,
        ptr_deref_1150_data_3,
        ptr_deref_1150_word_address_3,
        "ptr_deref_1150_data_3",
        "ptr_deref_1150_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1150_load_2_req_0,
        ptr_deref_1150_load_2_ack_0,
        ptr_deref_1150_load_2_req_1,
        ptr_deref_1150_load_2_ack_1,
        "ptr_deref_1150_load_2",
        "memory_space_5" ,
        ptr_deref_1150_data_2,
        ptr_deref_1150_word_address_2,
        "ptr_deref_1150_data_2",
        "ptr_deref_1150_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1134_load_2_req_0,
        ptr_deref_1134_load_2_ack_0,
        ptr_deref_1134_load_2_req_1,
        ptr_deref_1134_load_2_ack_1,
        "ptr_deref_1134_load_2",
        "memory_space_5" ,
        ptr_deref_1134_data_2,
        ptr_deref_1134_word_address_2,
        "ptr_deref_1134_data_2",
        "ptr_deref_1134_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1150_load_1_req_0,
        ptr_deref_1150_load_1_ack_0,
        ptr_deref_1150_load_1_req_1,
        ptr_deref_1150_load_1_ack_1,
        "ptr_deref_1150_load_1",
        "memory_space_5" ,
        ptr_deref_1150_data_1,
        ptr_deref_1150_word_address_1,
        "ptr_deref_1150_data_1",
        "ptr_deref_1150_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1150_load_0_req_0,
        ptr_deref_1150_load_0_ack_0,
        ptr_deref_1150_load_0_req_1,
        ptr_deref_1150_load_0_ack_1,
        "ptr_deref_1150_load_0",
        "memory_space_5" ,
        ptr_deref_1150_data_0,
        ptr_deref_1150_word_address_0,
        "ptr_deref_1150_data_0",
        "ptr_deref_1150_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1201_load_2_req_0,
        ptr_deref_1201_load_2_ack_0,
        ptr_deref_1201_load_2_req_1,
        ptr_deref_1201_load_2_ack_1,
        "ptr_deref_1201_load_2",
        "memory_space_5" ,
        ptr_deref_1201_data_2,
        ptr_deref_1201_word_address_2,
        "ptr_deref_1201_data_2",
        "ptr_deref_1201_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1134_load_1_req_0,
        ptr_deref_1134_load_1_ack_0,
        ptr_deref_1134_load_1_req_1,
        ptr_deref_1134_load_1_ack_1,
        "ptr_deref_1134_load_1",
        "memory_space_5" ,
        ptr_deref_1134_data_1,
        ptr_deref_1134_word_address_1,
        "ptr_deref_1134_data_1",
        "ptr_deref_1134_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1134_load_0_req_0,
        ptr_deref_1134_load_0_ack_0,
        ptr_deref_1134_load_0_req_1,
        ptr_deref_1134_load_0_ack_1,
        "ptr_deref_1134_load_0",
        "memory_space_5" ,
        ptr_deref_1134_data_0,
        ptr_deref_1134_word_address_0,
        "ptr_deref_1134_data_0",
        "ptr_deref_1134_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1134_load_3_req_0,
        ptr_deref_1134_load_3_ack_0,
        ptr_deref_1134_load_3_req_1,
        ptr_deref_1134_load_3_ack_1,
        "ptr_deref_1134_load_3",
        "memory_space_5" ,
        ptr_deref_1134_data_3,
        ptr_deref_1134_word_address_3,
        "ptr_deref_1134_data_3",
        "ptr_deref_1134_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1201_load_3_req_0,
        ptr_deref_1201_load_3_ack_0,
        ptr_deref_1201_load_3_req_1,
        ptr_deref_1201_load_3_ack_1,
        "ptr_deref_1201_load_3",
        "memory_space_5" ,
        ptr_deref_1201_data_3,
        ptr_deref_1201_word_address_3,
        "ptr_deref_1201_data_3",
        "ptr_deref_1201_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1461_load_0_req_0,
        ptr_deref_1461_load_0_ack_0,
        ptr_deref_1461_load_0_req_1,
        ptr_deref_1461_load_0_ack_1,
        "ptr_deref_1461_load_0",
        "memory_space_5" ,
        ptr_deref_1461_data_0,
        ptr_deref_1461_word_address_0,
        "ptr_deref_1461_data_0",
        "ptr_deref_1461_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1620_load_0_req_0,
        ptr_deref_1620_load_0_ack_0,
        ptr_deref_1620_load_0_req_1,
        ptr_deref_1620_load_0_ack_1,
        "ptr_deref_1620_load_0",
        "memory_space_5" ,
        ptr_deref_1620_data_0,
        ptr_deref_1620_word_address_0,
        "ptr_deref_1620_data_0",
        "ptr_deref_1620_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1382_load_1_req_0,
        ptr_deref_1382_load_1_ack_0,
        ptr_deref_1382_load_1_req_1,
        ptr_deref_1382_load_1_ack_1,
        "ptr_deref_1382_load_1",
        "memory_space_5" ,
        ptr_deref_1382_data_1,
        ptr_deref_1382_word_address_1,
        "ptr_deref_1382_data_1",
        "ptr_deref_1382_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1382_load_0_req_0,
        ptr_deref_1382_load_0_ack_0,
        ptr_deref_1382_load_0_req_1,
        ptr_deref_1382_load_0_ack_1,
        "ptr_deref_1382_load_0",
        "memory_space_5" ,
        ptr_deref_1382_data_0,
        ptr_deref_1382_word_address_0,
        "ptr_deref_1382_data_0",
        "ptr_deref_1382_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1201_load_1_req_0,
        ptr_deref_1201_load_1_ack_0,
        ptr_deref_1201_load_1_req_1,
        ptr_deref_1201_load_1_ack_1,
        "ptr_deref_1201_load_1",
        "memory_space_5" ,
        ptr_deref_1201_data_1,
        ptr_deref_1201_word_address_1,
        "ptr_deref_1201_data_1",
        "ptr_deref_1201_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1201_load_0_req_0,
        ptr_deref_1201_load_0_ack_0,
        ptr_deref_1201_load_0_req_1,
        ptr_deref_1201_load_0_ack_1,
        "ptr_deref_1201_load_0",
        "memory_space_5" ,
        ptr_deref_1201_data_0,
        ptr_deref_1201_word_address_0,
        "ptr_deref_1201_data_0",
        "ptr_deref_1201_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1620_load_1_req_0,
        ptr_deref_1620_load_1_ack_0,
        ptr_deref_1620_load_1_req_1,
        ptr_deref_1620_load_1_ack_1,
        "ptr_deref_1620_load_1",
        "memory_space_5" ,
        ptr_deref_1620_data_1,
        ptr_deref_1620_word_address_1,
        "ptr_deref_1620_data_1",
        "ptr_deref_1620_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1620_load_2_req_0,
        ptr_deref_1620_load_2_ack_0,
        ptr_deref_1620_load_2_req_1,
        ptr_deref_1620_load_2_ack_1,
        "ptr_deref_1620_load_2",
        "memory_space_5" ,
        ptr_deref_1620_data_2,
        ptr_deref_1620_word_address_2,
        "ptr_deref_1620_data_2",
        "ptr_deref_1620_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1620_load_3_req_0,
        ptr_deref_1620_load_3_ack_0,
        ptr_deref_1620_load_3_req_1,
        ptr_deref_1620_load_3_ack_1,
        "ptr_deref_1620_load_3",
        "memory_space_5" ,
        ptr_deref_1620_data_3,
        ptr_deref_1620_word_address_3,
        "ptr_deref_1620_data_3",
        "ptr_deref_1620_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1650_load_0_req_0,
        ptr_deref_1650_load_0_ack_0,
        ptr_deref_1650_load_0_req_1,
        ptr_deref_1650_load_0_ack_1,
        "ptr_deref_1650_load_0",
        "memory_space_5" ,
        ptr_deref_1650_data_0,
        ptr_deref_1650_word_address_0,
        "ptr_deref_1650_data_0",
        "ptr_deref_1650_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1650_load_1_req_0,
        ptr_deref_1650_load_1_ack_0,
        ptr_deref_1650_load_1_req_1,
        ptr_deref_1650_load_1_ack_1,
        "ptr_deref_1650_load_1",
        "memory_space_5" ,
        ptr_deref_1650_data_1,
        ptr_deref_1650_word_address_1,
        "ptr_deref_1650_data_1",
        "ptr_deref_1650_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1650_load_2_req_0,
        ptr_deref_1650_load_2_ack_0,
        ptr_deref_1650_load_2_req_1,
        ptr_deref_1650_load_2_ack_1,
        "ptr_deref_1650_load_2",
        "memory_space_5" ,
        ptr_deref_1650_data_2,
        ptr_deref_1650_word_address_2,
        "ptr_deref_1650_data_2",
        "ptr_deref_1650_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1650_load_3_req_0,
        ptr_deref_1650_load_3_ack_0,
        ptr_deref_1650_load_3_req_1,
        ptr_deref_1650_load_3_ack_1,
        "ptr_deref_1650_load_3",
        "memory_space_5" ,
        ptr_deref_1650_data_3,
        ptr_deref_1650_word_address_3,
        "ptr_deref_1650_data_3",
        "ptr_deref_1650_word_address_3" -- 
      );
      reqL(22) <= ptr_deref_1150_load_3_req_0;
      reqL(21) <= ptr_deref_1150_load_2_req_0;
      reqL(20) <= ptr_deref_1134_load_2_req_0;
      reqL(19) <= ptr_deref_1150_load_1_req_0;
      reqL(18) <= ptr_deref_1150_load_0_req_0;
      reqL(17) <= ptr_deref_1201_load_2_req_0;
      reqL(16) <= ptr_deref_1134_load_1_req_0;
      reqL(15) <= ptr_deref_1134_load_0_req_0;
      reqL(14) <= ptr_deref_1134_load_3_req_0;
      reqL(13) <= ptr_deref_1201_load_3_req_0;
      reqL(12) <= ptr_deref_1461_load_0_req_0;
      reqL(11) <= ptr_deref_1620_load_0_req_0;
      reqL(10) <= ptr_deref_1382_load_1_req_0;
      reqL(9) <= ptr_deref_1382_load_0_req_0;
      reqL(8) <= ptr_deref_1201_load_1_req_0;
      reqL(7) <= ptr_deref_1201_load_0_req_0;
      reqL(6) <= ptr_deref_1620_load_1_req_0;
      reqL(5) <= ptr_deref_1620_load_2_req_0;
      reqL(4) <= ptr_deref_1620_load_3_req_0;
      reqL(3) <= ptr_deref_1650_load_0_req_0;
      reqL(2) <= ptr_deref_1650_load_1_req_0;
      reqL(1) <= ptr_deref_1650_load_2_req_0;
      reqL(0) <= ptr_deref_1650_load_3_req_0;
      ptr_deref_1150_load_3_ack_0 <= ackL(22);
      ptr_deref_1150_load_2_ack_0 <= ackL(21);
      ptr_deref_1134_load_2_ack_0 <= ackL(20);
      ptr_deref_1150_load_1_ack_0 <= ackL(19);
      ptr_deref_1150_load_0_ack_0 <= ackL(18);
      ptr_deref_1201_load_2_ack_0 <= ackL(17);
      ptr_deref_1134_load_1_ack_0 <= ackL(16);
      ptr_deref_1134_load_0_ack_0 <= ackL(15);
      ptr_deref_1134_load_3_ack_0 <= ackL(14);
      ptr_deref_1201_load_3_ack_0 <= ackL(13);
      ptr_deref_1461_load_0_ack_0 <= ackL(12);
      ptr_deref_1620_load_0_ack_0 <= ackL(11);
      ptr_deref_1382_load_1_ack_0 <= ackL(10);
      ptr_deref_1382_load_0_ack_0 <= ackL(9);
      ptr_deref_1201_load_1_ack_0 <= ackL(8);
      ptr_deref_1201_load_0_ack_0 <= ackL(7);
      ptr_deref_1620_load_1_ack_0 <= ackL(6);
      ptr_deref_1620_load_2_ack_0 <= ackL(5);
      ptr_deref_1620_load_3_ack_0 <= ackL(4);
      ptr_deref_1650_load_0_ack_0 <= ackL(3);
      ptr_deref_1650_load_1_ack_0 <= ackL(2);
      ptr_deref_1650_load_2_ack_0 <= ackL(1);
      ptr_deref_1650_load_3_ack_0 <= ackL(0);
      reqR(22) <= ptr_deref_1150_load_3_req_1;
      reqR(21) <= ptr_deref_1150_load_2_req_1;
      reqR(20) <= ptr_deref_1134_load_2_req_1;
      reqR(19) <= ptr_deref_1150_load_1_req_1;
      reqR(18) <= ptr_deref_1150_load_0_req_1;
      reqR(17) <= ptr_deref_1201_load_2_req_1;
      reqR(16) <= ptr_deref_1134_load_1_req_1;
      reqR(15) <= ptr_deref_1134_load_0_req_1;
      reqR(14) <= ptr_deref_1134_load_3_req_1;
      reqR(13) <= ptr_deref_1201_load_3_req_1;
      reqR(12) <= ptr_deref_1461_load_0_req_1;
      reqR(11) <= ptr_deref_1620_load_0_req_1;
      reqR(10) <= ptr_deref_1382_load_1_req_1;
      reqR(9) <= ptr_deref_1382_load_0_req_1;
      reqR(8) <= ptr_deref_1201_load_1_req_1;
      reqR(7) <= ptr_deref_1201_load_0_req_1;
      reqR(6) <= ptr_deref_1620_load_1_req_1;
      reqR(5) <= ptr_deref_1620_load_2_req_1;
      reqR(4) <= ptr_deref_1620_load_3_req_1;
      reqR(3) <= ptr_deref_1650_load_0_req_1;
      reqR(2) <= ptr_deref_1650_load_1_req_1;
      reqR(1) <= ptr_deref_1650_load_2_req_1;
      reqR(0) <= ptr_deref_1650_load_3_req_1;
      ptr_deref_1150_load_3_ack_1 <= ackR(22);
      ptr_deref_1150_load_2_ack_1 <= ackR(21);
      ptr_deref_1134_load_2_ack_1 <= ackR(20);
      ptr_deref_1150_load_1_ack_1 <= ackR(19);
      ptr_deref_1150_load_0_ack_1 <= ackR(18);
      ptr_deref_1201_load_2_ack_1 <= ackR(17);
      ptr_deref_1134_load_1_ack_1 <= ackR(16);
      ptr_deref_1134_load_0_ack_1 <= ackR(15);
      ptr_deref_1134_load_3_ack_1 <= ackR(14);
      ptr_deref_1201_load_3_ack_1 <= ackR(13);
      ptr_deref_1461_load_0_ack_1 <= ackR(12);
      ptr_deref_1620_load_0_ack_1 <= ackR(11);
      ptr_deref_1382_load_1_ack_1 <= ackR(10);
      ptr_deref_1382_load_0_ack_1 <= ackR(9);
      ptr_deref_1201_load_1_ack_1 <= ackR(8);
      ptr_deref_1201_load_0_ack_1 <= ackR(7);
      ptr_deref_1620_load_1_ack_1 <= ackR(6);
      ptr_deref_1620_load_2_ack_1 <= ackR(5);
      ptr_deref_1620_load_3_ack_1 <= ackR(4);
      ptr_deref_1650_load_0_ack_1 <= ackR(3);
      ptr_deref_1650_load_1_ack_1 <= ackR(2);
      ptr_deref_1650_load_2_ack_1 <= ackR(1);
      ptr_deref_1650_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_1150_word_address_3 & ptr_deref_1150_word_address_2 & ptr_deref_1134_word_address_2 & ptr_deref_1150_word_address_1 & ptr_deref_1150_word_address_0 & ptr_deref_1201_word_address_2 & ptr_deref_1134_word_address_1 & ptr_deref_1134_word_address_0 & ptr_deref_1134_word_address_3 & ptr_deref_1201_word_address_3 & ptr_deref_1461_word_address_0 & ptr_deref_1620_word_address_0 & ptr_deref_1382_word_address_1 & ptr_deref_1382_word_address_0 & ptr_deref_1201_word_address_1 & ptr_deref_1201_word_address_0 & ptr_deref_1620_word_address_1 & ptr_deref_1620_word_address_2 & ptr_deref_1620_word_address_3 & ptr_deref_1650_word_address_0 & ptr_deref_1650_word_address_1 & ptr_deref_1650_word_address_2 & ptr_deref_1650_word_address_3;
      ptr_deref_1150_data_3 <= data_out(183 downto 176);
      ptr_deref_1150_data_2 <= data_out(175 downto 168);
      ptr_deref_1134_data_2 <= data_out(167 downto 160);
      ptr_deref_1150_data_1 <= data_out(159 downto 152);
      ptr_deref_1150_data_0 <= data_out(151 downto 144);
      ptr_deref_1201_data_2 <= data_out(143 downto 136);
      ptr_deref_1134_data_1 <= data_out(135 downto 128);
      ptr_deref_1134_data_0 <= data_out(127 downto 120);
      ptr_deref_1134_data_3 <= data_out(119 downto 112);
      ptr_deref_1201_data_3 <= data_out(111 downto 104);
      ptr_deref_1461_data_0 <= data_out(103 downto 96);
      ptr_deref_1620_data_0 <= data_out(95 downto 88);
      ptr_deref_1382_data_1 <= data_out(87 downto 80);
      ptr_deref_1382_data_0 <= data_out(79 downto 72);
      ptr_deref_1201_data_1 <= data_out(71 downto 64);
      ptr_deref_1201_data_0 <= data_out(63 downto 56);
      ptr_deref_1620_data_1 <= data_out(55 downto 48);
      ptr_deref_1620_data_2 <= data_out(47 downto 40);
      ptr_deref_1620_data_3 <= data_out(39 downto 32);
      ptr_deref_1650_data_0 <= data_out(31 downto 24);
      ptr_deref_1650_data_1 <= data_out(23 downto 16);
      ptr_deref_1650_data_2 <= data_out(15 downto 8);
      ptr_deref_1650_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 23,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 23,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_1564_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1564_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1564_word_address_0) &  " data ptr_deref_1564_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1564_data_0) severity note; --
        end if;
        if ptr_deref_1543_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1543_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1543_word_address_3) &  " data ptr_deref_1543_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1543_data_3) severity note; --
        end if;
        if ptr_deref_1543_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1543_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1543_word_address_2) &  " data ptr_deref_1543_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1543_data_2) severity note; --
        end if;
        if ptr_deref_1543_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1543_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1543_word_address_1) &  " data ptr_deref_1543_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1543_data_1) severity note; --
        end if;
        if ptr_deref_1543_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1543_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1543_word_address_0) &  " data ptr_deref_1543_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1543_data_0) severity note; --
        end if;
        if ptr_deref_1564_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1564_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1564_word_address_3) &  " data ptr_deref_1564_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1564_data_3) severity note; --
        end if;
        if ptr_deref_1564_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1564_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1564_word_address_2) &  " data ptr_deref_1564_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1564_data_2) severity note; --
        end if;
        if ptr_deref_1606_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1606_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1606_word_address_3) &  " data ptr_deref_1606_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1606_data_3) severity note; --
        end if;
        if ptr_deref_1606_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1606_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1606_word_address_2) &  " data ptr_deref_1606_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1606_data_2) severity note; --
        end if;
        if ptr_deref_1606_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1606_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1606_word_address_1) &  " data ptr_deref_1606_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1606_data_1) severity note; --
        end if;
        if ptr_deref_1564_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1564_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1564_word_address_1) &  " data ptr_deref_1564_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1564_data_1) severity note; --
        end if;
        if ptr_deref_1606_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1606_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1606_word_address_0) &  " data ptr_deref_1606_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1606_data_0) severity note; --
        end if;
        if ptr_deref_1634_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1634_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1634_word_address_0) &  " data ptr_deref_1634_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1634_data_0) severity note; --
        end if;
        if ptr_deref_1634_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1634_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1634_word_address_1) &  " data ptr_deref_1634_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1634_data_1) severity note; --
        end if;
        if ptr_deref_1634_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1634_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1634_word_address_2) &  " data ptr_deref_1634_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1634_data_2) severity note; --
        end if;
        if ptr_deref_1634_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1634_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1634_word_address_3) &  " data ptr_deref_1634_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1634_data_3) severity note; --
        end if;
        if ptr_deref_1664_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1664_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1664_word_address_0) &  " data ptr_deref_1664_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1664_data_0) severity note; --
        end if;
        if ptr_deref_1664_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1664_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1664_word_address_1) &  " data ptr_deref_1664_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1664_data_1) severity note; --
        end if;
        if ptr_deref_1664_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1664_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1664_word_address_2) &  " data ptr_deref_1664_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1664_data_2) severity note; --
        end if;
        if ptr_deref_1664_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_1664_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1664_word_address_3) &  " data ptr_deref_1664_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1664_data_3) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1564_store_0 ptr_deref_1543_store_3 ptr_deref_1543_store_2 ptr_deref_1543_store_1 ptr_deref_1543_store_0 ptr_deref_1564_store_3 ptr_deref_1564_store_2 ptr_deref_1606_store_3 ptr_deref_1606_store_2 ptr_deref_1606_store_1 ptr_deref_1564_store_1 ptr_deref_1606_store_0 ptr_deref_1634_store_0 ptr_deref_1634_store_1 ptr_deref_1634_store_2 ptr_deref_1634_store_3 ptr_deref_1664_store_0 ptr_deref_1664_store_1 ptr_deref_1664_store_2 ptr_deref_1664_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(319 downto 0);
      signal data_in: std_logic_vector(159 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 19 downto 0);
      -- 
    begin -- 
      reqL(19) <= ptr_deref_1564_store_0_req_0;
      reqL(18) <= ptr_deref_1543_store_3_req_0;
      reqL(17) <= ptr_deref_1543_store_2_req_0;
      reqL(16) <= ptr_deref_1543_store_1_req_0;
      reqL(15) <= ptr_deref_1543_store_0_req_0;
      reqL(14) <= ptr_deref_1564_store_3_req_0;
      reqL(13) <= ptr_deref_1564_store_2_req_0;
      reqL(12) <= ptr_deref_1606_store_3_req_0;
      reqL(11) <= ptr_deref_1606_store_2_req_0;
      reqL(10) <= ptr_deref_1606_store_1_req_0;
      reqL(9) <= ptr_deref_1564_store_1_req_0;
      reqL(8) <= ptr_deref_1606_store_0_req_0;
      reqL(7) <= ptr_deref_1634_store_0_req_0;
      reqL(6) <= ptr_deref_1634_store_1_req_0;
      reqL(5) <= ptr_deref_1634_store_2_req_0;
      reqL(4) <= ptr_deref_1634_store_3_req_0;
      reqL(3) <= ptr_deref_1664_store_0_req_0;
      reqL(2) <= ptr_deref_1664_store_1_req_0;
      reqL(1) <= ptr_deref_1664_store_2_req_0;
      reqL(0) <= ptr_deref_1664_store_3_req_0;
      ptr_deref_1564_store_0_ack_0 <= ackL(19);
      ptr_deref_1543_store_3_ack_0 <= ackL(18);
      ptr_deref_1543_store_2_ack_0 <= ackL(17);
      ptr_deref_1543_store_1_ack_0 <= ackL(16);
      ptr_deref_1543_store_0_ack_0 <= ackL(15);
      ptr_deref_1564_store_3_ack_0 <= ackL(14);
      ptr_deref_1564_store_2_ack_0 <= ackL(13);
      ptr_deref_1606_store_3_ack_0 <= ackL(12);
      ptr_deref_1606_store_2_ack_0 <= ackL(11);
      ptr_deref_1606_store_1_ack_0 <= ackL(10);
      ptr_deref_1564_store_1_ack_0 <= ackL(9);
      ptr_deref_1606_store_0_ack_0 <= ackL(8);
      ptr_deref_1634_store_0_ack_0 <= ackL(7);
      ptr_deref_1634_store_1_ack_0 <= ackL(6);
      ptr_deref_1634_store_2_ack_0 <= ackL(5);
      ptr_deref_1634_store_3_ack_0 <= ackL(4);
      ptr_deref_1664_store_0_ack_0 <= ackL(3);
      ptr_deref_1664_store_1_ack_0 <= ackL(2);
      ptr_deref_1664_store_2_ack_0 <= ackL(1);
      ptr_deref_1664_store_3_ack_0 <= ackL(0);
      reqR(19) <= ptr_deref_1564_store_0_req_1;
      reqR(18) <= ptr_deref_1543_store_3_req_1;
      reqR(17) <= ptr_deref_1543_store_2_req_1;
      reqR(16) <= ptr_deref_1543_store_1_req_1;
      reqR(15) <= ptr_deref_1543_store_0_req_1;
      reqR(14) <= ptr_deref_1564_store_3_req_1;
      reqR(13) <= ptr_deref_1564_store_2_req_1;
      reqR(12) <= ptr_deref_1606_store_3_req_1;
      reqR(11) <= ptr_deref_1606_store_2_req_1;
      reqR(10) <= ptr_deref_1606_store_1_req_1;
      reqR(9) <= ptr_deref_1564_store_1_req_1;
      reqR(8) <= ptr_deref_1606_store_0_req_1;
      reqR(7) <= ptr_deref_1634_store_0_req_1;
      reqR(6) <= ptr_deref_1634_store_1_req_1;
      reqR(5) <= ptr_deref_1634_store_2_req_1;
      reqR(4) <= ptr_deref_1634_store_3_req_1;
      reqR(3) <= ptr_deref_1664_store_0_req_1;
      reqR(2) <= ptr_deref_1664_store_1_req_1;
      reqR(1) <= ptr_deref_1664_store_2_req_1;
      reqR(0) <= ptr_deref_1664_store_3_req_1;
      ptr_deref_1564_store_0_ack_1 <= ackR(19);
      ptr_deref_1543_store_3_ack_1 <= ackR(18);
      ptr_deref_1543_store_2_ack_1 <= ackR(17);
      ptr_deref_1543_store_1_ack_1 <= ackR(16);
      ptr_deref_1543_store_0_ack_1 <= ackR(15);
      ptr_deref_1564_store_3_ack_1 <= ackR(14);
      ptr_deref_1564_store_2_ack_1 <= ackR(13);
      ptr_deref_1606_store_3_ack_1 <= ackR(12);
      ptr_deref_1606_store_2_ack_1 <= ackR(11);
      ptr_deref_1606_store_1_ack_1 <= ackR(10);
      ptr_deref_1564_store_1_ack_1 <= ackR(9);
      ptr_deref_1606_store_0_ack_1 <= ackR(8);
      ptr_deref_1634_store_0_ack_1 <= ackR(7);
      ptr_deref_1634_store_1_ack_1 <= ackR(6);
      ptr_deref_1634_store_2_ack_1 <= ackR(5);
      ptr_deref_1634_store_3_ack_1 <= ackR(4);
      ptr_deref_1664_store_0_ack_1 <= ackR(3);
      ptr_deref_1664_store_1_ack_1 <= ackR(2);
      ptr_deref_1664_store_2_ack_1 <= ackR(1);
      ptr_deref_1664_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1564_word_address_0 & ptr_deref_1543_word_address_3 & ptr_deref_1543_word_address_2 & ptr_deref_1543_word_address_1 & ptr_deref_1543_word_address_0 & ptr_deref_1564_word_address_3 & ptr_deref_1564_word_address_2 & ptr_deref_1606_word_address_3 & ptr_deref_1606_word_address_2 & ptr_deref_1606_word_address_1 & ptr_deref_1564_word_address_1 & ptr_deref_1606_word_address_0 & ptr_deref_1634_word_address_0 & ptr_deref_1634_word_address_1 & ptr_deref_1634_word_address_2 & ptr_deref_1634_word_address_3 & ptr_deref_1664_word_address_0 & ptr_deref_1664_word_address_1 & ptr_deref_1664_word_address_2 & ptr_deref_1664_word_address_3;
      data_in <= ptr_deref_1564_data_0 & ptr_deref_1543_data_3 & ptr_deref_1543_data_2 & ptr_deref_1543_data_1 & ptr_deref_1543_data_0 & ptr_deref_1564_data_3 & ptr_deref_1564_data_2 & ptr_deref_1606_data_3 & ptr_deref_1606_data_2 & ptr_deref_1606_data_1 & ptr_deref_1564_data_1 & ptr_deref_1606_data_0 & ptr_deref_1634_data_0 & ptr_deref_1634_data_1 & ptr_deref_1634_data_2 & ptr_deref_1634_data_3 & ptr_deref_1664_data_0 & ptr_deref_1664_data_1 & ptr_deref_1664_data_2 & ptr_deref_1664_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 20,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 20,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_1118_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1118_inst_ack_0 then -- 
            assert false report " ReadPipe chk_in0 to wire simple_obj_ref_1118_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1118_inst_req_0;
      simple_obj_ref_1118_inst_ack_0 <= ack(0);
      simple_obj_ref_1118_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => chk_in0_pipe_read_req(0),
          oack => chk_in0_pipe_read_ack(0),
          odata => chk_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1267_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_1270_wire value="  &  convert_slv_to_hex_string(binary_1270_wire) severity note; --
        end if;
        if simple_obj_ref_1305_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_1308_wire value="  &  convert_slv_to_hex_string(binary_1308_wire) severity note; --
        end if;
        if simple_obj_ref_1233_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_1236_wire value="  &  convert_slv_to_hex_string(binary_1236_wire) severity note; --
        end if;
        if simple_obj_ref_1527_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_1530_wire value="  &  convert_slv_to_hex_string(binary_1530_wire) severity note; --
        end if;
        if simple_obj_ref_1187_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_1190_wire value="  &  convert_slv_to_hex_string(binary_1190_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_1267_inst simple_obj_ref_1305_inst simple_obj_ref_1233_inst simple_obj_ref_1527_inst simple_obj_ref_1187_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(159 downto 0);
      signal req, ack : BooleanArray( 4 downto 0);
      -- 
    begin -- 
      req(4) <= simple_obj_ref_1267_inst_req_0;
      req(3) <= simple_obj_ref_1305_inst_req_0;
      req(2) <= simple_obj_ref_1233_inst_req_0;
      req(1) <= simple_obj_ref_1527_inst_req_0;
      req(0) <= simple_obj_ref_1187_inst_req_0;
      simple_obj_ref_1267_inst_ack_0 <= ack(4);
      simple_obj_ref_1305_inst_ack_0 <= ack(3);
      simple_obj_ref_1233_inst_ack_0 <= ack(2);
      simple_obj_ref_1527_inst_ack_0 <= ack(1);
      simple_obj_ref_1187_inst_ack_0 <= ack(0);
      data_in <= binary_1270_wire & binary_1308_wire & binary_1236_wire & binary_1530_wire & binary_1190_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 5,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1684_inst_ack_0 then -- 
          assert false report " WritePipe rtt_in0 from wire type_cast_1686_wire value="  &  convert_slv_to_hex_string(type_cast_1686_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_1684_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_1684_inst_req_0;
      simple_obj_ref_1684_inst_ack_0 <= ack(0);
      data_in <= type_cast_1686_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => rtt_in0_pipe_write_req(0),
          oack => rtt_in0_pipe_write_ack(0),
          odata => rtt_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_1277_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_1277_call_req_0;
      call_stmt_1277_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_1277_call_req_1;
      call_stmt_1277_call_ack_1 <= ackR(0);
      data_in <= tmp35x_xi_1224;
      tmp32_1277 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 16,
        owidth => 16,
        twidth => 2,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 16, twidth => 2, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_rtt is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(4 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_lr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_3_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
    memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_3_sr_tag :  out  std_logic_vector(7 downto 0);
    memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
    memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
    memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    rtt_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    to0_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to0_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to0_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to1_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to1_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to1_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to2_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to2_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to2_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    to3_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    to3_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    to3_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_rtt;
architecture Default of ahir_glue_rtt is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_rtt_CP_7287_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_1888_index_0_scale_req_0 : boolean;
  signal binary_1823_inst_ack_1 : boolean;
  signal ptr_deref_1869_load_0_ack_1 : boolean;
  signal type_cast_1788_inst_ack_0 : boolean;
  signal binary_1823_inst_req_0 : boolean;
  signal binary_1761_inst_ack_1 : boolean;
  signal binary_1823_inst_req_1 : boolean;
  signal if_stmt_1877_branch_ack_0 : boolean;
  signal binary_1761_inst_ack_0 : boolean;
  signal ptr_deref_1869_root_address_inst_ack_0 : boolean;
  signal type_cast_1788_inst_req_0 : boolean;
  signal binary_1761_inst_req_1 : boolean;
  signal binary_1807_inst_req_0 : boolean;
  signal ptr_deref_1869_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_1825_gather_scatter_ack_0 : boolean;
  signal if_stmt_1763_branch_req_0 : boolean;
  signal ptr_deref_2042_load_0_req_0 : boolean;
  signal if_stmt_1763_branch_ack_0 : boolean;
  signal ptr_deref_1869_gather_scatter_req_0 : boolean;
  signal ptr_deref_1869_load_0_ack_0 : boolean;
  signal ptr_deref_1869_load_0_req_0 : boolean;
  signal simple_obj_ref_1825_store_0_ack_0 : boolean;
  signal addr_of_1889_final_reg_req_0 : boolean;
  signal ptr_deref_2042_load_1_req_1 : boolean;
  signal binary_1761_inst_req_0 : boolean;
  signal ptr_deref_1869_load_0_req_1 : boolean;
  signal simple_obj_ref_1825_gather_scatter_req_0 : boolean;
  signal binary_1792_inst_ack_1 : boolean;
  signal ptr_deref_1869_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_1825_store_0_req_0 : boolean;
  signal binary_1823_inst_ack_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_req_0 : boolean;
  signal binary_1792_inst_req_1 : boolean;
  signal array_obj_ref_1888_index_0_scale_ack_0 : boolean;
  signal binary_1755_inst_ack_1 : boolean;
  signal array_obj_ref_1888_offset_inst_ack_0 : boolean;
  signal ptr_deref_2046_load_3_ack_0 : boolean;
  signal ptr_deref_1869_addr_0_req_0 : boolean;
  signal ptr_deref_2042_load_1_ack_1 : boolean;
  signal ptr_deref_2042_load_0_ack_0 : boolean;
  signal binary_1834_inst_req_1 : boolean;
  signal ptr_deref_1869_addr_0_ack_0 : boolean;
  signal if_stmt_1763_branch_ack_1 : boolean;
  signal array_obj_ref_1888_index_0_scale_req_1 : boolean;
  signal binary_1875_inst_req_1 : boolean;
  signal array_obj_ref_1937_offset_inst_ack_0 : boolean;
  signal binary_1792_inst_ack_0 : boolean;
  signal array_obj_ref_1888_index_0_scale_ack_1 : boolean;
  signal if_stmt_1794_branch_req_0 : boolean;
  signal array_obj_ref_1888_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1888_index_sum_1_ack_0 : boolean;
  signal if_stmt_1794_branch_ack_1 : boolean;
  signal binary_1792_inst_req_0 : boolean;
  signal ptr_deref_2046_load_3_req_0 : boolean;
  signal array_obj_ref_1888_index_sum_1_req_1 : boolean;
  signal binary_1875_inst_ack_1 : boolean;
  signal if_stmt_1925_branch_req_0 : boolean;
  signal array_obj_ref_1888_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1888_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1888_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1869_base_resize_req_0 : boolean;
  signal array_obj_ref_1888_offset_inst_req_0 : boolean;
  signal ptr_deref_1869_base_resize_ack_0 : boolean;
  signal if_stmt_1794_branch_ack_0 : boolean;
  signal binary_1834_inst_ack_1 : boolean;
  signal binary_1755_inst_req_1 : boolean;
  signal if_stmt_1912_branch_ack_1 : boolean;
  signal binary_1755_inst_req_0 : boolean;
  signal simple_obj_ref_1817_gather_scatter_ack_0 : boolean;
  signal binary_1807_inst_ack_1 : boolean;
  signal simple_obj_ref_1697_inst_ack_0 : boolean;
  signal simple_obj_ref_1697_inst_req_0 : boolean;
  signal array_obj_ref_1709_final_reg_ack_0 : boolean;
  signal array_obj_ref_1888_index_0_resize_ack_0 : boolean;
  signal binary_1875_inst_ack_0 : boolean;
  signal binary_1774_inst_req_0 : boolean;
  signal binary_1755_inst_ack_0 : boolean;
  signal array_obj_ref_1709_root_address_inst_req_0 : boolean;
  signal binary_1834_inst_req_0 : boolean;
  signal simple_obj_ref_1825_store_0_ack_1 : boolean;
  signal simple_obj_ref_1817_load_0_req_0 : boolean;
  signal ptr_deref_2046_load_1_req_0 : boolean;
  signal binary_1875_inst_req_0 : boolean;
  signal simple_obj_ref_1825_store_0_req_1 : boolean;
  signal type_cast_1702_inst_req_0 : boolean;
  signal type_cast_1698_inst_ack_0 : boolean;
  signal array_obj_ref_1864_index_0_scale_ack_1 : boolean;
  signal ptr_deref_1717_addr_3_ack_1 : boolean;
  signal binary_1807_inst_req_1 : boolean;
  signal array_obj_ref_1864_index_sum_1_req_0 : boolean;
  signal ptr_deref_1717_addr_2_req_1 : boolean;
  signal ptr_deref_1717_addr_2_ack_1 : boolean;
  signal type_cast_1702_inst_ack_0 : boolean;
  signal addr_of_1889_final_reg_ack_0 : boolean;
  signal array_obj_ref_1709_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1709_base_resize_req_0 : boolean;
  signal binary_1834_inst_ack_0 : boolean;
  signal array_obj_ref_1937_base_resize_req_0 : boolean;
  signal array_obj_ref_1709_base_resize_ack_0 : boolean;
  signal ptr_deref_2046_load_2_ack_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_ack_0 : boolean;
  signal binary_1904_inst_ack_0 : boolean;
  signal binary_1807_inst_ack_0 : boolean;
  signal if_stmt_1912_branch_req_0 : boolean;
  signal if_stmt_1877_branch_ack_1 : boolean;
  signal ptr_deref_2046_load_1_ack_0 : boolean;
  signal type_cast_1803_inst_req_0 : boolean;
  signal array_obj_ref_1864_index_sum_1_ack_1 : boolean;
  signal ptr_deref_1717_addr_1_req_0 : boolean;
  signal addr_of_1865_final_reg_ack_0 : boolean;
  signal array_obj_ref_1864_root_address_inst_req_0 : boolean;
  signal ptr_deref_1717_base_resize_req_0 : boolean;
  signal type_cast_1803_inst_ack_0 : boolean;
  signal addr_of_1865_final_reg_req_0 : boolean;
  signal type_cast_1713_inst_req_0 : boolean;
  signal ptr_deref_2046_base_resize_req_0 : boolean;
  signal simple_obj_ref_1817_load_0_ack_1 : boolean;
  signal ptr_deref_1717_addr_1_ack_0 : boolean;
  signal array_obj_ref_1864_index_sum_1_req_1 : boolean;
  signal ptr_deref_1717_addr_1_req_1 : boolean;
  signal array_obj_ref_1709_final_reg_req_0 : boolean;
  signal type_cast_1713_inst_ack_0 : boolean;
  signal binary_1923_inst_req_1 : boolean;
  signal array_obj_ref_1864_offset_inst_req_0 : boolean;
  signal ptr_deref_1717_addr_0_ack_1 : boolean;
  signal ptr_deref_1717_addr_2_req_0 : boolean;
  signal array_obj_ref_1864_index_sum_1_ack_0 : boolean;
  signal ptr_deref_1717_addr_2_ack_0 : boolean;
  signal ptr_deref_1717_base_resize_ack_0 : boolean;
  signal simple_obj_ref_1817_load_0_req_1 : boolean;
  signal type_cast_1698_inst_req_0 : boolean;
  signal ptr_deref_1717_root_address_inst_req_0 : boolean;
  signal type_cast_1830_inst_ack_0 : boolean;
  signal simple_obj_ref_1817_load_0_ack_0 : boolean;
  signal array_obj_ref_1709_root_address_inst_ack_1 : boolean;
  signal ptr_deref_1717_addr_3_ack_0 : boolean;
  signal ptr_deref_1717_addr_3_req_1 : boolean;
  signal ptr_deref_1717_addr_1_ack_1 : boolean;
  signal array_obj_ref_1709_root_address_inst_req_1 : boolean;
  signal if_stmt_1912_branch_ack_0 : boolean;
  signal ptr_deref_1717_addr_3_req_0 : boolean;
  signal ptr_deref_1717_load_1_ack_0 : boolean;
  signal ptr_deref_1717_load_2_req_0 : boolean;
  signal array_obj_ref_1864_index_0_scale_req_0 : boolean;
  signal ptr_deref_1717_load_2_ack_0 : boolean;
  signal ptr_deref_1717_addr_0_ack_0 : boolean;
  signal array_obj_ref_1864_offset_inst_ack_0 : boolean;
  signal ptr_deref_1717_addr_0_req_1 : boolean;
  signal binary_1923_inst_ack_1 : boolean;
  signal ptr_deref_1717_load_3_req_0 : boolean;
  signal ptr_deref_1717_load_3_ack_0 : boolean;
  signal ptr_deref_1717_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_1817_gather_scatter_req_0 : boolean;
  signal array_obj_ref_1864_index_0_scale_ack_0 : boolean;
  signal ptr_deref_1717_load_1_req_0 : boolean;
  signal ptr_deref_1717_addr_0_req_0 : boolean;
  signal type_cast_1830_inst_req_0 : boolean;
  signal ptr_deref_1717_load_0_req_0 : boolean;
  signal array_obj_ref_1864_index_0_scale_req_1 : boolean;
  signal ptr_deref_1717_load_0_ack_0 : boolean;
  signal binary_1910_inst_req_1 : boolean;
  signal binary_1910_inst_ack_1 : boolean;
  signal binary_1904_inst_ack_1 : boolean;
  signal binary_1923_inst_ack_0 : boolean;
  signal ptr_deref_1717_load_0_req_1 : boolean;
  signal array_obj_ref_1864_index_0_resize_ack_0 : boolean;
  signal ptr_deref_1717_load_0_ack_1 : boolean;
  signal binary_1910_inst_ack_0 : boolean;
  signal ptr_deref_1940_store_0_ack_0 : boolean;
  signal ptr_deref_1940_store_0_req_1 : boolean;
  signal ptr_deref_1940_store_0_ack_1 : boolean;
  signal ptr_deref_1940_base_resize_req_0 : boolean;
  signal ptr_deref_1940_base_resize_ack_0 : boolean;
  signal ptr_deref_1940_root_address_inst_req_0 : boolean;
  signal ptr_deref_1940_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1940_addr_0_req_0 : boolean;
  signal ptr_deref_1940_addr_0_ack_0 : boolean;
  signal ptr_deref_1940_gather_scatter_req_0 : boolean;
  signal ptr_deref_1940_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1940_store_0_req_0 : boolean;
  signal if_stmt_1925_branch_ack_0 : boolean;
  signal ptr_deref_2042_load_3_ack_0 : boolean;
  signal array_obj_ref_1937_root_address_inst_ack_0 : boolean;
  signal if_stmt_1925_branch_ack_1 : boolean;
  signal binary_1904_inst_req_1 : boolean;
  signal ptr_deref_2046_base_resize_ack_0 : boolean;
  signal binary_1774_inst_ack_0 : boolean;
  signal array_obj_ref_1937_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1937_root_address_inst_ack_1 : boolean;
  signal if_stmt_1836_branch_req_0 : boolean;
  signal array_obj_ref_1937_final_reg_req_0 : boolean;
  signal array_obj_ref_1937_final_reg_ack_0 : boolean;
  signal phi_stmt_1845_req_1 : boolean;
  signal array_obj_ref_1937_root_address_inst_req_0 : boolean;
  signal ptr_deref_1717_load_1_req_1 : boolean;
  signal array_obj_ref_1864_index_0_resize_req_0 : boolean;
  signal ptr_deref_1717_load_1_ack_1 : boolean;
  signal ptr_deref_1717_load_2_req_1 : boolean;
  signal ptr_deref_1717_load_2_ack_1 : boolean;
  signal binary_1923_inst_req_0 : boolean;
  signal ptr_deref_1717_load_3_req_1 : boolean;
  signal ptr_deref_1717_load_3_ack_1 : boolean;
  signal ptr_deref_2046_addr_2_req_1 : boolean;
  signal ptr_deref_1717_gather_scatter_req_0 : boolean;
  signal ptr_deref_1717_gather_scatter_ack_0 : boolean;
  signal binary_1910_inst_req_0 : boolean;
  signal if_stmt_1877_branch_req_0 : boolean;
  signal ptr_deref_2046_addr_3_ack_1 : boolean;
  signal ptr_deref_2046_load_0_req_0 : boolean;
  signal ptr_deref_2046_load_1_req_1 : boolean;
  signal if_stmt_1809_branch_ack_0 : boolean;
  signal if_stmt_1809_branch_ack_1 : boolean;
  signal binary_1904_inst_req_0 : boolean;
  signal binary_1774_inst_ack_1 : boolean;
  signal array_obj_ref_1937_offset_inst_req_0 : boolean;
  signal array_obj_ref_1727_index_0_resize_req_0 : boolean;
  signal if_stmt_1836_branch_ack_0 : boolean;
  signal array_obj_ref_1727_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_1937_base_resize_ack_0 : boolean;
  signal binary_1774_inst_req_1 : boolean;
  signal array_obj_ref_1727_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1727_index_0_scale_ack_0 : boolean;
  signal if_stmt_1809_branch_req_0 : boolean;
  signal array_obj_ref_1727_index_0_scale_req_1 : boolean;
  signal if_stmt_1836_branch_ack_1 : boolean;
  signal array_obj_ref_1727_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_1727_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1727_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1727_index_sum_1_req_1 : boolean;
  signal array_obj_ref_1727_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_1727_offset_inst_req_0 : boolean;
  signal array_obj_ref_1727_offset_inst_ack_0 : boolean;
  signal array_obj_ref_1727_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1727_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2046_load_2_ack_1 : boolean;
  signal ptr_deref_2046_load_2_req_1 : boolean;
  signal addr_of_1728_final_reg_req_0 : boolean;
  signal addr_of_1728_final_reg_ack_0 : boolean;
  signal ptr_deref_2046_load_0_req_1 : boolean;
  signal ptr_deref_2046_addr_2_ack_1 : boolean;
  signal ptr_deref_2046_load_0_ack_1 : boolean;
  signal ptr_deref_2046_load_2_req_0 : boolean;
  signal ptr_deref_2046_root_address_inst_req_0 : boolean;
  signal ptr_deref_2042_load_2_req_1 : boolean;
  signal ptr_deref_2046_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2042_load_2_ack_1 : boolean;
  signal array_obj_ref_1736_index_0_resize_req_0 : boolean;
  signal array_obj_ref_1736_index_0_resize_ack_0 : boolean;
  signal ptr_deref_2046_load_1_ack_1 : boolean;
  signal array_obj_ref_1736_index_0_scale_req_0 : boolean;
  signal array_obj_ref_1736_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_1736_index_0_scale_req_1 : boolean;
  signal array_obj_ref_1736_index_0_scale_ack_1 : boolean;
  signal ptr_deref_2042_load_3_req_0 : boolean;
  signal ptr_deref_2046_addr_2_ack_0 : boolean;
  signal ptr_deref_2042_load_1_req_0 : boolean;
  signal array_obj_ref_1736_index_sum_1_req_0 : boolean;
  signal array_obj_ref_1736_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_1736_index_sum_1_req_1 : boolean;
  signal ptr_deref_2042_load_1_ack_0 : boolean;
  signal array_obj_ref_1736_index_sum_1_ack_1 : boolean;
  signal ptr_deref_2042_load_3_req_1 : boolean;
  signal array_obj_ref_1736_offset_inst_req_0 : boolean;
  signal array_obj_ref_1736_offset_inst_ack_0 : boolean;
  signal ptr_deref_2046_load_0_ack_0 : boolean;
  signal array_obj_ref_1736_root_address_inst_req_0 : boolean;
  signal ptr_deref_2042_load_3_ack_1 : boolean;
  signal array_obj_ref_1736_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2046_gather_scatter_req_0 : boolean;
  signal ptr_deref_2046_gather_scatter_ack_0 : boolean;
  signal addr_of_1737_final_reg_req_0 : boolean;
  signal ptr_deref_2042_gather_scatter_req_0 : boolean;
  signal addr_of_1737_final_reg_ack_0 : boolean;
  signal ptr_deref_2046_addr_3_ack_0 : boolean;
  signal ptr_deref_2046_addr_2_req_0 : boolean;
  signal ptr_deref_2046_addr_0_req_0 : boolean;
  signal ptr_deref_2042_load_2_req_0 : boolean;
  signal ptr_deref_2042_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2046_addr_0_ack_0 : boolean;
  signal ptr_deref_2042_load_2_ack_0 : boolean;
  signal ptr_deref_2046_addr_0_req_1 : boolean;
  signal ptr_deref_2042_load_0_req_1 : boolean;
  signal ptr_deref_2046_addr_0_ack_1 : boolean;
  signal ptr_deref_2046_addr_3_req_1 : boolean;
  signal ptr_deref_2042_load_0_ack_1 : boolean;
  signal ptr_deref_1741_base_resize_req_0 : boolean;
  signal ptr_deref_1741_base_resize_ack_0 : boolean;
  signal ptr_deref_2046_addr_1_req_0 : boolean;
  signal ptr_deref_1741_root_address_inst_req_0 : boolean;
  signal ptr_deref_1741_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2046_addr_3_req_0 : boolean;
  signal ptr_deref_1741_addr_0_req_0 : boolean;
  signal ptr_deref_1741_addr_0_ack_0 : boolean;
  signal ptr_deref_2046_load_3_req_1 : boolean;
  signal ptr_deref_2046_load_3_ack_1 : boolean;
  signal ptr_deref_2046_addr_1_ack_0 : boolean;
  signal ptr_deref_1741_load_0_req_0 : boolean;
  signal ptr_deref_1741_load_0_ack_0 : boolean;
  signal ptr_deref_2046_addr_1_req_1 : boolean;
  signal ptr_deref_2046_addr_1_ack_1 : boolean;
  signal ptr_deref_1741_load_0_req_1 : boolean;
  signal ptr_deref_1741_load_0_ack_1 : boolean;
  signal ptr_deref_1741_gather_scatter_req_0 : boolean;
  signal ptr_deref_1741_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1745_base_resize_req_0 : boolean;
  signal ptr_deref_1745_base_resize_ack_0 : boolean;
  signal ptr_deref_1745_root_address_inst_req_0 : boolean;
  signal ptr_deref_1745_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1745_addr_0_req_0 : boolean;
  signal ptr_deref_1745_addr_0_ack_0 : boolean;
  signal ptr_deref_1745_load_0_req_0 : boolean;
  signal ptr_deref_1745_load_0_ack_0 : boolean;
  signal ptr_deref_1745_load_0_req_1 : boolean;
  signal ptr_deref_1745_load_0_ack_1 : boolean;
  signal ptr_deref_1745_gather_scatter_req_0 : boolean;
  signal ptr_deref_1745_gather_scatter_ack_0 : boolean;
  signal binary_1750_inst_req_0 : boolean;
  signal binary_1750_inst_ack_0 : boolean;
  signal binary_1750_inst_req_1 : boolean;
  signal binary_1750_inst_ack_1 : boolean;
  signal type_cast_1848_inst_req_0 : boolean;
  signal array_obj_ref_1947_base_resize_req_0 : boolean;
  signal array_obj_ref_1947_base_resize_ack_0 : boolean;
  signal array_obj_ref_1947_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1947_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1947_root_address_inst_req_1 : boolean;
  signal array_obj_ref_1947_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1947_final_reg_req_0 : boolean;
  signal array_obj_ref_1947_final_reg_ack_0 : boolean;
  signal type_cast_1951_inst_req_0 : boolean;
  signal type_cast_1951_inst_ack_0 : boolean;
  signal ptr_deref_1954_base_resize_req_0 : boolean;
  signal ptr_deref_1954_base_resize_ack_0 : boolean;
  signal type_cast_1898_inst_req_0 : boolean;
  signal ptr_deref_1954_root_address_inst_req_0 : boolean;
  signal ptr_deref_1954_root_address_inst_ack_0 : boolean;
  signal phi_stmt_1852_req_1 : boolean;
  signal ptr_deref_1954_addr_0_req_0 : boolean;
  signal type_cast_1898_inst_ack_0 : boolean;
  signal ptr_deref_1954_addr_0_ack_0 : boolean;
  signal ptr_deref_1954_addr_0_req_1 : boolean;
  signal phi_stmt_1893_req_1 : boolean;
  signal ptr_deref_1954_addr_0_ack_1 : boolean;
  signal ptr_deref_1954_addr_1_req_0 : boolean;
  signal ptr_deref_1954_addr_1_ack_0 : boolean;
  signal ptr_deref_1954_addr_1_req_1 : boolean;
  signal ptr_deref_1954_addr_1_ack_1 : boolean;
  signal ptr_deref_1954_addr_2_req_0 : boolean;
  signal ptr_deref_1954_addr_2_ack_0 : boolean;
  signal ptr_deref_1954_addr_2_req_1 : boolean;
  signal ptr_deref_1954_addr_2_ack_1 : boolean;
  signal ptr_deref_1954_addr_3_req_0 : boolean;
  signal ptr_deref_1954_addr_3_ack_0 : boolean;
  signal ptr_deref_1954_addr_3_req_1 : boolean;
  signal ptr_deref_1954_addr_3_ack_1 : boolean;
  signal ptr_deref_1954_gather_scatter_req_0 : boolean;
  signal ptr_deref_1954_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1954_store_0_req_0 : boolean;
  signal ptr_deref_1954_store_0_ack_0 : boolean;
  signal ptr_deref_1954_store_1_req_0 : boolean;
  signal ptr_deref_1954_store_1_ack_0 : boolean;
  signal ptr_deref_1954_store_2_req_0 : boolean;
  signal ptr_deref_1954_store_2_ack_0 : boolean;
  signal ptr_deref_1954_store_3_req_0 : boolean;
  signal ptr_deref_1954_store_3_ack_0 : boolean;
  signal ptr_deref_1954_store_0_req_1 : boolean;
  signal ptr_deref_1954_store_0_ack_1 : boolean;
  signal ptr_deref_1954_store_1_req_1 : boolean;
  signal ptr_deref_1954_store_1_ack_1 : boolean;
  signal ptr_deref_1954_store_2_req_1 : boolean;
  signal ptr_deref_1954_store_2_ack_1 : boolean;
  signal ptr_deref_1954_store_3_req_1 : boolean;
  signal ptr_deref_1954_store_3_ack_1 : boolean;
  signal type_cast_1848_inst_ack_0 : boolean;
  signal array_obj_ref_1961_base_resize_req_0 : boolean;
  signal array_obj_ref_1961_base_resize_ack_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_req_1 : boolean;
  signal phi_stmt_1845_req_0 : boolean;
  signal array_obj_ref_1961_root_address_inst_ack_1 : boolean;
  signal type_cast_1896_inst_req_0 : boolean;
  signal array_obj_ref_1961_final_reg_req_0 : boolean;
  signal array_obj_ref_1961_final_reg_ack_0 : boolean;
  signal type_cast_1896_inst_ack_0 : boolean;
  signal type_cast_1965_inst_req_0 : boolean;
  signal type_cast_1965_inst_ack_0 : boolean;
  signal type_cast_1969_inst_req_0 : boolean;
  signal type_cast_1969_inst_ack_0 : boolean;
  signal ptr_deref_1972_base_resize_req_0 : boolean;
  signal ptr_deref_1972_base_resize_ack_0 : boolean;
  signal phi_stmt_1893_req_0 : boolean;
  signal ptr_deref_1972_root_address_inst_req_0 : boolean;
  signal ptr_deref_1972_root_address_inst_ack_0 : boolean;
  signal ptr_deref_1972_addr_0_req_0 : boolean;
  signal ptr_deref_1972_addr_0_ack_0 : boolean;
  signal ptr_deref_1972_addr_0_req_1 : boolean;
  signal ptr_deref_1972_addr_0_ack_1 : boolean;
  signal ptr_deref_1972_addr_1_req_0 : boolean;
  signal ptr_deref_1972_addr_1_ack_0 : boolean;
  signal ptr_deref_1972_addr_1_req_1 : boolean;
  signal ptr_deref_1972_addr_1_ack_1 : boolean;
  signal ptr_deref_1972_addr_2_req_0 : boolean;
  signal ptr_deref_1972_addr_2_ack_0 : boolean;
  signal ptr_deref_1972_addr_2_req_1 : boolean;
  signal ptr_deref_1972_addr_2_ack_1 : boolean;
  signal ptr_deref_1972_addr_3_req_0 : boolean;
  signal ptr_deref_1972_addr_3_ack_0 : boolean;
  signal ptr_deref_1972_addr_3_req_1 : boolean;
  signal type_cast_1855_inst_req_0 : boolean;
  signal ptr_deref_1972_addr_3_ack_1 : boolean;
  signal ptr_deref_1972_gather_scatter_req_0 : boolean;
  signal ptr_deref_1972_gather_scatter_ack_0 : boolean;
  signal ptr_deref_1972_store_0_req_0 : boolean;
  signal ptr_deref_1972_store_0_ack_0 : boolean;
  signal ptr_deref_1972_store_1_req_0 : boolean;
  signal phi_stmt_1893_ack_0 : boolean;
  signal ptr_deref_1972_store_1_ack_0 : boolean;
  signal ptr_deref_1972_store_2_req_0 : boolean;
  signal ptr_deref_1972_store_2_ack_0 : boolean;
  signal ptr_deref_1972_store_3_req_0 : boolean;
  signal ptr_deref_1972_store_3_ack_0 : boolean;
  signal ptr_deref_1972_store_0_req_1 : boolean;
  signal ptr_deref_1972_store_0_ack_1 : boolean;
  signal ptr_deref_1972_store_1_req_1 : boolean;
  signal ptr_deref_1972_store_1_ack_1 : boolean;
  signal ptr_deref_1972_store_2_req_1 : boolean;
  signal ptr_deref_1972_store_2_ack_1 : boolean;
  signal type_cast_1855_inst_ack_0 : boolean;
  signal ptr_deref_1972_store_3_req_1 : boolean;
  signal ptr_deref_1972_store_3_ack_1 : boolean;
  signal phi_stmt_1852_req_0 : boolean;
  signal type_cast_1978_inst_req_0 : boolean;
  signal type_cast_1978_inst_ack_0 : boolean;
  signal array_obj_ref_1987_base_resize_req_0 : boolean;
  signal array_obj_ref_1987_base_resize_ack_0 : boolean;
  signal phi_stmt_1845_ack_0 : boolean;
  signal array_obj_ref_1987_root_address_inst_req_0 : boolean;
  signal array_obj_ref_1987_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_1987_root_address_inst_req_1 : boolean;
  signal phi_stmt_1852_ack_0 : boolean;
  signal array_obj_ref_1987_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_1987_final_reg_req_0 : boolean;
  signal array_obj_ref_1987_final_reg_ack_0 : boolean;
  signal binary_1993_inst_req_0 : boolean;
  signal binary_1993_inst_ack_0 : boolean;
  signal binary_1993_inst_req_1 : boolean;
  signal binary_1993_inst_ack_1 : boolean;
  signal if_stmt_1995_branch_req_0 : boolean;
  signal if_stmt_1995_branch_ack_1 : boolean;
  signal if_stmt_1995_branch_ack_0 : boolean;
  signal ptr_deref_2003_base_resize_req_0 : boolean;
  signal ptr_deref_2003_base_resize_ack_0 : boolean;
  signal ptr_deref_2003_root_address_inst_req_0 : boolean;
  signal ptr_deref_2003_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2003_addr_0_req_0 : boolean;
  signal ptr_deref_2003_addr_0_ack_0 : boolean;
  signal ptr_deref_2003_gather_scatter_req_0 : boolean;
  signal ptr_deref_2003_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2003_store_0_req_0 : boolean;
  signal ptr_deref_2003_store_0_ack_0 : boolean;
  signal ptr_deref_2003_store_0_req_1 : boolean;
  signal ptr_deref_2003_store_0_ack_1 : boolean;
  signal ptr_deref_2011_base_resize_req_0 : boolean;
  signal ptr_deref_2011_base_resize_ack_0 : boolean;
  signal ptr_deref_2011_root_address_inst_req_0 : boolean;
  signal ptr_deref_2011_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2011_addr_0_req_0 : boolean;
  signal ptr_deref_2011_addr_0_ack_0 : boolean;
  signal ptr_deref_2011_addr_0_req_1 : boolean;
  signal ptr_deref_2011_addr_0_ack_1 : boolean;
  signal ptr_deref_2011_addr_1_req_0 : boolean;
  signal ptr_deref_2011_addr_1_ack_0 : boolean;
  signal ptr_deref_2011_addr_1_req_1 : boolean;
  signal ptr_deref_2011_addr_1_ack_1 : boolean;
  signal ptr_deref_2011_addr_2_req_0 : boolean;
  signal ptr_deref_2011_addr_2_ack_0 : boolean;
  signal ptr_deref_2011_addr_2_req_1 : boolean;
  signal ptr_deref_2011_addr_2_ack_1 : boolean;
  signal ptr_deref_2011_addr_3_req_0 : boolean;
  signal ptr_deref_2011_addr_3_ack_0 : boolean;
  signal ptr_deref_2011_addr_3_req_1 : boolean;
  signal ptr_deref_2011_addr_3_ack_1 : boolean;
  signal ptr_deref_2011_load_0_req_0 : boolean;
  signal ptr_deref_2011_load_0_ack_0 : boolean;
  signal ptr_deref_2011_load_1_req_0 : boolean;
  signal ptr_deref_2011_load_1_ack_0 : boolean;
  signal ptr_deref_2011_load_2_req_0 : boolean;
  signal ptr_deref_2011_load_2_ack_0 : boolean;
  signal ptr_deref_2011_load_3_req_0 : boolean;
  signal ptr_deref_2011_load_3_ack_0 : boolean;
  signal ptr_deref_2011_load_0_req_1 : boolean;
  signal ptr_deref_2011_load_0_ack_1 : boolean;
  signal ptr_deref_2011_load_1_req_1 : boolean;
  signal ptr_deref_2011_load_1_ack_1 : boolean;
  signal ptr_deref_2011_load_2_req_1 : boolean;
  signal ptr_deref_2011_load_2_ack_1 : boolean;
  signal ptr_deref_2011_load_3_req_1 : boolean;
  signal ptr_deref_2011_load_3_ack_1 : boolean;
  signal ptr_deref_2011_gather_scatter_req_0 : boolean;
  signal ptr_deref_2011_gather_scatter_ack_0 : boolean;
  signal binary_2017_inst_req_0 : boolean;
  signal binary_2017_inst_ack_0 : boolean;
  signal binary_2017_inst_req_1 : boolean;
  signal binary_2017_inst_ack_1 : boolean;
  signal ptr_deref_2020_base_resize_req_0 : boolean;
  signal ptr_deref_2020_base_resize_ack_0 : boolean;
  signal ptr_deref_2020_root_address_inst_req_0 : boolean;
  signal ptr_deref_2020_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2020_addr_0_req_0 : boolean;
  signal ptr_deref_2020_addr_0_ack_0 : boolean;
  signal ptr_deref_2020_addr_0_req_1 : boolean;
  signal ptr_deref_2020_addr_0_ack_1 : boolean;
  signal ptr_deref_2020_addr_1_req_0 : boolean;
  signal ptr_deref_2020_addr_1_ack_0 : boolean;
  signal ptr_deref_2020_addr_1_req_1 : boolean;
  signal ptr_deref_2020_addr_1_ack_1 : boolean;
  signal ptr_deref_2020_addr_2_req_0 : boolean;
  signal ptr_deref_2020_addr_2_ack_0 : boolean;
  signal ptr_deref_2020_addr_2_req_1 : boolean;
  signal ptr_deref_2020_addr_2_ack_1 : boolean;
  signal ptr_deref_2020_addr_3_req_0 : boolean;
  signal ptr_deref_2020_addr_3_ack_0 : boolean;
  signal ptr_deref_2020_addr_3_req_1 : boolean;
  signal ptr_deref_2020_addr_3_ack_1 : boolean;
  signal ptr_deref_2020_gather_scatter_req_0 : boolean;
  signal ptr_deref_2020_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2020_store_0_req_0 : boolean;
  signal ptr_deref_2020_store_0_ack_0 : boolean;
  signal ptr_deref_2020_store_1_req_0 : boolean;
  signal ptr_deref_2020_store_1_ack_0 : boolean;
  signal ptr_deref_2020_store_2_req_0 : boolean;
  signal ptr_deref_2020_store_2_ack_0 : boolean;
  signal ptr_deref_2020_store_3_req_0 : boolean;
  signal ptr_deref_2020_store_3_ack_0 : boolean;
  signal ptr_deref_2020_store_0_req_1 : boolean;
  signal ptr_deref_2020_store_0_ack_1 : boolean;
  signal ptr_deref_2020_store_1_req_1 : boolean;
  signal ptr_deref_2020_store_1_ack_1 : boolean;
  signal ptr_deref_2020_store_2_req_1 : boolean;
  signal ptr_deref_2020_store_2_ack_1 : boolean;
  signal ptr_deref_2020_store_3_req_1 : boolean;
  signal ptr_deref_2020_store_3_ack_1 : boolean;
  signal ptr_deref_2025_base_resize_req_0 : boolean;
  signal ptr_deref_2025_base_resize_ack_0 : boolean;
  signal ptr_deref_2025_root_address_inst_req_0 : boolean;
  signal ptr_deref_2025_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2025_addr_0_req_0 : boolean;
  signal ptr_deref_2025_addr_0_ack_0 : boolean;
  signal ptr_deref_2025_addr_0_req_1 : boolean;
  signal ptr_deref_2025_addr_0_ack_1 : boolean;
  signal ptr_deref_2025_addr_1_req_0 : boolean;
  signal ptr_deref_2025_addr_1_ack_0 : boolean;
  signal ptr_deref_2025_addr_1_req_1 : boolean;
  signal ptr_deref_2025_addr_1_ack_1 : boolean;
  signal ptr_deref_2025_addr_2_req_0 : boolean;
  signal ptr_deref_2025_addr_2_ack_0 : boolean;
  signal ptr_deref_2025_addr_2_req_1 : boolean;
  signal ptr_deref_2025_addr_2_ack_1 : boolean;
  signal ptr_deref_2025_addr_3_req_0 : boolean;
  signal ptr_deref_2025_addr_3_ack_0 : boolean;
  signal ptr_deref_2025_addr_3_req_1 : boolean;
  signal ptr_deref_2025_addr_3_ack_1 : boolean;
  signal ptr_deref_2025_load_0_req_0 : boolean;
  signal ptr_deref_2025_load_0_ack_0 : boolean;
  signal ptr_deref_2025_load_1_req_0 : boolean;
  signal ptr_deref_2025_load_1_ack_0 : boolean;
  signal ptr_deref_2025_load_2_req_0 : boolean;
  signal ptr_deref_2025_load_2_ack_0 : boolean;
  signal ptr_deref_2025_load_3_req_0 : boolean;
  signal ptr_deref_2025_load_3_ack_0 : boolean;
  signal ptr_deref_2025_load_0_req_1 : boolean;
  signal ptr_deref_2025_load_0_ack_1 : boolean;
  signal ptr_deref_2025_load_1_req_1 : boolean;
  signal ptr_deref_2025_load_1_ack_1 : boolean;
  signal ptr_deref_2025_load_2_req_1 : boolean;
  signal ptr_deref_2025_load_2_ack_1 : boolean;
  signal ptr_deref_2025_load_3_req_1 : boolean;
  signal ptr_deref_2025_load_3_ack_1 : boolean;
  signal ptr_deref_2025_gather_scatter_req_0 : boolean;
  signal ptr_deref_2025_gather_scatter_ack_0 : boolean;
  signal binary_2031_inst_req_0 : boolean;
  signal binary_2031_inst_ack_0 : boolean;
  signal binary_2031_inst_req_1 : boolean;
  signal binary_2031_inst_ack_1 : boolean;
  signal if_stmt_2033_branch_req_0 : boolean;
  signal if_stmt_2033_branch_ack_1 : boolean;
  signal if_stmt_2033_branch_ack_0 : boolean;
  signal ptr_deref_2042_base_resize_req_0 : boolean;
  signal ptr_deref_2042_base_resize_ack_0 : boolean;
  signal ptr_deref_2042_root_address_inst_req_0 : boolean;
  signal ptr_deref_2042_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2042_addr_0_req_0 : boolean;
  signal ptr_deref_2042_addr_0_ack_0 : boolean;
  signal ptr_deref_2042_addr_0_req_1 : boolean;
  signal ptr_deref_2042_addr_0_ack_1 : boolean;
  signal ptr_deref_2042_addr_1_req_0 : boolean;
  signal ptr_deref_2042_addr_1_ack_0 : boolean;
  signal ptr_deref_2042_addr_1_req_1 : boolean;
  signal ptr_deref_2042_addr_1_ack_1 : boolean;
  signal ptr_deref_2042_addr_2_req_0 : boolean;
  signal ptr_deref_2042_addr_2_ack_0 : boolean;
  signal ptr_deref_2042_addr_2_req_1 : boolean;
  signal ptr_deref_2042_addr_2_ack_1 : boolean;
  signal ptr_deref_2042_addr_3_req_0 : boolean;
  signal ptr_deref_2042_addr_3_ack_0 : boolean;
  signal ptr_deref_2042_addr_3_req_1 : boolean;
  signal ptr_deref_2042_addr_3_ack_1 : boolean;
  signal binary_2051_inst_req_0 : boolean;
  signal binary_2051_inst_ack_0 : boolean;
  signal binary_2051_inst_req_1 : boolean;
  signal binary_2051_inst_ack_1 : boolean;
  signal if_stmt_2053_branch_req_0 : boolean;
  signal if_stmt_2053_branch_ack_1 : boolean;
  signal if_stmt_2053_branch_ack_0 : boolean;
  signal ptr_deref_2062_base_resize_req_0 : boolean;
  signal ptr_deref_2062_base_resize_ack_0 : boolean;
  signal ptr_deref_2062_root_address_inst_req_0 : boolean;
  signal ptr_deref_2062_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2062_addr_0_req_0 : boolean;
  signal ptr_deref_2062_addr_0_ack_0 : boolean;
  signal ptr_deref_2062_addr_0_req_1 : boolean;
  signal ptr_deref_2062_addr_0_ack_1 : boolean;
  signal ptr_deref_2062_addr_1_req_0 : boolean;
  signal ptr_deref_2062_addr_1_ack_0 : boolean;
  signal ptr_deref_2062_addr_1_req_1 : boolean;
  signal ptr_deref_2062_addr_1_ack_1 : boolean;
  signal ptr_deref_2062_addr_2_req_0 : boolean;
  signal ptr_deref_2062_addr_2_ack_0 : boolean;
  signal ptr_deref_2062_addr_2_req_1 : boolean;
  signal ptr_deref_2062_addr_2_ack_1 : boolean;
  signal ptr_deref_2062_addr_3_req_0 : boolean;
  signal ptr_deref_2062_addr_3_ack_0 : boolean;
  signal ptr_deref_2062_addr_3_req_1 : boolean;
  signal ptr_deref_2062_addr_3_ack_1 : boolean;
  signal ptr_deref_2062_load_0_req_0 : boolean;
  signal ptr_deref_2062_load_0_ack_0 : boolean;
  signal ptr_deref_2062_load_1_req_0 : boolean;
  signal ptr_deref_2062_load_1_ack_0 : boolean;
  signal ptr_deref_2062_load_2_req_0 : boolean;
  signal ptr_deref_2062_load_2_ack_0 : boolean;
  signal ptr_deref_2062_load_3_req_0 : boolean;
  signal ptr_deref_2062_load_3_ack_0 : boolean;
  signal ptr_deref_2062_load_0_req_1 : boolean;
  signal ptr_deref_2062_load_0_ack_1 : boolean;
  signal ptr_deref_2062_load_1_req_1 : boolean;
  signal ptr_deref_2062_load_1_ack_1 : boolean;
  signal ptr_deref_2062_load_2_req_1 : boolean;
  signal ptr_deref_2062_load_2_ack_1 : boolean;
  signal ptr_deref_2062_load_3_req_1 : boolean;
  signal ptr_deref_2062_load_3_ack_1 : boolean;
  signal ptr_deref_2062_gather_scatter_req_0 : boolean;
  signal ptr_deref_2062_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2067_base_resize_req_0 : boolean;
  signal ptr_deref_2067_base_resize_ack_0 : boolean;
  signal ptr_deref_2067_root_address_inst_req_0 : boolean;
  signal ptr_deref_2067_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2067_addr_0_req_0 : boolean;
  signal ptr_deref_2067_addr_0_ack_0 : boolean;
  signal ptr_deref_2067_gather_scatter_req_0 : boolean;
  signal ptr_deref_2067_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2067_store_0_req_0 : boolean;
  signal ptr_deref_2067_store_0_ack_0 : boolean;
  signal ptr_deref_2067_store_0_req_1 : boolean;
  signal ptr_deref_2067_store_0_ack_1 : boolean;
  signal binary_2077_inst_req_0 : boolean;
  signal binary_2077_inst_ack_0 : boolean;
  signal binary_2077_inst_req_1 : boolean;
  signal binary_2077_inst_ack_1 : boolean;
  signal simple_obj_ref_2074_inst_req_0 : boolean;
  signal simple_obj_ref_2074_inst_ack_0 : boolean;
  signal array_obj_ref_2086_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2086_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2086_index_0_scale_req_0 : boolean;
  signal array_obj_ref_2086_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_2086_index_0_scale_req_1 : boolean;
  signal array_obj_ref_2086_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_2086_index_sum_1_req_0 : boolean;
  signal array_obj_ref_2086_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_2086_index_sum_1_req_1 : boolean;
  signal array_obj_ref_2086_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_2086_offset_inst_req_0 : boolean;
  signal array_obj_ref_2086_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2086_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2086_root_address_inst_ack_0 : boolean;
  signal addr_of_2087_final_reg_req_0 : boolean;
  signal addr_of_2087_final_reg_ack_0 : boolean;
  signal ptr_deref_2091_base_resize_req_0 : boolean;
  signal ptr_deref_2091_base_resize_ack_0 : boolean;
  signal ptr_deref_2091_root_address_inst_req_0 : boolean;
  signal ptr_deref_2091_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2091_addr_0_req_0 : boolean;
  signal ptr_deref_2091_addr_0_ack_0 : boolean;
  signal ptr_deref_2091_load_0_req_0 : boolean;
  signal ptr_deref_2091_load_0_ack_0 : boolean;
  signal ptr_deref_2091_load_0_req_1 : boolean;
  signal ptr_deref_2091_load_0_ack_1 : boolean;
  signal ptr_deref_2091_gather_scatter_req_0 : boolean;
  signal ptr_deref_2091_gather_scatter_ack_0 : boolean;
  signal binary_2097_inst_req_0 : boolean;
  signal binary_2097_inst_ack_0 : boolean;
  signal binary_2097_inst_req_1 : boolean;
  signal binary_2097_inst_ack_1 : boolean;
  signal array_obj_ref_2105_index_2_resize_req_0 : boolean;
  signal array_obj_ref_2105_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_2105_index_2_rename_req_0 : boolean;
  signal array_obj_ref_2105_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_2105_index_sum_1_req_0 : boolean;
  signal array_obj_ref_2105_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_2105_index_sum_1_req_1 : boolean;
  signal array_obj_ref_2105_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_2105_offset_inst_req_0 : boolean;
  signal array_obj_ref_2105_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2105_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2105_root_address_inst_ack_0 : boolean;
  signal addr_of_2106_final_reg_req_0 : boolean;
  signal addr_of_2106_final_reg_ack_0 : boolean;
  signal ptr_deref_2110_base_resize_req_0 : boolean;
  signal ptr_deref_2110_base_resize_ack_0 : boolean;
  signal ptr_deref_2110_root_address_inst_req_0 : boolean;
  signal ptr_deref_2110_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2110_addr_0_req_0 : boolean;
  signal ptr_deref_2110_addr_0_ack_0 : boolean;
  signal ptr_deref_2110_load_0_req_0 : boolean;
  signal ptr_deref_2110_load_0_ack_0 : boolean;
  signal ptr_deref_2110_load_0_req_1 : boolean;
  signal ptr_deref_2110_load_0_ack_1 : boolean;
  signal ptr_deref_2110_gather_scatter_req_0 : boolean;
  signal ptr_deref_2110_gather_scatter_ack_0 : boolean;
  signal binary_2116_inst_req_0 : boolean;
  signal binary_2116_inst_ack_0 : boolean;
  signal binary_2116_inst_req_1 : boolean;
  signal binary_2116_inst_ack_1 : boolean;
  signal if_stmt_2118_branch_req_0 : boolean;
  signal if_stmt_2118_branch_ack_1 : boolean;
  signal if_stmt_2118_branch_ack_0 : boolean;
  signal binary_2129_inst_req_0 : boolean;
  signal binary_2129_inst_ack_0 : boolean;
  signal binary_2129_inst_req_1 : boolean;
  signal binary_2129_inst_ack_1 : boolean;
  signal array_obj_ref_2137_index_2_resize_req_0 : boolean;
  signal array_obj_ref_2137_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_2137_index_2_rename_req_0 : boolean;
  signal array_obj_ref_2137_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_2137_index_sum_1_req_0 : boolean;
  signal array_obj_ref_2137_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_2137_index_sum_1_req_1 : boolean;
  signal array_obj_ref_2137_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_2137_offset_inst_req_0 : boolean;
  signal array_obj_ref_2137_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2137_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2137_root_address_inst_ack_0 : boolean;
  signal addr_of_2138_final_reg_req_0 : boolean;
  signal addr_of_2138_final_reg_ack_0 : boolean;
  signal ptr_deref_2142_base_resize_req_0 : boolean;
  signal ptr_deref_2142_base_resize_ack_0 : boolean;
  signal ptr_deref_2142_root_address_inst_req_0 : boolean;
  signal ptr_deref_2142_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2142_addr_0_req_0 : boolean;
  signal ptr_deref_2142_addr_0_ack_0 : boolean;
  signal ptr_deref_2142_load_0_req_0 : boolean;
  signal ptr_deref_2142_load_0_ack_0 : boolean;
  signal ptr_deref_2142_load_0_req_1 : boolean;
  signal ptr_deref_2142_load_0_ack_1 : boolean;
  signal ptr_deref_2142_gather_scatter_req_0 : boolean;
  signal ptr_deref_2142_gather_scatter_ack_0 : boolean;
  signal binary_2148_inst_req_0 : boolean;
  signal binary_2148_inst_ack_0 : boolean;
  signal binary_2148_inst_req_1 : boolean;
  signal binary_2148_inst_ack_1 : boolean;
  signal if_stmt_2150_branch_req_0 : boolean;
  signal if_stmt_2150_branch_ack_1 : boolean;
  signal if_stmt_2150_branch_ack_0 : boolean;
  signal binary_2161_inst_req_0 : boolean;
  signal binary_2161_inst_ack_0 : boolean;
  signal binary_2161_inst_req_1 : boolean;
  signal binary_2161_inst_ack_1 : boolean;
  signal array_obj_ref_2169_index_2_resize_req_0 : boolean;
  signal array_obj_ref_2169_index_2_resize_ack_0 : boolean;
  signal array_obj_ref_2169_index_2_rename_req_0 : boolean;
  signal array_obj_ref_2169_index_2_rename_ack_0 : boolean;
  signal array_obj_ref_2169_index_sum_1_req_0 : boolean;
  signal array_obj_ref_2169_index_sum_1_ack_0 : boolean;
  signal array_obj_ref_2169_index_sum_1_req_1 : boolean;
  signal array_obj_ref_2169_index_sum_1_ack_1 : boolean;
  signal array_obj_ref_2169_offset_inst_req_0 : boolean;
  signal array_obj_ref_2169_offset_inst_ack_0 : boolean;
  signal array_obj_ref_2169_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2169_root_address_inst_ack_0 : boolean;
  signal addr_of_2170_final_reg_req_0 : boolean;
  signal addr_of_2170_final_reg_ack_0 : boolean;
  signal ptr_deref_2174_base_resize_req_0 : boolean;
  signal ptr_deref_2174_base_resize_ack_0 : boolean;
  signal ptr_deref_2174_root_address_inst_req_0 : boolean;
  signal ptr_deref_2174_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2174_addr_0_req_0 : boolean;
  signal ptr_deref_2174_addr_0_ack_0 : boolean;
  signal ptr_deref_2174_load_0_req_0 : boolean;
  signal ptr_deref_2174_load_0_ack_0 : boolean;
  signal ptr_deref_2174_load_0_req_1 : boolean;
  signal ptr_deref_2174_load_0_ack_1 : boolean;
  signal ptr_deref_2174_gather_scatter_req_0 : boolean;
  signal ptr_deref_2174_gather_scatter_ack_0 : boolean;
  signal type_cast_2179_inst_req_0 : boolean;
  signal type_cast_2179_inst_ack_0 : boolean;
  signal binary_2183_inst_req_0 : boolean;
  signal binary_2183_inst_ack_0 : boolean;
  signal binary_2183_inst_req_1 : boolean;
  signal binary_2183_inst_ack_1 : boolean;
  signal if_stmt_2185_branch_req_0 : boolean;
  signal if_stmt_2185_branch_ack_1 : boolean;
  signal if_stmt_2185_branch_ack_0 : boolean;
  signal type_cast_2194_inst_req_0 : boolean;
  signal type_cast_2194_inst_ack_0 : boolean;
  signal binary_2198_inst_req_0 : boolean;
  signal binary_2198_inst_ack_0 : boolean;
  signal binary_2198_inst_req_1 : boolean;
  signal binary_2198_inst_ack_1 : boolean;
  signal if_stmt_2200_branch_req_0 : boolean;
  signal if_stmt_2200_branch_ack_1 : boolean;
  signal if_stmt_2200_branch_ack_0 : boolean;
  signal binary_2211_inst_req_0 : boolean;
  signal binary_2211_inst_ack_0 : boolean;
  signal binary_2211_inst_req_1 : boolean;
  signal binary_2211_inst_ack_1 : boolean;
  signal if_stmt_2213_branch_req_0 : boolean;
  signal if_stmt_2213_branch_ack_1 : boolean;
  signal if_stmt_2213_branch_ack_0 : boolean;
  signal binary_2224_inst_req_0 : boolean;
  signal binary_2224_inst_ack_0 : boolean;
  signal binary_2224_inst_req_1 : boolean;
  signal binary_2224_inst_ack_1 : boolean;
  signal if_stmt_2226_branch_req_0 : boolean;
  signal if_stmt_2226_branch_ack_1 : boolean;
  signal if_stmt_2226_branch_ack_0 : boolean;
  signal type_cast_2235_inst_req_0 : boolean;
  signal type_cast_2235_inst_ack_0 : boolean;
  signal binary_2239_inst_req_0 : boolean;
  signal binary_2239_inst_ack_0 : boolean;
  signal binary_2239_inst_req_1 : boolean;
  signal binary_2239_inst_ack_1 : boolean;
  signal if_stmt_2241_branch_req_0 : boolean;
  signal if_stmt_2241_branch_ack_1 : boolean;
  signal if_stmt_2241_branch_ack_0 : boolean;
  signal binary_2252_inst_req_0 : boolean;
  signal binary_2252_inst_ack_0 : boolean;
  signal binary_2252_inst_req_1 : boolean;
  signal binary_2252_inst_ack_1 : boolean;
  signal if_stmt_2254_branch_req_0 : boolean;
  signal if_stmt_2254_branch_ack_1 : boolean;
  signal if_stmt_2254_branch_ack_0 : boolean;
  signal binary_2265_inst_req_0 : boolean;
  signal binary_2265_inst_ack_0 : boolean;
  signal binary_2265_inst_req_1 : boolean;
  signal binary_2265_inst_ack_1 : boolean;
  signal if_stmt_2267_branch_req_0 : boolean;
  signal if_stmt_2267_branch_ack_1 : boolean;
  signal if_stmt_2267_branch_ack_0 : boolean;
  signal type_cast_2276_inst_req_0 : boolean;
  signal type_cast_2276_inst_ack_0 : boolean;
  signal simple_obj_ref_2274_inst_req_0 : boolean;
  signal simple_obj_ref_2274_inst_ack_0 : boolean;
  signal type_cast_2282_inst_req_0 : boolean;
  signal type_cast_2282_inst_ack_0 : boolean;
  signal simple_obj_ref_2280_inst_req_0 : boolean;
  signal simple_obj_ref_2280_inst_ack_0 : boolean;
  signal type_cast_2288_inst_req_0 : boolean;
  signal type_cast_2288_inst_ack_0 : boolean;
  signal simple_obj_ref_2286_inst_req_0 : boolean;
  signal simple_obj_ref_2286_inst_ack_0 : boolean;
  signal type_cast_2294_inst_req_0 : boolean;
  signal type_cast_2294_inst_ack_0 : boolean;
  signal simple_obj_ref_2292_inst_req_0 : boolean;
  signal simple_obj_ref_2292_inst_ack_0 : boolean;
  signal type_cast_2300_inst_req_0 : boolean;
  signal type_cast_2300_inst_ack_0 : boolean;
  signal simple_obj_ref_2298_inst_req_0 : boolean;
  signal simple_obj_ref_2298_inst_ack_0 : boolean;
  signal phi_stmt_1778_req_1 : boolean;
  signal type_cast_1781_inst_req_0 : boolean;
  signal type_cast_1781_inst_ack_0 : boolean;
  signal phi_stmt_1778_req_0 : boolean;
  signal phi_stmt_1778_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_rtt_CP_7287: Block -- control-path 
    signal cp_elements: BooleanArray(1031 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1031);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(1031), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(134) & cp_elements(953));
    cp_elements(2) <= OrReduce(cp_elements(132) & cp_elements(959));
    cp_elements(3) <= OrReduce(cp_elements(961) & cp_elements(963));
    cp_elements(4) <= cp_elements(200);
    cp_elements(5) <= OrReduce(cp_elements(207) & cp_elements(965));
    cp_elements(6) <= cp_elements(980);
    cp_elements(7) <= OrReduce(cp_elements(238) & cp_elements(982));
    cp_elements(8) <= OrReduce(cp_elements(269) & cp_elements(995));
    cp_elements(9) <= OrReduce(cp_elements(284) & cp_elements(997));
    cp_elements(10) <= cp_elements(420);
    cp_elements(11) <= OrReduce(cp_elements(429) & cp_elements(999));
    cp_elements(12) <= cp_elements(560);
    cp_elements(13) <= OrReduce(cp_elements(567) & cp_elements(1003));
    cp_elements(14) <= OrReduce(cp_elements(651) & cp_elements(1005));
    base_resize_req_9436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => ptr_deref_2062_base_resize_req_0); -- 
    cp_elements(15) <= OrReduce(cp_elements(752) & cp_elements(1011));
    cp_elements(16) <= OrReduce(cp_elements(786) & cp_elements(1013));
    cp_elements(17) <= OrReduce(cp_elements(825) & cp_elements(1015));
    cp_elements(18) <= OrReduce(cp_elements(843) & cp_elements(1017));
    cp_elements(19) <= OrReduce(cp_elements(841) & cp_elements(1019));
    cp_elements(20) <= OrReduce(cp_elements(823) & cp_elements(1021));
    cp_elements(21) <= OrReduce(cp_elements(891) & cp_elements(1023));
    cp_elements(22) <= OrReduce(cp_elements(889) & cp_elements(1025));
    cp_elements(23) <= OrReduce(cp_elements(919) & cp_elements(1027));
    cp_elements(24) <= cp_elements(0);
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(26) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => type_cast_1698_inst_req_0); -- 
    cp_elements(26) <= cp_elements(24);
    cp_elements(27) <= cp_elements(24);
    req_7476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => simple_obj_ref_1697_inst_req_0); -- 
    ack_7477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1697_inst_ack_0, ack => cp_elements(28)); -- 
    ack_7482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1698_inst_ack_0, ack => cp_elements(29)); -- 
    cp_elements(30) <= cp_elements(29);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(33));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7494_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => type_cast_1702_inst_req_0); -- 
    cp_elements(32) <= cp_elements(30);
    cp_elements(33) <= cp_elements(30);
    ack_7495_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1702_inst_ack_0, ack => cp_elements(34)); -- 
    base_resize_req_7506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => array_obj_ref_1709_base_resize_req_0); -- 
    cp_elements(35) <= cp_elements(30);
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_1709_final_reg_req_0); -- 
    base_resize_ack_7507_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1709_base_resize_ack_0, ack => cp_elements(37)); -- 
    plus_base_rr_7512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_1709_root_address_inst_req_0); -- 
    plus_base_ra_7513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1709_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    plus_base_cr_7514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_1709_root_address_inst_req_1); -- 
    plus_base_ca_7515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1709_root_address_inst_ack_1, ack => cp_elements(39)); -- 
    final_reg_ack_7520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1709_final_reg_ack_0, ack => cp_elements(40)); -- 
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(40) & cp_elements(42));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => type_cast_1713_inst_req_0); -- 
    cp_elements(42) <= cp_elements(30);
    ack_7530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1713_inst_ack_0, ack => cp_elements(43)); -- 
    base_resize_req_7543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_1717_base_resize_req_0); -- 
    base_resize_ack_7544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_base_resize_ack_0, ack => cp_elements(44)); -- 
    sum_rename_req_7548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_1717_root_address_inst_req_0); -- 
    cp_elements(45) <= ptr_deref_1717_root_address_inst_ack_0;
    cp_elements(46) <= cp_elements(45);
    rr_7556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => ptr_deref_1717_addr_0_req_0); -- 
    ra_7557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_0_ack_0, ack => cp_elements(47)); -- 
    cr_7558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_1717_addr_0_req_1); -- 
    ca_7559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(45);
    rr_7563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_1717_addr_1_req_0); -- 
    ra_7564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_1_ack_0, ack => cp_elements(50)); -- 
    cr_7565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => ptr_deref_1717_addr_1_req_1); -- 
    ca_7566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_1_ack_1, ack => cp_elements(51)); -- 
    cp_elements(52) <= cp_elements(45);
    rr_7570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => ptr_deref_1717_addr_2_req_0); -- 
    ra_7571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_2_ack_0, ack => cp_elements(53)); -- 
    cr_7572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => ptr_deref_1717_addr_2_req_1); -- 
    ca_7573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_2_ack_1, ack => cp_elements(54)); -- 
    cp_elements(55) <= cp_elements(45);
    rr_7577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_1717_addr_3_req_0); -- 
    ra_7578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_3_ack_0, ack => cp_elements(56)); -- 
    cr_7579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_1717_addr_3_req_1); -- 
    ca_7580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_addr_3_ack_1, ack => cp_elements(57)); -- 
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(51) & cp_elements(54) & cp_elements(57));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(59) <= cp_elements(58);
    rr_7590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_1717_load_0_req_0); -- 
    ra_7591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_0, ack => cp_elements(60)); -- 
    cp_elements(61) <= cp_elements(58);
    rr_7595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_1717_load_1_req_0); -- 
    ra_7596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_1_ack_0, ack => cp_elements(62)); -- 
    cp_elements(63) <= cp_elements(58);
    rr_7600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => ptr_deref_1717_load_2_req_0); -- 
    ra_7601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_2_ack_0, ack => cp_elements(64)); -- 
    cp_elements(65) <= cp_elements(58);
    rr_7605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_1717_load_3_req_0); -- 
    ra_7606_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_3_ack_0, ack => cp_elements(66)); -- 
    cpelement_group_67 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(62) & cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(67),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(68) <= cp_elements(67);
    cr_7616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_1717_load_0_req_1); -- 
    ca_7617_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_0_ack_1, ack => cp_elements(69)); -- 
    cp_elements(70) <= cp_elements(67);
    cr_7621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_1717_load_1_req_1); -- 
    ca_7622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_1_ack_1, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(67);
    cr_7626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_1717_load_2_req_1); -- 
    ca_7627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_2_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= cp_elements(67);
    cr_7631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_1717_load_3_req_1); -- 
    ca_7632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_load_3_ack_1, ack => cp_elements(75)); -- 
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(69) & cp_elements(71) & cp_elements(73) & cp_elements(75));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_7633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_1717_gather_scatter_req_0); -- 
    merge_ack_7634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1717_gather_scatter_ack_0, ack => cp_elements(77)); -- 
    phi_stmt_1778_req_10445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => phi_stmt_1778_req_1); -- 
    cp_elements(78) <= cp_elements(156);
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(80) & cp_elements(88));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => addr_of_1728_final_reg_req_0); -- 
    cp_elements(80) <= cp_elements(78);
    cp_elements(81) <= cp_elements(78);
    index_resize_req_7651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => array_obj_ref_1727_index_0_resize_req_0); -- 
    index_resize_ack_7652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_index_0_resize_ack_0, ack => cp_elements(82)); -- 
    scale_rr_7656_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => array_obj_ref_1727_index_0_scale_req_0); -- 
    scale_ra_7657_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_index_0_scale_ack_0, ack => cp_elements(83)); -- 
    scale_cr_7658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => array_obj_ref_1727_index_0_scale_req_1); -- 
    scale_ca_7659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_index_0_scale_ack_1, ack => cp_elements(84)); -- 
    partial_sum_1_rr_7663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => array_obj_ref_1727_index_sum_1_req_0); -- 
    partial_sum_1_ra_7664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_index_sum_1_ack_0, ack => cp_elements(85)); -- 
    partial_sum_1_cr_7665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => array_obj_ref_1727_index_sum_1_req_1); -- 
    partial_sum_1_ca_7666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_index_sum_1_ack_1, ack => cp_elements(86)); -- 
    final_index_req_7667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => array_obj_ref_1727_offset_inst_req_0); -- 
    final_index_ack_7668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_offset_inst_ack_0, ack => cp_elements(87)); -- 
    sum_rename_req_7672_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => array_obj_ref_1727_root_address_inst_req_0); -- 
    sum_rename_ack_7673_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1727_root_address_inst_ack_0, ack => cp_elements(88)); -- 
    final_reg_ack_7678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1728_final_reg_ack_0, ack => cp_elements(89)); -- 
    base_resize_req_7732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_1741_base_resize_req_0); -- 
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_7718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => addr_of_1737_final_reg_req_0); -- 
    cp_elements(91) <= cp_elements(78);
    cp_elements(92) <= cp_elements(78);
    index_resize_req_7692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => array_obj_ref_1736_index_0_resize_req_0); -- 
    index_resize_ack_7693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_0_resize_ack_0, ack => cp_elements(93)); -- 
    scale_rr_7697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => array_obj_ref_1736_index_0_scale_req_0); -- 
    scale_ra_7698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_0_scale_ack_0, ack => cp_elements(94)); -- 
    scale_cr_7699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => array_obj_ref_1736_index_0_scale_req_1); -- 
    scale_ca_7700_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_0_scale_ack_1, ack => cp_elements(95)); -- 
    partial_sum_1_rr_7704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_1736_index_sum_1_req_0); -- 
    partial_sum_1_ra_7705_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_sum_1_ack_0, ack => cp_elements(96)); -- 
    partial_sum_1_cr_7706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_1736_index_sum_1_req_1); -- 
    partial_sum_1_ca_7707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_index_sum_1_ack_1, ack => cp_elements(97)); -- 
    final_index_req_7708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => array_obj_ref_1736_offset_inst_req_0); -- 
    final_index_ack_7709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_offset_inst_ack_0, ack => cp_elements(98)); -- 
    sum_rename_req_7713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_1736_root_address_inst_req_0); -- 
    sum_rename_ack_7714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1736_root_address_inst_ack_0, ack => cp_elements(99)); -- 
    final_reg_ack_7719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1737_final_reg_ack_0, ack => cp_elements(100)); -- 
    base_resize_req_7780_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_1745_base_resize_req_0); -- 
    base_resize_ack_7733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_base_resize_ack_0, ack => cp_elements(101)); -- 
    sum_rename_req_7737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_1741_root_address_inst_req_0); -- 
    sum_rename_ack_7738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_root_address_inst_ack_0, ack => cp_elements(102)); -- 
    root_rename_req_7742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => ptr_deref_1741_addr_0_req_0); -- 
    root_rename_ack_7743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_addr_0_ack_0, ack => cp_elements(103)); -- 
    rr_7753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_1741_load_0_req_0); -- 
    ra_7754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_load_0_ack_0, ack => cp_elements(104)); -- 
    cr_7764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => ptr_deref_1741_load_0_req_1); -- 
    ca_7765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_load_0_ack_1, ack => cp_elements(105)); -- 
    merge_req_7766_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_1741_gather_scatter_req_0); -- 
    merge_ack_7767_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1741_gather_scatter_ack_0, ack => cp_elements(106)); -- 
    base_resize_ack_7781_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_base_resize_ack_0, ack => cp_elements(107)); -- 
    sum_rename_req_7785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_1745_root_address_inst_req_0); -- 
    sum_rename_ack_7786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_root_address_inst_ack_0, ack => cp_elements(108)); -- 
    root_rename_req_7790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => ptr_deref_1745_addr_0_req_0); -- 
    root_rename_ack_7791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_addr_0_ack_0, ack => cp_elements(109)); -- 
    rr_7801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_1745_load_0_req_0); -- 
    ra_7802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_load_0_ack_0, ack => cp_elements(110)); -- 
    cr_7812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_1745_load_0_req_1); -- 
    ca_7813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_load_0_ack_1, ack => cp_elements(111)); -- 
    merge_req_7814_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_1745_gather_scatter_req_0); -- 
    merge_ack_7815_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1745_gather_scatter_ack_0, ack => cp_elements(112)); -- 
    cpelement_group_113 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(106) & cp_elements(114) & cp_elements(115));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(113),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7825_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => binary_1750_inst_req_0); -- 
    cp_elements(114) <= cp_elements(78);
    cp_elements(115) <= cp_elements(78);
    ra_7826_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1750_inst_ack_0, ack => cp_elements(116)); -- 
    cr_7827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => binary_1750_inst_req_1); -- 
    ca_7828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1750_inst_ack_1, ack => cp_elements(117)); -- 
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(112) & cp_elements(117) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => binary_1755_inst_req_0); -- 
    cp_elements(119) <= cp_elements(78);
    ra_7839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1755_inst_ack_0, ack => cp_elements(120)); -- 
    cr_7840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => binary_1755_inst_req_1); -- 
    ca_7841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1755_inst_ack_1, ack => cp_elements(121)); -- 
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(121) & cp_elements(123));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => binary_1761_inst_req_0); -- 
    cp_elements(123) <= cp_elements(78);
    ra_7851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1761_inst_ack_0, ack => cp_elements(124)); -- 
    cr_7852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => binary_1761_inst_req_1); -- 
    ca_7853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1761_inst_ack_1, ack => cp_elements(125)); -- 
    cp_elements(126) <= cp_elements(125);
    cp_elements(127) <= false;
    cp_elements(128) <= cp_elements(127);
    cp_elements(129) <= cp_elements(125);
    branch_req_7861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => if_stmt_1763_branch_req_0); -- 
    cp_elements(130) <= cp_elements(129);
    cp_elements(131) <= cp_elements(130);
    if_choice_transition_7866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1763_branch_ack_1, ack => cp_elements(132)); -- 
    cp_elements(133) <= cp_elements(130);
    else_choice_transition_7870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1763_branch_ack_0, ack => cp_elements(134)); -- 
    cp_elements(135) <= cp_elements(1);
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(138));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => binary_1774_inst_req_0); -- 
    cp_elements(137) <= cp_elements(135);
    cp_elements(138) <= cp_elements(135);
    ra_7885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1774_inst_ack_0, ack => cp_elements(139)); -- 
    cr_7886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => binary_1774_inst_req_1); -- 
    ca_7887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1774_inst_ack_1, ack => cp_elements(140)); -- 
    req_10458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => type_cast_1781_inst_req_0); -- 
    cp_elements(141) <= cp_elements(957);
    cpelement_group_142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(147));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => binary_1792_inst_req_0); -- 
    cp_elements(143) <= cp_elements(141);
    cpelement_group_144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(145) & cp_elements(146));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => type_cast_1788_inst_req_0); -- 
    cp_elements(145) <= cp_elements(141);
    cp_elements(146) <= cp_elements(141);
    ack_7902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1788_inst_ack_0, ack => cp_elements(147)); -- 
    ra_7907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1792_inst_ack_0, ack => cp_elements(148)); -- 
    cr_7908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => binary_1792_inst_req_1); -- 
    ca_7909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1792_inst_ack_1, ack => cp_elements(149)); -- 
    cp_elements(150) <= cp_elements(149);
    cp_elements(151) <= false;
    cp_elements(152) <= cp_elements(151);
    cp_elements(153) <= cp_elements(149);
    branch_req_7917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => if_stmt_1794_branch_req_0); -- 
    cp_elements(154) <= cp_elements(153);
    cp_elements(155) <= cp_elements(154);
    if_choice_transition_7922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1794_branch_ack_1, ack => cp_elements(156)); -- 
    cp_elements(157) <= cp_elements(154);
    else_choice_transition_7926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1794_branch_ack_0, ack => cp_elements(158)); -- 
    cp_elements(159) <= cp_elements(2);
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(161) & cp_elements(165));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_7947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_1807_inst_req_0); -- 
    cp_elements(161) <= cp_elements(159);
    cpelement_group_162 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(163) & cp_elements(164));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(162),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_7942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => type_cast_1803_inst_req_0); -- 
    cp_elements(163) <= cp_elements(159);
    cp_elements(164) <= cp_elements(159);
    ack_7943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1803_inst_ack_0, ack => cp_elements(165)); -- 
    ra_7948_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1807_inst_ack_0, ack => cp_elements(166)); -- 
    cr_7949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => binary_1807_inst_req_1); -- 
    ca_7950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1807_inst_ack_1, ack => cp_elements(167)); -- 
    cp_elements(168) <= cp_elements(167);
    cp_elements(169) <= false;
    cp_elements(170) <= cp_elements(169);
    cp_elements(171) <= cp_elements(167);
    branch_req_7958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => if_stmt_1809_branch_req_0); -- 
    cp_elements(172) <= cp_elements(171);
    cp_elements(173) <= cp_elements(172);
    if_choice_transition_7963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_1, ack => cp_elements(174)); -- 
    cp_elements(175) <= cp_elements(172);
    else_choice_transition_7967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1809_branch_ack_0, ack => cp_elements(176)); -- 
    cp_elements(177) <= cp_elements(3);
    cp_elements(178) <= cp_elements(177);
    rr_7988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => simple_obj_ref_1817_load_0_req_0); -- 
    ra_7989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1817_load_0_ack_0, ack => cp_elements(179)); -- 
    cr_7999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => simple_obj_ref_1817_load_0_req_1); -- 
    ca_8000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1817_load_0_ack_1, ack => cp_elements(180)); -- 
    merge_req_8001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => simple_obj_ref_1817_gather_scatter_req_0); -- 
    merge_ack_8002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1817_gather_scatter_ack_0, ack => cp_elements(181)); -- 
    cpelement_group_182 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(183));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(182),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(182), ack => binary_1823_inst_req_0); -- 
    cp_elements(183) <= cp_elements(177);
    ra_8012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1823_inst_ack_0, ack => cp_elements(184)); -- 
    cr_8013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(184), ack => binary_1823_inst_req_1); -- 
    cp_elements(185) <= binary_1823_inst_ack_1;
    cp_elements(186) <= cp_elements(185);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => simple_obj_ref_1825_gather_scatter_req_0); -- 
    cp_elements(188) <= cp_elements(177);
    split_ack_8026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1825_gather_scatter_ack_0, ack => cp_elements(189)); -- 
    rr_8033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => simple_obj_ref_1825_store_0_req_0); -- 
    ra_8034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1825_store_0_ack_0, ack => cp_elements(190)); -- 
    cr_8044_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => simple_obj_ref_1825_store_0_req_1); -- 
    ca_8045_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_1825_store_0_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(193) & cp_elements(197));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => binary_1834_inst_req_0); -- 
    cp_elements(193) <= cp_elements(177);
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(195) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => type_cast_1830_inst_req_0); -- 
    cp_elements(195) <= cp_elements(177);
    cp_elements(196) <= cp_elements(185);
    ack_8057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1830_inst_ack_0, ack => cp_elements(197)); -- 
    ra_8062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1834_inst_ack_0, ack => cp_elements(198)); -- 
    cr_8063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => binary_1834_inst_req_1); -- 
    ca_8064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1834_inst_ack_1, ack => cp_elements(199)); -- 
    cpelement_group_200 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(199));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(200),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(201) <= cp_elements(4);
    cp_elements(202) <= false;
    cp_elements(203) <= cp_elements(202);
    cp_elements(204) <= cp_elements(4);
    branch_req_8072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => if_stmt_1836_branch_req_0); -- 
    cp_elements(205) <= cp_elements(204);
    cp_elements(206) <= cp_elements(205);
    if_choice_transition_8077_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1836_branch_ack_1, ack => cp_elements(207)); -- 
    cp_elements(208) <= cp_elements(205);
    else_choice_transition_8081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1836_branch_ack_0, ack => cp_elements(209)); -- 
    cp_elements(210) <= cp_elements(6);
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(212) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => addr_of_1865_final_reg_req_0); -- 
    cp_elements(212) <= cp_elements(210);
    cp_elements(213) <= cp_elements(210);
    index_resize_req_8100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => array_obj_ref_1864_index_0_resize_req_0); -- 
    index_resize_ack_8101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_index_0_resize_ack_0, ack => cp_elements(214)); -- 
    scale_rr_8105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(214), ack => array_obj_ref_1864_index_0_scale_req_0); -- 
    scale_ra_8106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_index_0_scale_ack_0, ack => cp_elements(215)); -- 
    scale_cr_8107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => array_obj_ref_1864_index_0_scale_req_1); -- 
    scale_ca_8108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_index_0_scale_ack_1, ack => cp_elements(216)); -- 
    partial_sum_1_rr_8112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(216), ack => array_obj_ref_1864_index_sum_1_req_0); -- 
    partial_sum_1_ra_8113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_index_sum_1_ack_0, ack => cp_elements(217)); -- 
    partial_sum_1_cr_8114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => array_obj_ref_1864_index_sum_1_req_1); -- 
    partial_sum_1_ca_8115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_index_sum_1_ack_1, ack => cp_elements(218)); -- 
    final_index_req_8116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => array_obj_ref_1864_offset_inst_req_0); -- 
    final_index_ack_8117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_offset_inst_ack_0, ack => cp_elements(219)); -- 
    sum_rename_req_8121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => array_obj_ref_1864_root_address_inst_req_0); -- 
    sum_rename_ack_8122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1864_root_address_inst_ack_0, ack => cp_elements(220)); -- 
    final_reg_ack_8127_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_1865_final_reg_ack_0, ack => cp_elements(221)); -- 
    base_resize_req_8140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => ptr_deref_1869_base_resize_req_0); -- 
    base_resize_ack_8141_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_base_resize_ack_0, ack => cp_elements(222)); -- 
    sum_rename_req_8145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_1869_root_address_inst_req_0); -- 
    sum_rename_ack_8146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_root_address_inst_ack_0, ack => cp_elements(223)); -- 
    root_rename_req_8150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => ptr_deref_1869_addr_0_req_0); -- 
    root_rename_ack_8151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_addr_0_ack_0, ack => cp_elements(224)); -- 
    rr_8161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_1869_load_0_req_0); -- 
    ra_8162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_load_0_ack_0, ack => cp_elements(225)); -- 
    cr_8172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => ptr_deref_1869_load_0_req_1); -- 
    ca_8173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_load_0_ack_1, ack => cp_elements(226)); -- 
    merge_req_8174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => ptr_deref_1869_gather_scatter_req_0); -- 
    merge_ack_8175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1869_gather_scatter_ack_0, ack => cp_elements(227)); -- 
    cpelement_group_228 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(227) & cp_elements(229));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(228),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_1875_inst_req_0); -- 
    cp_elements(229) <= cp_elements(210);
    ra_8185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_0, ack => cp_elements(230)); -- 
    cr_8186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => binary_1875_inst_req_1); -- 
    ca_8187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1875_inst_ack_1, ack => cp_elements(231)); -- 
    cp_elements(232) <= cp_elements(231);
    cp_elements(233) <= false;
    cp_elements(234) <= cp_elements(233);
    cp_elements(235) <= cp_elements(231);
    branch_req_8195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => if_stmt_1877_branch_req_0); -- 
    cp_elements(236) <= cp_elements(235);
    cp_elements(237) <= cp_elements(236);
    if_choice_transition_8200_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1877_branch_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(236);
    cp_elements(240) <= if_stmt_1877_branch_ack_0;
    cp_elements(241) <= cp_elements(7);
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(243) & cp_elements(251));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => addr_of_1889_final_reg_req_0); -- 
    cp_elements(243) <= cp_elements(241);
    cp_elements(244) <= cp_elements(241);
    index_resize_req_8223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => array_obj_ref_1888_index_0_resize_req_0); -- 
    index_resize_ack_8224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_index_0_resize_ack_0, ack => cp_elements(245)); -- 
    scale_rr_8228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(245), ack => array_obj_ref_1888_index_0_scale_req_0); -- 
    scale_ra_8229_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_index_0_scale_ack_0, ack => cp_elements(246)); -- 
    scale_cr_8230_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => array_obj_ref_1888_index_0_scale_req_1); -- 
    scale_ca_8231_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_index_0_scale_ack_1, ack => cp_elements(247)); -- 
    partial_sum_1_rr_8235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(247), ack => array_obj_ref_1888_index_sum_1_req_0); -- 
    partial_sum_1_ra_8236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_index_sum_1_ack_0, ack => cp_elements(248)); -- 
    partial_sum_1_cr_8237_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => array_obj_ref_1888_index_sum_1_req_1); -- 
    partial_sum_1_ca_8238_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_index_sum_1_ack_1, ack => cp_elements(249)); -- 
    final_index_req_8239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => array_obj_ref_1888_offset_inst_req_0); -- 
    final_index_ack_8240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_offset_inst_ack_0, ack => cp_elements(250)); -- 
    sum_rename_req_8244_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => array_obj_ref_1888_root_address_inst_req_0); -- 
    sum_rename_ack_8245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1888_root_address_inst_ack_0, ack => cp_elements(251)); -- 
    cp_elements(252) <= addr_of_1889_final_reg_ack_0;
    cp_elements(253) <= cp_elements(993);
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(255) & cp_elements(256));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8262_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => binary_1904_inst_req_0); -- 
    cp_elements(255) <= cp_elements(253);
    cp_elements(256) <= cp_elements(253);
    ra_8263_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1904_inst_ack_0, ack => cp_elements(257)); -- 
    cr_8264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => binary_1904_inst_req_1); -- 
    ca_8265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1904_inst_ack_1, ack => cp_elements(258)); -- 
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(258) & cp_elements(260));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => binary_1910_inst_req_0); -- 
    cp_elements(260) <= cp_elements(253);
    ra_8275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1910_inst_ack_0, ack => cp_elements(261)); -- 
    cr_8276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => binary_1910_inst_req_1); -- 
    ca_8277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1910_inst_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(262);
    cp_elements(264) <= false;
    cp_elements(265) <= cp_elements(264);
    cp_elements(266) <= cp_elements(262);
    branch_req_8285_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => if_stmt_1912_branch_req_0); -- 
    cp_elements(267) <= cp_elements(266);
    cp_elements(268) <= cp_elements(267);
    if_choice_transition_8290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1912_branch_ack_1, ack => cp_elements(269)); -- 
    cp_elements(270) <= cp_elements(267);
    else_choice_transition_8294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1912_branch_ack_0, ack => cp_elements(271)); -- 
    cp_elements(272) <= cp_elements(8);
    cpelement_group_273 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(275));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(273),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => binary_1923_inst_req_0); -- 
    cp_elements(274) <= cp_elements(272);
    cp_elements(275) <= cp_elements(272);
    ra_8309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1923_inst_ack_0, ack => cp_elements(276)); -- 
    cr_8310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(276), ack => binary_1923_inst_req_1); -- 
    ca_8311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1923_inst_ack_1, ack => cp_elements(277)); -- 
    cp_elements(278) <= cp_elements(277);
    cp_elements(279) <= false;
    cp_elements(280) <= cp_elements(279);
    cp_elements(281) <= cp_elements(277);
    branch_req_8319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => if_stmt_1925_branch_req_0); -- 
    cp_elements(282) <= cp_elements(281);
    cp_elements(283) <= cp_elements(282);
    if_choice_transition_8324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1925_branch_ack_1, ack => cp_elements(284)); -- 
    cp_elements(285) <= cp_elements(282);
    else_choice_transition_8328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1925_branch_ack_0, ack => cp_elements(286)); -- 
    cp_elements(287) <= cp_elements(286);
    cp_elements(288) <= cp_elements(287);
    cpelement_group_289 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(288) & cp_elements(296));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(289),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => array_obj_ref_1937_final_reg_req_0); -- 
    cp_elements(290) <= cp_elements(287);
    base_resize_req_8351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => array_obj_ref_1937_base_resize_req_0); -- 
    cp_elements(291) <= cp_elements(287);
    final_index_req_8345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(291), ack => array_obj_ref_1937_offset_inst_req_0); -- 
    final_index_ack_8346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1937_offset_inst_ack_0, ack => cp_elements(292)); -- 
    base_resize_ack_8352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1937_base_resize_ack_0, ack => cp_elements(293)); -- 
    cpelement_group_294 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(292) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(294),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_8357_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => array_obj_ref_1937_root_address_inst_req_0); -- 
    plus_base_ra_8358_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1937_root_address_inst_ack_0, ack => cp_elements(295)); -- 
    plus_base_cr_8359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => array_obj_ref_1937_root_address_inst_req_1); -- 
    plus_base_ca_8360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1937_root_address_inst_ack_1, ack => cp_elements(296)); -- 
    final_reg_ack_8365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1937_final_reg_ack_0, ack => cp_elements(297)); -- 
    base_resize_req_8378_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(297), ack => ptr_deref_1940_base_resize_req_0); -- 
    cp_elements(298) <= cp_elements(287);
    cpelement_group_299 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(298) & cp_elements(302));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(299),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(299), ack => ptr_deref_1940_gather_scatter_req_0); -- 
    base_resize_ack_8379_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1940_base_resize_ack_0, ack => cp_elements(300)); -- 
    sum_rename_req_8383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => ptr_deref_1940_root_address_inst_req_0); -- 
    sum_rename_ack_8384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1940_root_address_inst_ack_0, ack => cp_elements(301)); -- 
    root_rename_req_8388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => ptr_deref_1940_addr_0_req_0); -- 
    root_rename_ack_8389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1940_addr_0_ack_0, ack => cp_elements(302)); -- 
    split_ack_8394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1940_gather_scatter_ack_0, ack => cp_elements(303)); -- 
    rr_8401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(303), ack => ptr_deref_1940_store_0_req_0); -- 
    cp_elements(304) <= ptr_deref_1940_store_0_ack_0;
    cp_elements(305) <= cp_elements(304);
    cr_8412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(305), ack => ptr_deref_1940_store_0_req_1); -- 
    ca_8413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1940_store_0_ack_1, ack => cp_elements(306)); -- 
    cp_elements(307) <= cp_elements(287);
    cpelement_group_308 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(307) & cp_elements(312));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(308),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => array_obj_ref_1947_final_reg_req_0); -- 
    cp_elements(309) <= cp_elements(287);
    base_resize_req_8424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => array_obj_ref_1947_base_resize_req_0); -- 
    base_resize_ack_8425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1947_base_resize_ack_0, ack => cp_elements(310)); -- 
    plus_base_rr_8430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(310), ack => array_obj_ref_1947_root_address_inst_req_0); -- 
    plus_base_ra_8431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1947_root_address_inst_ack_0, ack => cp_elements(311)); -- 
    plus_base_cr_8432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => array_obj_ref_1947_root_address_inst_req_1); -- 
    plus_base_ca_8433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1947_root_address_inst_ack_1, ack => cp_elements(312)); -- 
    final_reg_ack_8438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1947_final_reg_ack_0, ack => cp_elements(313)); -- 
    cpelement_group_314 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(313) & cp_elements(315));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(314),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8447_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(314), ack => type_cast_1951_inst_req_0); -- 
    cp_elements(315) <= cp_elements(287);
    cp_elements(316) <= type_cast_1951_inst_ack_0;
    cp_elements(317) <= cp_elements(287);
    cpelement_group_318 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(304) & cp_elements(316) & cp_elements(317) & cp_elements(334));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(318),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(318), ack => ptr_deref_1954_gather_scatter_req_0); -- 
    cp_elements(319) <= cp_elements(316);
    base_resize_req_8461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => ptr_deref_1954_base_resize_req_0); -- 
    base_resize_ack_8462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_base_resize_ack_0, ack => cp_elements(320)); -- 
    sum_rename_req_8466_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(320), ack => ptr_deref_1954_root_address_inst_req_0); -- 
    cp_elements(321) <= ptr_deref_1954_root_address_inst_ack_0;
    cp_elements(322) <= cp_elements(321);
    rr_8474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => ptr_deref_1954_addr_0_req_0); -- 
    ra_8475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_0_ack_0, ack => cp_elements(323)); -- 
    cr_8476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => ptr_deref_1954_addr_0_req_1); -- 
    ca_8477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_0_ack_1, ack => cp_elements(324)); -- 
    cp_elements(325) <= cp_elements(321);
    rr_8481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => ptr_deref_1954_addr_1_req_0); -- 
    ra_8482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_1_ack_0, ack => cp_elements(326)); -- 
    cr_8483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(326), ack => ptr_deref_1954_addr_1_req_1); -- 
    ca_8484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_1_ack_1, ack => cp_elements(327)); -- 
    cp_elements(328) <= cp_elements(321);
    rr_8488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(328), ack => ptr_deref_1954_addr_2_req_0); -- 
    ra_8489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_2_ack_0, ack => cp_elements(329)); -- 
    cr_8490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(329), ack => ptr_deref_1954_addr_2_req_1); -- 
    ca_8491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_2_ack_1, ack => cp_elements(330)); -- 
    cp_elements(331) <= cp_elements(321);
    rr_8495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => ptr_deref_1954_addr_3_req_0); -- 
    ra_8496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_3_ack_0, ack => cp_elements(332)); -- 
    cr_8497_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(332), ack => ptr_deref_1954_addr_3_req_1); -- 
    ca_8498_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_addr_3_ack_1, ack => cp_elements(333)); -- 
    cpelement_group_334 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(324) & cp_elements(327) & cp_elements(330) & cp_elements(333));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(334),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(335) <= ptr_deref_1954_gather_scatter_ack_0;
    cp_elements(336) <= cp_elements(335);
    rr_8510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(336), ack => ptr_deref_1954_store_0_req_0); -- 
    ra_8511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_0_ack_0, ack => cp_elements(337)); -- 
    cp_elements(338) <= cp_elements(335);
    rr_8515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(338), ack => ptr_deref_1954_store_1_req_0); -- 
    ra_8516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_1_ack_0, ack => cp_elements(339)); -- 
    cp_elements(340) <= cp_elements(335);
    rr_8520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(340), ack => ptr_deref_1954_store_2_req_0); -- 
    ra_8521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_2_ack_0, ack => cp_elements(341)); -- 
    cp_elements(342) <= cp_elements(335);
    rr_8525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => ptr_deref_1954_store_3_req_0); -- 
    ra_8526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_3_ack_0, ack => cp_elements(343)); -- 
    cpelement_group_344 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(337) & cp_elements(339) & cp_elements(341) & cp_elements(343));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(344),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(345) <= cp_elements(344);
    cp_elements(346) <= cp_elements(345);
    cr_8536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(346), ack => ptr_deref_1954_store_0_req_1); -- 
    ca_8537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_0_ack_1, ack => cp_elements(347)); -- 
    cp_elements(348) <= cp_elements(345);
    cr_8541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(348), ack => ptr_deref_1954_store_1_req_1); -- 
    ca_8542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_1_ack_1, ack => cp_elements(349)); -- 
    cp_elements(350) <= cp_elements(345);
    cr_8546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => ptr_deref_1954_store_2_req_1); -- 
    ca_8547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_2_ack_1, ack => cp_elements(351)); -- 
    cp_elements(352) <= cp_elements(345);
    cr_8551_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(352), ack => ptr_deref_1954_store_3_req_1); -- 
    ca_8552_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1954_store_3_ack_1, ack => cp_elements(353)); -- 
    cpelement_group_354 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(347) & cp_elements(349) & cp_elements(351) & cp_elements(353));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(354),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(355) <= cp_elements(287);
    cpelement_group_356 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(355) & cp_elements(360));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(356),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(356), ack => array_obj_ref_1961_final_reg_req_0); -- 
    cp_elements(357) <= cp_elements(287);
    base_resize_req_8563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => array_obj_ref_1961_base_resize_req_0); -- 
    base_resize_ack_8564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_base_resize_ack_0, ack => cp_elements(358)); -- 
    plus_base_rr_8569_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => array_obj_ref_1961_root_address_inst_req_0); -- 
    plus_base_ra_8570_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_root_address_inst_ack_0, ack => cp_elements(359)); -- 
    plus_base_cr_8571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(359), ack => array_obj_ref_1961_root_address_inst_req_1); -- 
    plus_base_ca_8572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_root_address_inst_ack_1, ack => cp_elements(360)); -- 
    final_reg_ack_8577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1961_final_reg_ack_0, ack => cp_elements(361)); -- 
    cpelement_group_362 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(361) & cp_elements(363));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(362),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(362), ack => type_cast_1965_inst_req_0); -- 
    cp_elements(363) <= cp_elements(287);
    ack_8587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1965_inst_ack_0, ack => cp_elements(364)); -- 
    cpelement_group_365 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(366) & cp_elements(367));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(365),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(365), ack => type_cast_1969_inst_req_0); -- 
    cp_elements(366) <= cp_elements(287);
    cp_elements(367) <= cp_elements(287);
    cp_elements(368) <= type_cast_1969_inst_ack_0;
    cp_elements(369) <= cp_elements(287);
    cpelement_group_370 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(344) & cp_elements(368) & cp_elements(369) & cp_elements(386));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(370),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(370), ack => ptr_deref_1972_gather_scatter_req_0); -- 
    cp_elements(371) <= cp_elements(368);
    base_resize_req_8610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(371), ack => ptr_deref_1972_base_resize_req_0); -- 
    base_resize_ack_8611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_base_resize_ack_0, ack => cp_elements(372)); -- 
    sum_rename_req_8615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(372), ack => ptr_deref_1972_root_address_inst_req_0); -- 
    cp_elements(373) <= ptr_deref_1972_root_address_inst_ack_0;
    cp_elements(374) <= cp_elements(373);
    rr_8623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(374), ack => ptr_deref_1972_addr_0_req_0); -- 
    ra_8624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_0_ack_0, ack => cp_elements(375)); -- 
    cr_8625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(375), ack => ptr_deref_1972_addr_0_req_1); -- 
    ca_8626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_0_ack_1, ack => cp_elements(376)); -- 
    cp_elements(377) <= cp_elements(373);
    rr_8630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(377), ack => ptr_deref_1972_addr_1_req_0); -- 
    ra_8631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_1_ack_0, ack => cp_elements(378)); -- 
    cr_8632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(378), ack => ptr_deref_1972_addr_1_req_1); -- 
    ca_8633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_1_ack_1, ack => cp_elements(379)); -- 
    cp_elements(380) <= cp_elements(373);
    rr_8637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => ptr_deref_1972_addr_2_req_0); -- 
    ra_8638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_2_ack_0, ack => cp_elements(381)); -- 
    cr_8639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => ptr_deref_1972_addr_2_req_1); -- 
    ca_8640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_2_ack_1, ack => cp_elements(382)); -- 
    cp_elements(383) <= cp_elements(373);
    rr_8644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(383), ack => ptr_deref_1972_addr_3_req_0); -- 
    ra_8645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_3_ack_0, ack => cp_elements(384)); -- 
    cr_8646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => ptr_deref_1972_addr_3_req_1); -- 
    ca_8647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_addr_3_ack_1, ack => cp_elements(385)); -- 
    cpelement_group_386 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(376) & cp_elements(379) & cp_elements(382) & cp_elements(385));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(386),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(387) <= ptr_deref_1972_gather_scatter_ack_0;
    cp_elements(388) <= cp_elements(387);
    rr_8659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(388), ack => ptr_deref_1972_store_0_req_0); -- 
    ra_8660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_0_ack_0, ack => cp_elements(389)); -- 
    cp_elements(390) <= cp_elements(387);
    rr_8664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(390), ack => ptr_deref_1972_store_1_req_0); -- 
    ra_8665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_1_ack_0, ack => cp_elements(391)); -- 
    cp_elements(392) <= cp_elements(387);
    rr_8669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(392), ack => ptr_deref_1972_store_2_req_0); -- 
    ra_8670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_2_ack_0, ack => cp_elements(393)); -- 
    cp_elements(394) <= cp_elements(387);
    rr_8674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => ptr_deref_1972_store_3_req_0); -- 
    ra_8675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_3_ack_0, ack => cp_elements(395)); -- 
    cpelement_group_396 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(389) & cp_elements(391) & cp_elements(393) & cp_elements(395));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(396),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(397) <= cp_elements(396);
    cr_8685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(397), ack => ptr_deref_1972_store_0_req_1); -- 
    ca_8686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_0_ack_1, ack => cp_elements(398)); -- 
    cp_elements(399) <= cp_elements(396);
    cr_8690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(399), ack => ptr_deref_1972_store_1_req_1); -- 
    ca_8691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_1_ack_1, ack => cp_elements(400)); -- 
    cp_elements(401) <= cp_elements(396);
    cr_8695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(401), ack => ptr_deref_1972_store_2_req_1); -- 
    ca_8696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_2_ack_1, ack => cp_elements(402)); -- 
    cp_elements(403) <= cp_elements(396);
    cr_8700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(403), ack => ptr_deref_1972_store_3_req_1); -- 
    ca_8701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_1972_store_3_ack_1, ack => cp_elements(404)); -- 
    cpelement_group_405 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(398) & cp_elements(400) & cp_elements(402) & cp_elements(404));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(405),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_406 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(407) & cp_elements(408));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(406),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_8710_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(406), ack => type_cast_1978_inst_req_0); -- 
    cp_elements(407) <= cp_elements(287);
    cp_elements(408) <= cp_elements(287);
    ack_8711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1978_inst_ack_0, ack => cp_elements(409)); -- 
    base_resize_req_8722_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(409), ack => array_obj_ref_1987_base_resize_req_0); -- 
    cp_elements(410) <= cp_elements(287);
    cpelement_group_411 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(410) & cp_elements(414));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(411),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_8735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(411), ack => array_obj_ref_1987_final_reg_req_0); -- 
    base_resize_ack_8723_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1987_base_resize_ack_0, ack => cp_elements(412)); -- 
    plus_base_rr_8728_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(412), ack => array_obj_ref_1987_root_address_inst_req_0); -- 
    plus_base_ra_8729_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1987_root_address_inst_ack_0, ack => cp_elements(413)); -- 
    plus_base_cr_8730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(413), ack => array_obj_ref_1987_root_address_inst_req_1); -- 
    plus_base_ca_8731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1987_root_address_inst_ack_1, ack => cp_elements(414)); -- 
    final_reg_ack_8736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1987_final_reg_ack_0, ack => cp_elements(415)); -- 
    cpelement_group_416 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(415) & cp_elements(417));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(416),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8745_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(416), ack => binary_1993_inst_req_0); -- 
    cp_elements(417) <= cp_elements(287);
    ra_8746_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1993_inst_ack_0, ack => cp_elements(418)); -- 
    cr_8747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(418), ack => binary_1993_inst_req_1); -- 
    ca_8748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_1993_inst_ack_1, ack => cp_elements(419)); -- 
    cpelement_group_420 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(306) & cp_elements(354) & cp_elements(364) & cp_elements(405) & cp_elements(419));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(420),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(421) <= cp_elements(10);
    cp_elements(422) <= false;
    cp_elements(423) <= cp_elements(422);
    cp_elements(424) <= cp_elements(10);
    branch_req_8756_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(424), ack => if_stmt_1995_branch_req_0); -- 
    cp_elements(425) <= cp_elements(424);
    cp_elements(426) <= cp_elements(425);
    if_choice_transition_8761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1995_branch_ack_1, ack => cp_elements(427)); -- 
    cp_elements(428) <= cp_elements(425);
    else_choice_transition_8765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1995_branch_ack_0, ack => cp_elements(429)); -- 
    cp_elements(430) <= cp_elements(11);
    cp_elements(431) <= cp_elements(430);
    cpelement_group_432 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(431) & cp_elements(433) & cp_elements(437));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(432),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8798_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(432), ack => ptr_deref_2003_gather_scatter_req_0); -- 
    cp_elements(433) <= cp_elements(430);
    cp_elements(434) <= cp_elements(433);
    base_resize_req_8783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(434), ack => ptr_deref_2003_base_resize_req_0); -- 
    base_resize_ack_8784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_base_resize_ack_0, ack => cp_elements(435)); -- 
    sum_rename_req_8788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(435), ack => ptr_deref_2003_root_address_inst_req_0); -- 
    sum_rename_ack_8789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_root_address_inst_ack_0, ack => cp_elements(436)); -- 
    root_rename_req_8793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(436), ack => ptr_deref_2003_addr_0_req_0); -- 
    root_rename_ack_8794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_addr_0_ack_0, ack => cp_elements(437)); -- 
    split_ack_8799_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_gather_scatter_ack_0, ack => cp_elements(438)); -- 
    rr_8806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(438), ack => ptr_deref_2003_store_0_req_0); -- 
    ra_8807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_store_0_ack_0, ack => cp_elements(439)); -- 
    cr_8817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(439), ack => ptr_deref_2003_store_0_req_1); -- 
    ca_8818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2003_store_0_ack_1, ack => cp_elements(440)); -- 
    cp_elements(441) <= cp_elements(1001);
    cp_elements(442) <= cp_elements(441);
    base_resize_req_8834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(442), ack => ptr_deref_2011_base_resize_req_0); -- 
    base_resize_ack_8835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_base_resize_ack_0, ack => cp_elements(443)); -- 
    sum_rename_req_8839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(443), ack => ptr_deref_2011_root_address_inst_req_0); -- 
    cp_elements(444) <= ptr_deref_2011_root_address_inst_ack_0;
    cp_elements(445) <= cp_elements(444);
    rr_8847_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => ptr_deref_2011_addr_0_req_0); -- 
    ra_8848_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_0_ack_0, ack => cp_elements(446)); -- 
    cr_8849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(446), ack => ptr_deref_2011_addr_0_req_1); -- 
    ca_8850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_0_ack_1, ack => cp_elements(447)); -- 
    cp_elements(448) <= cp_elements(444);
    rr_8854_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(448), ack => ptr_deref_2011_addr_1_req_0); -- 
    ra_8855_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_1_ack_0, ack => cp_elements(449)); -- 
    cr_8856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => ptr_deref_2011_addr_1_req_1); -- 
    ca_8857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_1_ack_1, ack => cp_elements(450)); -- 
    cp_elements(451) <= cp_elements(444);
    rr_8861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(451), ack => ptr_deref_2011_addr_2_req_0); -- 
    ra_8862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_2_ack_0, ack => cp_elements(452)); -- 
    cr_8863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(452), ack => ptr_deref_2011_addr_2_req_1); -- 
    ca_8864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_2_ack_1, ack => cp_elements(453)); -- 
    cp_elements(454) <= cp_elements(444);
    rr_8868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(454), ack => ptr_deref_2011_addr_3_req_0); -- 
    ra_8869_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_3_ack_0, ack => cp_elements(455)); -- 
    cr_8870_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(455), ack => ptr_deref_2011_addr_3_req_1); -- 
    ca_8871_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_addr_3_ack_1, ack => cp_elements(456)); -- 
    cpelement_group_457 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(447) & cp_elements(450) & cp_elements(453) & cp_elements(456));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(457),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(458) <= cp_elements(457);
    rr_8881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(458), ack => ptr_deref_2011_load_0_req_0); -- 
    ra_8882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_0_ack_0, ack => cp_elements(459)); -- 
    cp_elements(460) <= cp_elements(457);
    rr_8886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(460), ack => ptr_deref_2011_load_1_req_0); -- 
    ra_8887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_1_ack_0, ack => cp_elements(461)); -- 
    cp_elements(462) <= cp_elements(457);
    rr_8891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(462), ack => ptr_deref_2011_load_2_req_0); -- 
    ra_8892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_2_ack_0, ack => cp_elements(463)); -- 
    cp_elements(464) <= cp_elements(457);
    rr_8896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(464), ack => ptr_deref_2011_load_3_req_0); -- 
    ra_8897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_3_ack_0, ack => cp_elements(465)); -- 
    cpelement_group_466 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(459) & cp_elements(461) & cp_elements(463) & cp_elements(465));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(466),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(467) <= cp_elements(466);
    cr_8907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => ptr_deref_2011_load_0_req_1); -- 
    ca_8908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_0_ack_1, ack => cp_elements(468)); -- 
    cp_elements(469) <= cp_elements(466);
    cr_8912_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => ptr_deref_2011_load_1_req_1); -- 
    ca_8913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_1_ack_1, ack => cp_elements(470)); -- 
    cp_elements(471) <= cp_elements(466);
    cr_8917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(471), ack => ptr_deref_2011_load_2_req_1); -- 
    ca_8918_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_2_ack_1, ack => cp_elements(472)); -- 
    cp_elements(473) <= cp_elements(466);
    cr_8922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(473), ack => ptr_deref_2011_load_3_req_1); -- 
    ca_8923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_load_3_ack_1, ack => cp_elements(474)); -- 
    cpelement_group_475 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(468) & cp_elements(470) & cp_elements(472) & cp_elements(474));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(475),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_8924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(475), ack => ptr_deref_2011_gather_scatter_req_0); -- 
    merge_ack_8925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2011_gather_scatter_ack_0, ack => cp_elements(476)); -- 
    cpelement_group_477 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(476) & cp_elements(478));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(477),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_8934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(477), ack => binary_2017_inst_req_0); -- 
    cp_elements(478) <= cp_elements(441);
    ra_8935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2017_inst_ack_0, ack => cp_elements(479)); -- 
    cr_8936_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(479), ack => binary_2017_inst_req_1); -- 
    ca_8937_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2017_inst_ack_1, ack => cp_elements(480)); -- 
    cpelement_group_481 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(480) & cp_elements(482) & cp_elements(498));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(481),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_8992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(481), ack => ptr_deref_2020_gather_scatter_req_0); -- 
    cp_elements(482) <= cp_elements(441);
    cp_elements(483) <= cp_elements(482);
    base_resize_req_8951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(483), ack => ptr_deref_2020_base_resize_req_0); -- 
    base_resize_ack_8952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_base_resize_ack_0, ack => cp_elements(484)); -- 
    sum_rename_req_8956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(484), ack => ptr_deref_2020_root_address_inst_req_0); -- 
    cp_elements(485) <= ptr_deref_2020_root_address_inst_ack_0;
    cp_elements(486) <= cp_elements(485);
    rr_8964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(486), ack => ptr_deref_2020_addr_0_req_0); -- 
    ra_8965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_0_ack_0, ack => cp_elements(487)); -- 
    cr_8966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(487), ack => ptr_deref_2020_addr_0_req_1); -- 
    ca_8967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_0_ack_1, ack => cp_elements(488)); -- 
    cp_elements(489) <= cp_elements(485);
    rr_8971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(489), ack => ptr_deref_2020_addr_1_req_0); -- 
    ra_8972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_1_ack_0, ack => cp_elements(490)); -- 
    cr_8973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(490), ack => ptr_deref_2020_addr_1_req_1); -- 
    ca_8974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_1_ack_1, ack => cp_elements(491)); -- 
    cp_elements(492) <= cp_elements(485);
    rr_8978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(492), ack => ptr_deref_2020_addr_2_req_0); -- 
    ra_8979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_2_ack_0, ack => cp_elements(493)); -- 
    cr_8980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(493), ack => ptr_deref_2020_addr_2_req_1); -- 
    ca_8981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_2_ack_1, ack => cp_elements(494)); -- 
    cp_elements(495) <= cp_elements(485);
    rr_8985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(495), ack => ptr_deref_2020_addr_3_req_0); -- 
    ra_8986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_3_ack_0, ack => cp_elements(496)); -- 
    cr_8987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(496), ack => ptr_deref_2020_addr_3_req_1); -- 
    ca_8988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_addr_3_ack_1, ack => cp_elements(497)); -- 
    cpelement_group_498 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(488) & cp_elements(491) & cp_elements(494) & cp_elements(497));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(498),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(499) <= ptr_deref_2020_gather_scatter_ack_0;
    cp_elements(500) <= cp_elements(499);
    rr_9000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(500), ack => ptr_deref_2020_store_0_req_0); -- 
    ra_9001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_0_ack_0, ack => cp_elements(501)); -- 
    cp_elements(502) <= cp_elements(499);
    rr_9005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(502), ack => ptr_deref_2020_store_1_req_0); -- 
    ra_9006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_1_ack_0, ack => cp_elements(503)); -- 
    cp_elements(504) <= cp_elements(499);
    rr_9010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(504), ack => ptr_deref_2020_store_2_req_0); -- 
    ra_9011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_2_ack_0, ack => cp_elements(505)); -- 
    cp_elements(506) <= cp_elements(499);
    rr_9015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(506), ack => ptr_deref_2020_store_3_req_0); -- 
    ra_9016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_3_ack_0, ack => cp_elements(507)); -- 
    cpelement_group_508 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(501) & cp_elements(503) & cp_elements(505) & cp_elements(507));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(508),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(509) <= cp_elements(508);
    cp_elements(510) <= cp_elements(509);
    cr_9026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(510), ack => ptr_deref_2020_store_0_req_1); -- 
    ca_9027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_0_ack_1, ack => cp_elements(511)); -- 
    cp_elements(512) <= cp_elements(509);
    cr_9031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(512), ack => ptr_deref_2020_store_1_req_1); -- 
    ca_9032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_1_ack_1, ack => cp_elements(513)); -- 
    cp_elements(514) <= cp_elements(509);
    cr_9036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(514), ack => ptr_deref_2020_store_2_req_1); -- 
    ca_9037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_2_ack_1, ack => cp_elements(515)); -- 
    cp_elements(516) <= cp_elements(509);
    cr_9041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(516), ack => ptr_deref_2020_store_3_req_1); -- 
    ca_9042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2020_store_3_ack_1, ack => cp_elements(517)); -- 
    cpelement_group_518 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(511) & cp_elements(513) & cp_elements(515) & cp_elements(517));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(518),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_519 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(508) & cp_elements(520) & cp_elements(536));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(519),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(520) <= cp_elements(441);
    cp_elements(521) <= cp_elements(520);
    base_resize_req_9055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(521), ack => ptr_deref_2025_base_resize_req_0); -- 
    base_resize_ack_9056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_base_resize_ack_0, ack => cp_elements(522)); -- 
    sum_rename_req_9060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(522), ack => ptr_deref_2025_root_address_inst_req_0); -- 
    cp_elements(523) <= ptr_deref_2025_root_address_inst_ack_0;
    cp_elements(524) <= cp_elements(523);
    rr_9068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(524), ack => ptr_deref_2025_addr_0_req_0); -- 
    ra_9069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_0_ack_0, ack => cp_elements(525)); -- 
    cr_9070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(525), ack => ptr_deref_2025_addr_0_req_1); -- 
    ca_9071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_0_ack_1, ack => cp_elements(526)); -- 
    cp_elements(527) <= cp_elements(523);
    rr_9075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(527), ack => ptr_deref_2025_addr_1_req_0); -- 
    ra_9076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_1_ack_0, ack => cp_elements(528)); -- 
    cr_9077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(528), ack => ptr_deref_2025_addr_1_req_1); -- 
    ca_9078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_1_ack_1, ack => cp_elements(529)); -- 
    cp_elements(530) <= cp_elements(523);
    rr_9082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(530), ack => ptr_deref_2025_addr_2_req_0); -- 
    ra_9083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_2_ack_0, ack => cp_elements(531)); -- 
    cr_9084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(531), ack => ptr_deref_2025_addr_2_req_1); -- 
    ca_9085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_2_ack_1, ack => cp_elements(532)); -- 
    cp_elements(533) <= cp_elements(523);
    rr_9089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(533), ack => ptr_deref_2025_addr_3_req_0); -- 
    ra_9090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_3_ack_0, ack => cp_elements(534)); -- 
    cr_9091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(534), ack => ptr_deref_2025_addr_3_req_1); -- 
    ca_9092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_addr_3_ack_1, ack => cp_elements(535)); -- 
    cpelement_group_536 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(526) & cp_elements(529) & cp_elements(532) & cp_elements(535));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(536),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(537) <= cp_elements(519);
    rr_9102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(537), ack => ptr_deref_2025_load_0_req_0); -- 
    ra_9103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_0_ack_0, ack => cp_elements(538)); -- 
    cp_elements(539) <= cp_elements(519);
    rr_9107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(539), ack => ptr_deref_2025_load_1_req_0); -- 
    ra_9108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_1_ack_0, ack => cp_elements(540)); -- 
    cp_elements(541) <= cp_elements(519);
    rr_9112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => ptr_deref_2025_load_2_req_0); -- 
    ra_9113_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_2_ack_0, ack => cp_elements(542)); -- 
    cp_elements(543) <= cp_elements(519);
    rr_9117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(543), ack => ptr_deref_2025_load_3_req_0); -- 
    ra_9118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_3_ack_0, ack => cp_elements(544)); -- 
    cpelement_group_545 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(538) & cp_elements(540) & cp_elements(542) & cp_elements(544));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(545),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(546) <= cp_elements(545);
    cr_9128_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(546), ack => ptr_deref_2025_load_0_req_1); -- 
    ca_9129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_0_ack_1, ack => cp_elements(547)); -- 
    cp_elements(548) <= cp_elements(545);
    cr_9133_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => ptr_deref_2025_load_1_req_1); -- 
    ca_9134_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_1_ack_1, ack => cp_elements(549)); -- 
    cp_elements(550) <= cp_elements(545);
    cr_9138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => ptr_deref_2025_load_2_req_1); -- 
    ca_9139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_2_ack_1, ack => cp_elements(551)); -- 
    cp_elements(552) <= cp_elements(545);
    cr_9143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => ptr_deref_2025_load_3_req_1); -- 
    ca_9144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_load_3_ack_1, ack => cp_elements(553)); -- 
    cpelement_group_554 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(547) & cp_elements(549) & cp_elements(551) & cp_elements(553));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(554),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => ptr_deref_2025_gather_scatter_req_0); -- 
    merge_ack_9146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2025_gather_scatter_ack_0, ack => cp_elements(555)); -- 
    cpelement_group_556 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(555) & cp_elements(557));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(556),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9155_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => binary_2031_inst_req_0); -- 
    cp_elements(557) <= cp_elements(441);
    ra_9156_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2031_inst_ack_0, ack => cp_elements(558)); -- 
    cr_9157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(558), ack => binary_2031_inst_req_1); -- 
    ca_9158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2031_inst_ack_1, ack => cp_elements(559)); -- 
    cpelement_group_560 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(518) & cp_elements(559));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(560),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(561) <= cp_elements(12);
    cp_elements(562) <= false;
    cp_elements(563) <= cp_elements(562);
    cp_elements(564) <= cp_elements(12);
    branch_req_9166_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => if_stmt_2033_branch_req_0); -- 
    cp_elements(565) <= cp_elements(564);
    cp_elements(566) <= cp_elements(565);
    if_choice_transition_9171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2033_branch_ack_1, ack => cp_elements(567)); -- 
    cp_elements(568) <= cp_elements(565);
    else_choice_transition_9175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2033_branch_ack_0, ack => cp_elements(569)); -- 
    cp_elements(570) <= cp_elements(13);
    cp_elements(571) <= cp_elements(570);
    base_resize_req_9193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(571), ack => ptr_deref_2042_base_resize_req_0); -- 
    base_resize_ack_9194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_base_resize_ack_0, ack => cp_elements(572)); -- 
    sum_rename_req_9198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(572), ack => ptr_deref_2042_root_address_inst_req_0); -- 
    cp_elements(573) <= ptr_deref_2042_root_address_inst_ack_0;
    cp_elements(574) <= cp_elements(573);
    rr_9206_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(574), ack => ptr_deref_2042_addr_0_req_0); -- 
    ra_9207_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_0_ack_0, ack => cp_elements(575)); -- 
    cr_9208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(575), ack => ptr_deref_2042_addr_0_req_1); -- 
    ca_9209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_0_ack_1, ack => cp_elements(576)); -- 
    cp_elements(577) <= cp_elements(573);
    rr_9213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(577), ack => ptr_deref_2042_addr_1_req_0); -- 
    ra_9214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_1_ack_0, ack => cp_elements(578)); -- 
    cr_9215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(578), ack => ptr_deref_2042_addr_1_req_1); -- 
    ca_9216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_1_ack_1, ack => cp_elements(579)); -- 
    cp_elements(580) <= cp_elements(573);
    rr_9220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(580), ack => ptr_deref_2042_addr_2_req_0); -- 
    ra_9221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_2_ack_0, ack => cp_elements(581)); -- 
    cr_9222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(581), ack => ptr_deref_2042_addr_2_req_1); -- 
    ca_9223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_2_ack_1, ack => cp_elements(582)); -- 
    cp_elements(583) <= cp_elements(573);
    rr_9227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(583), ack => ptr_deref_2042_addr_3_req_0); -- 
    ra_9228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_3_ack_0, ack => cp_elements(584)); -- 
    cr_9229_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => ptr_deref_2042_addr_3_req_1); -- 
    ca_9230_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_addr_3_ack_1, ack => cp_elements(585)); -- 
    cpelement_group_586 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(576) & cp_elements(579) & cp_elements(582) & cp_elements(585));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(586),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(587) <= cp_elements(586);
    rr_9240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(587), ack => ptr_deref_2042_load_0_req_0); -- 
    ra_9241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_0_ack_0, ack => cp_elements(588)); -- 
    cp_elements(589) <= cp_elements(586);
    rr_9245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(589), ack => ptr_deref_2042_load_1_req_0); -- 
    ra_9246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_1_ack_0, ack => cp_elements(590)); -- 
    cp_elements(591) <= cp_elements(586);
    rr_9250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => ptr_deref_2042_load_2_req_0); -- 
    ra_9251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_2_ack_0, ack => cp_elements(592)); -- 
    cp_elements(593) <= cp_elements(586);
    rr_9255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_2042_load_3_req_0); -- 
    ra_9256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_3_ack_0, ack => cp_elements(594)); -- 
    cpelement_group_595 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(588) & cp_elements(590) & cp_elements(592) & cp_elements(594));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(595),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(596) <= cp_elements(595);
    cr_9266_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(596), ack => ptr_deref_2042_load_0_req_1); -- 
    ca_9267_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_0_ack_1, ack => cp_elements(597)); -- 
    cp_elements(598) <= cp_elements(595);
    cr_9271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(598), ack => ptr_deref_2042_load_1_req_1); -- 
    ca_9272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_1_ack_1, ack => cp_elements(599)); -- 
    cp_elements(600) <= cp_elements(595);
    cr_9276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => ptr_deref_2042_load_2_req_1); -- 
    ca_9277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_2_ack_1, ack => cp_elements(601)); -- 
    cp_elements(602) <= cp_elements(595);
    cr_9281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(602), ack => ptr_deref_2042_load_3_req_1); -- 
    ca_9282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_load_3_ack_1, ack => cp_elements(603)); -- 
    cpelement_group_604 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(597) & cp_elements(599) & cp_elements(601) & cp_elements(603));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(604),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9283_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(604), ack => ptr_deref_2042_gather_scatter_req_0); -- 
    merge_ack_9284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2042_gather_scatter_ack_0, ack => cp_elements(605)); -- 
    cp_elements(606) <= cp_elements(570);
    base_resize_req_9297_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(606), ack => ptr_deref_2046_base_resize_req_0); -- 
    base_resize_ack_9298_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_base_resize_ack_0, ack => cp_elements(607)); -- 
    sum_rename_req_9302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(607), ack => ptr_deref_2046_root_address_inst_req_0); -- 
    cp_elements(608) <= ptr_deref_2046_root_address_inst_ack_0;
    cp_elements(609) <= cp_elements(608);
    rr_9310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(609), ack => ptr_deref_2046_addr_0_req_0); -- 
    ra_9311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_0_ack_0, ack => cp_elements(610)); -- 
    cr_9312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(610), ack => ptr_deref_2046_addr_0_req_1); -- 
    ca_9313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_0_ack_1, ack => cp_elements(611)); -- 
    cp_elements(612) <= cp_elements(608);
    rr_9317_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(612), ack => ptr_deref_2046_addr_1_req_0); -- 
    ra_9318_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_1_ack_0, ack => cp_elements(613)); -- 
    cr_9319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => ptr_deref_2046_addr_1_req_1); -- 
    ca_9320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_1_ack_1, ack => cp_elements(614)); -- 
    cp_elements(615) <= cp_elements(608);
    rr_9324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(615), ack => ptr_deref_2046_addr_2_req_0); -- 
    ra_9325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_2_ack_0, ack => cp_elements(616)); -- 
    cr_9326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(616), ack => ptr_deref_2046_addr_2_req_1); -- 
    ca_9327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_2_ack_1, ack => cp_elements(617)); -- 
    cp_elements(618) <= cp_elements(608);
    rr_9331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(618), ack => ptr_deref_2046_addr_3_req_0); -- 
    ra_9332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_3_ack_0, ack => cp_elements(619)); -- 
    cr_9333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(619), ack => ptr_deref_2046_addr_3_req_1); -- 
    ca_9334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_addr_3_ack_1, ack => cp_elements(620)); -- 
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(611) & cp_elements(614) & cp_elements(617) & cp_elements(620));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(622) <= cp_elements(621);
    rr_9344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(622), ack => ptr_deref_2046_load_0_req_0); -- 
    ra_9345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_0_ack_0, ack => cp_elements(623)); -- 
    cp_elements(624) <= cp_elements(621);
    rr_9349_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(624), ack => ptr_deref_2046_load_1_req_0); -- 
    ra_9350_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_1_ack_0, ack => cp_elements(625)); -- 
    cp_elements(626) <= cp_elements(621);
    rr_9354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(626), ack => ptr_deref_2046_load_2_req_0); -- 
    ra_9355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_2_ack_0, ack => cp_elements(627)); -- 
    cp_elements(628) <= cp_elements(621);
    rr_9359_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(628), ack => ptr_deref_2046_load_3_req_0); -- 
    ra_9360_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_3_ack_0, ack => cp_elements(629)); -- 
    cpelement_group_630 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(623) & cp_elements(625) & cp_elements(627) & cp_elements(629));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(630),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(631) <= cp_elements(630);
    cr_9370_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(631), ack => ptr_deref_2046_load_0_req_1); -- 
    ca_9371_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_0_ack_1, ack => cp_elements(632)); -- 
    cp_elements(633) <= cp_elements(630);
    cr_9375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(633), ack => ptr_deref_2046_load_1_req_1); -- 
    ca_9376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_1_ack_1, ack => cp_elements(634)); -- 
    cp_elements(635) <= cp_elements(630);
    cr_9380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(635), ack => ptr_deref_2046_load_2_req_1); -- 
    ca_9381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_2_ack_1, ack => cp_elements(636)); -- 
    cp_elements(637) <= cp_elements(630);
    cr_9385_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(637), ack => ptr_deref_2046_load_3_req_1); -- 
    ca_9386_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_load_3_ack_1, ack => cp_elements(638)); -- 
    cpelement_group_639 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(632) & cp_elements(634) & cp_elements(636) & cp_elements(638));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(639),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(639), ack => ptr_deref_2046_gather_scatter_req_0); -- 
    merge_ack_9388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2046_gather_scatter_ack_0, ack => cp_elements(640)); -- 
    cpelement_group_641 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(605) & cp_elements(640) & cp_elements(642));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(641),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(641), ack => binary_2051_inst_req_0); -- 
    cp_elements(642) <= cp_elements(570);
    ra_9399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2051_inst_ack_0, ack => cp_elements(643)); -- 
    cr_9400_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => binary_2051_inst_req_1); -- 
    ca_9401_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2051_inst_ack_1, ack => cp_elements(644)); -- 
    cp_elements(645) <= cp_elements(644);
    cp_elements(646) <= false;
    cp_elements(647) <= cp_elements(646);
    cp_elements(648) <= cp_elements(644);
    branch_req_9409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(648), ack => if_stmt_2053_branch_req_0); -- 
    cp_elements(649) <= cp_elements(648);
    cp_elements(650) <= cp_elements(649);
    if_choice_transition_9414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2053_branch_ack_1, ack => cp_elements(651)); -- 
    cp_elements(652) <= cp_elements(649);
    else_choice_transition_9418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2053_branch_ack_0, ack => cp_elements(653)); -- 
    base_resize_ack_9437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_base_resize_ack_0, ack => cp_elements(654)); -- 
    sum_rename_req_9441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_2062_root_address_inst_req_0); -- 
    cp_elements(655) <= ptr_deref_2062_root_address_inst_ack_0;
    cp_elements(656) <= cp_elements(655);
    rr_9449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => ptr_deref_2062_addr_0_req_0); -- 
    ra_9450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_0_ack_0, ack => cp_elements(657)); -- 
    cr_9451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(657), ack => ptr_deref_2062_addr_0_req_1); -- 
    ca_9452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_0_ack_1, ack => cp_elements(658)); -- 
    cp_elements(659) <= cp_elements(655);
    rr_9456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(659), ack => ptr_deref_2062_addr_1_req_0); -- 
    ra_9457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_1_ack_0, ack => cp_elements(660)); -- 
    cr_9458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(660), ack => ptr_deref_2062_addr_1_req_1); -- 
    ca_9459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_1_ack_1, ack => cp_elements(661)); -- 
    cp_elements(662) <= cp_elements(655);
    rr_9463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(662), ack => ptr_deref_2062_addr_2_req_0); -- 
    ra_9464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_2_ack_0, ack => cp_elements(663)); -- 
    cr_9465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(663), ack => ptr_deref_2062_addr_2_req_1); -- 
    ca_9466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_2_ack_1, ack => cp_elements(664)); -- 
    cp_elements(665) <= cp_elements(655);
    rr_9470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(665), ack => ptr_deref_2062_addr_3_req_0); -- 
    ra_9471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_3_ack_0, ack => cp_elements(666)); -- 
    cr_9472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(666), ack => ptr_deref_2062_addr_3_req_1); -- 
    ca_9473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_addr_3_ack_1, ack => cp_elements(667)); -- 
    cpelement_group_668 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(658) & cp_elements(661) & cp_elements(664) & cp_elements(667));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(668),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(669) <= cp_elements(668);
    rr_9483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(669), ack => ptr_deref_2062_load_0_req_0); -- 
    ra_9484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_0_ack_0, ack => cp_elements(670)); -- 
    cp_elements(671) <= cp_elements(668);
    rr_9488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(671), ack => ptr_deref_2062_load_1_req_0); -- 
    ra_9489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_1_ack_0, ack => cp_elements(672)); -- 
    cp_elements(673) <= cp_elements(668);
    rr_9493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(673), ack => ptr_deref_2062_load_2_req_0); -- 
    ra_9494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_2_ack_0, ack => cp_elements(674)); -- 
    cp_elements(675) <= cp_elements(668);
    rr_9498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(675), ack => ptr_deref_2062_load_3_req_0); -- 
    ra_9499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_3_ack_0, ack => cp_elements(676)); -- 
    cpelement_group_677 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(670) & cp_elements(672) & cp_elements(674) & cp_elements(676));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(677),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(678) <= cp_elements(677);
    cr_9509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(678), ack => ptr_deref_2062_load_0_req_1); -- 
    ca_9510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_0_ack_1, ack => cp_elements(679)); -- 
    cp_elements(680) <= cp_elements(677);
    cr_9514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(680), ack => ptr_deref_2062_load_1_req_1); -- 
    ca_9515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_1_ack_1, ack => cp_elements(681)); -- 
    cp_elements(682) <= cp_elements(677);
    cr_9519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(682), ack => ptr_deref_2062_load_2_req_1); -- 
    ca_9520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_2_ack_1, ack => cp_elements(683)); -- 
    cp_elements(684) <= cp_elements(677);
    cr_9524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(684), ack => ptr_deref_2062_load_3_req_1); -- 
    ca_9525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_load_3_ack_1, ack => cp_elements(685)); -- 
    cpelement_group_686 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(679) & cp_elements(681) & cp_elements(683) & cp_elements(685));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(686),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_9526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => ptr_deref_2062_gather_scatter_req_0); -- 
    merge_ack_9527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2062_gather_scatter_ack_0, ack => cp_elements(687)); -- 
    cp_elements(688) <= cp_elements(1007);
    cp_elements(689) <= cp_elements(688);
    cpelement_group_690 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(689) & cp_elements(691) & cp_elements(695));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(690),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_9558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(690), ack => ptr_deref_2067_gather_scatter_req_0); -- 
    cp_elements(691) <= cp_elements(688);
    cp_elements(692) <= cp_elements(691);
    base_resize_req_9543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(692), ack => ptr_deref_2067_base_resize_req_0); -- 
    base_resize_ack_9544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_base_resize_ack_0, ack => cp_elements(693)); -- 
    sum_rename_req_9548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => ptr_deref_2067_root_address_inst_req_0); -- 
    sum_rename_ack_9549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_root_address_inst_ack_0, ack => cp_elements(694)); -- 
    root_rename_req_9553_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(694), ack => ptr_deref_2067_addr_0_req_0); -- 
    root_rename_ack_9554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_addr_0_ack_0, ack => cp_elements(695)); -- 
    split_ack_9559_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_gather_scatter_ack_0, ack => cp_elements(696)); -- 
    rr_9566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(696), ack => ptr_deref_2067_store_0_req_0); -- 
    ra_9567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_store_0_ack_0, ack => cp_elements(697)); -- 
    cr_9577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => ptr_deref_2067_store_0_req_1); -- 
    ca_9578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2067_store_0_ack_1, ack => cp_elements(698)); -- 
    cpelement_group_699 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(700) & cp_elements(701));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(699),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => binary_2077_inst_req_0); -- 
    cp_elements(700) <= cp_elements(1009);
    cp_elements(701) <= cp_elements(1009);
    ra_9594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2077_inst_ack_0, ack => cp_elements(702)); -- 
    cr_9595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => binary_2077_inst_req_1); -- 
    ca_9596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2077_inst_ack_1, ack => cp_elements(703)); -- 
    pipe_wreq_9601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(703), ack => simple_obj_ref_2074_inst_req_0); -- 
    pipe_wack_9602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2074_inst_ack_0, ack => cp_elements(704)); -- 
    cp_elements(705) <= cp_elements(174);
    cpelement_group_706 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(707) & cp_elements(715));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(706),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(706), ack => addr_of_2087_final_reg_req_0); -- 
    cp_elements(707) <= cp_elements(705);
    cp_elements(708) <= cp_elements(705);
    index_resize_req_9619_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(708), ack => array_obj_ref_2086_index_0_resize_req_0); -- 
    index_resize_ack_9620_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_index_0_resize_ack_0, ack => cp_elements(709)); -- 
    scale_rr_9624_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(709), ack => array_obj_ref_2086_index_0_scale_req_0); -- 
    scale_ra_9625_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_index_0_scale_ack_0, ack => cp_elements(710)); -- 
    scale_cr_9626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(710), ack => array_obj_ref_2086_index_0_scale_req_1); -- 
    scale_ca_9627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_index_0_scale_ack_1, ack => cp_elements(711)); -- 
    partial_sum_1_rr_9631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => array_obj_ref_2086_index_sum_1_req_0); -- 
    partial_sum_1_ra_9632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_index_sum_1_ack_0, ack => cp_elements(712)); -- 
    partial_sum_1_cr_9633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(712), ack => array_obj_ref_2086_index_sum_1_req_1); -- 
    partial_sum_1_ca_9634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_index_sum_1_ack_1, ack => cp_elements(713)); -- 
    final_index_req_9635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(713), ack => array_obj_ref_2086_offset_inst_req_0); -- 
    final_index_ack_9636_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_offset_inst_ack_0, ack => cp_elements(714)); -- 
    sum_rename_req_9640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(714), ack => array_obj_ref_2086_root_address_inst_req_0); -- 
    sum_rename_ack_9641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2086_root_address_inst_ack_0, ack => cp_elements(715)); -- 
    final_reg_ack_9646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2087_final_reg_ack_0, ack => cp_elements(716)); -- 
    base_resize_req_9659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(716), ack => ptr_deref_2091_base_resize_req_0); -- 
    base_resize_ack_9660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_base_resize_ack_0, ack => cp_elements(717)); -- 
    sum_rename_req_9664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(717), ack => ptr_deref_2091_root_address_inst_req_0); -- 
    sum_rename_ack_9665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_root_address_inst_ack_0, ack => cp_elements(718)); -- 
    root_rename_req_9669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(718), ack => ptr_deref_2091_addr_0_req_0); -- 
    root_rename_ack_9670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_addr_0_ack_0, ack => cp_elements(719)); -- 
    rr_9680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(719), ack => ptr_deref_2091_load_0_req_0); -- 
    ra_9681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_load_0_ack_0, ack => cp_elements(720)); -- 
    cr_9691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => ptr_deref_2091_load_0_req_1); -- 
    ca_9692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_load_0_ack_1, ack => cp_elements(721)); -- 
    merge_req_9693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(721), ack => ptr_deref_2091_gather_scatter_req_0); -- 
    merge_ack_9694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2091_gather_scatter_ack_0, ack => cp_elements(722)); -- 
    cpelement_group_723 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(722) & cp_elements(724));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(723),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(723), ack => binary_2097_inst_req_0); -- 
    cp_elements(724) <= cp_elements(705);
    ra_9704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2097_inst_ack_0, ack => cp_elements(725)); -- 
    cr_9705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(725), ack => binary_2097_inst_req_1); -- 
    ca_9706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2097_inst_ack_1, ack => cp_elements(726)); -- 
    index_resize_req_9720_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(726), ack => array_obj_ref_2105_index_2_resize_req_0); -- 
    cpelement_group_727 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(728) & cp_elements(734));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(727),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(727), ack => addr_of_2106_final_reg_req_0); -- 
    cp_elements(728) <= cp_elements(705);
    index_resize_ack_9721_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_index_2_resize_ack_0, ack => cp_elements(729)); -- 
    scale_rename_req_9725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => array_obj_ref_2105_index_2_rename_req_0); -- 
    scale_rename_ack_9726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_index_2_rename_ack_0, ack => cp_elements(730)); -- 
    partial_sum_1_rr_9730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(730), ack => array_obj_ref_2105_index_sum_1_req_0); -- 
    partial_sum_1_ra_9731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_index_sum_1_ack_0, ack => cp_elements(731)); -- 
    partial_sum_1_cr_9732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(731), ack => array_obj_ref_2105_index_sum_1_req_1); -- 
    partial_sum_1_ca_9733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_index_sum_1_ack_1, ack => cp_elements(732)); -- 
    final_index_req_9734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(732), ack => array_obj_ref_2105_offset_inst_req_0); -- 
    final_index_ack_9735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_offset_inst_ack_0, ack => cp_elements(733)); -- 
    sum_rename_req_9739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(733), ack => array_obj_ref_2105_root_address_inst_req_0); -- 
    sum_rename_ack_9740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2105_root_address_inst_ack_0, ack => cp_elements(734)); -- 
    final_reg_ack_9745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2106_final_reg_ack_0, ack => cp_elements(735)); -- 
    base_resize_req_9758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(735), ack => ptr_deref_2110_base_resize_req_0); -- 
    base_resize_ack_9759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_base_resize_ack_0, ack => cp_elements(736)); -- 
    sum_rename_req_9763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => ptr_deref_2110_root_address_inst_req_0); -- 
    sum_rename_ack_9764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_root_address_inst_ack_0, ack => cp_elements(737)); -- 
    root_rename_req_9768_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(737), ack => ptr_deref_2110_addr_0_req_0); -- 
    root_rename_ack_9769_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_addr_0_ack_0, ack => cp_elements(738)); -- 
    rr_9779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(738), ack => ptr_deref_2110_load_0_req_0); -- 
    ra_9780_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_load_0_ack_0, ack => cp_elements(739)); -- 
    cr_9790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(739), ack => ptr_deref_2110_load_0_req_1); -- 
    ca_9791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_load_0_ack_1, ack => cp_elements(740)); -- 
    merge_req_9792_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => ptr_deref_2110_gather_scatter_req_0); -- 
    merge_ack_9793_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2110_gather_scatter_ack_0, ack => cp_elements(741)); -- 
    cpelement_group_742 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(741) & cp_elements(743));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(742),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => binary_2116_inst_req_0); -- 
    cp_elements(743) <= cp_elements(705);
    ra_9803_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2116_inst_ack_0, ack => cp_elements(744)); -- 
    cr_9804_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => binary_2116_inst_req_1); -- 
    ca_9805_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2116_inst_ack_1, ack => cp_elements(745)); -- 
    cp_elements(746) <= cp_elements(745);
    cp_elements(747) <= false;
    cp_elements(748) <= cp_elements(747);
    cp_elements(749) <= cp_elements(745);
    branch_req_9813_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(749), ack => if_stmt_2118_branch_req_0); -- 
    cp_elements(750) <= cp_elements(749);
    cp_elements(751) <= cp_elements(750);
    if_choice_transition_9818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2118_branch_ack_1, ack => cp_elements(752)); -- 
    cp_elements(753) <= cp_elements(750);
    else_choice_transition_9822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2118_branch_ack_0, ack => cp_elements(754)); -- 
    cp_elements(755) <= cp_elements(15);
    cpelement_group_756 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(757) & cp_elements(758));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(756),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9836_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => binary_2129_inst_req_0); -- 
    cp_elements(757) <= cp_elements(755);
    cp_elements(758) <= cp_elements(755);
    ra_9837_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2129_inst_ack_0, ack => cp_elements(759)); -- 
    cr_9838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(759), ack => binary_2129_inst_req_1); -- 
    ca_9839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2129_inst_ack_1, ack => cp_elements(760)); -- 
    index_resize_req_9853_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(760), ack => array_obj_ref_2137_index_2_resize_req_0); -- 
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(762) & cp_elements(768));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_9877_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(761), ack => addr_of_2138_final_reg_req_0); -- 
    cp_elements(762) <= cp_elements(755);
    index_resize_ack_9854_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_index_2_resize_ack_0, ack => cp_elements(763)); -- 
    scale_rename_req_9858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => array_obj_ref_2137_index_2_rename_req_0); -- 
    scale_rename_ack_9859_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_index_2_rename_ack_0, ack => cp_elements(764)); -- 
    partial_sum_1_rr_9863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(764), ack => array_obj_ref_2137_index_sum_1_req_0); -- 
    partial_sum_1_ra_9864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_index_sum_1_ack_0, ack => cp_elements(765)); -- 
    partial_sum_1_cr_9865_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => array_obj_ref_2137_index_sum_1_req_1); -- 
    partial_sum_1_ca_9866_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_index_sum_1_ack_1, ack => cp_elements(766)); -- 
    final_index_req_9867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(766), ack => array_obj_ref_2137_offset_inst_req_0); -- 
    final_index_ack_9868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_offset_inst_ack_0, ack => cp_elements(767)); -- 
    sum_rename_req_9872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => array_obj_ref_2137_root_address_inst_req_0); -- 
    sum_rename_ack_9873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2137_root_address_inst_ack_0, ack => cp_elements(768)); -- 
    final_reg_ack_9878_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2138_final_reg_ack_0, ack => cp_elements(769)); -- 
    base_resize_req_9891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(769), ack => ptr_deref_2142_base_resize_req_0); -- 
    base_resize_ack_9892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_base_resize_ack_0, ack => cp_elements(770)); -- 
    sum_rename_req_9896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(770), ack => ptr_deref_2142_root_address_inst_req_0); -- 
    sum_rename_ack_9897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_root_address_inst_ack_0, ack => cp_elements(771)); -- 
    root_rename_req_9901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(771), ack => ptr_deref_2142_addr_0_req_0); -- 
    root_rename_ack_9902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_addr_0_ack_0, ack => cp_elements(772)); -- 
    rr_9912_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => ptr_deref_2142_load_0_req_0); -- 
    ra_9913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_load_0_ack_0, ack => cp_elements(773)); -- 
    cr_9923_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(773), ack => ptr_deref_2142_load_0_req_1); -- 
    ca_9924_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_load_0_ack_1, ack => cp_elements(774)); -- 
    merge_req_9925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(774), ack => ptr_deref_2142_gather_scatter_req_0); -- 
    merge_ack_9926_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2142_gather_scatter_ack_0, ack => cp_elements(775)); -- 
    cpelement_group_776 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(775) & cp_elements(777));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(776),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(776), ack => binary_2148_inst_req_0); -- 
    cp_elements(777) <= cp_elements(755);
    ra_9936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2148_inst_ack_0, ack => cp_elements(778)); -- 
    cr_9937_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(778), ack => binary_2148_inst_req_1); -- 
    ca_9938_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2148_inst_ack_1, ack => cp_elements(779)); -- 
    cp_elements(780) <= cp_elements(779);
    cp_elements(781) <= false;
    cp_elements(782) <= cp_elements(781);
    cp_elements(783) <= cp_elements(779);
    branch_req_9946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => if_stmt_2150_branch_req_0); -- 
    cp_elements(784) <= cp_elements(783);
    cp_elements(785) <= cp_elements(784);
    if_choice_transition_9951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2150_branch_ack_1, ack => cp_elements(786)); -- 
    cp_elements(787) <= cp_elements(784);
    else_choice_transition_9955_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2150_branch_ack_0, ack => cp_elements(788)); -- 
    cp_elements(789) <= cp_elements(16);
    cpelement_group_790 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(791) & cp_elements(792));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(790),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_9969_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(790), ack => binary_2161_inst_req_0); -- 
    cp_elements(791) <= cp_elements(789);
    cp_elements(792) <= cp_elements(789);
    ra_9970_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2161_inst_ack_0, ack => cp_elements(793)); -- 
    cr_9971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(793), ack => binary_2161_inst_req_1); -- 
    ca_9972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2161_inst_ack_1, ack => cp_elements(794)); -- 
    index_resize_req_9986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(794), ack => array_obj_ref_2169_index_2_resize_req_0); -- 
    cpelement_group_795 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(796) & cp_elements(802));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(795),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_10010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(795), ack => addr_of_2170_final_reg_req_0); -- 
    cp_elements(796) <= cp_elements(789);
    index_resize_ack_9987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_index_2_resize_ack_0, ack => cp_elements(797)); -- 
    scale_rename_req_9991_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => array_obj_ref_2169_index_2_rename_req_0); -- 
    scale_rename_ack_9992_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_index_2_rename_ack_0, ack => cp_elements(798)); -- 
    partial_sum_1_rr_9996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(798), ack => array_obj_ref_2169_index_sum_1_req_0); -- 
    partial_sum_1_ra_9997_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_index_sum_1_ack_0, ack => cp_elements(799)); -- 
    partial_sum_1_cr_9998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => array_obj_ref_2169_index_sum_1_req_1); -- 
    partial_sum_1_ca_9999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_index_sum_1_ack_1, ack => cp_elements(800)); -- 
    final_index_req_10000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(800), ack => array_obj_ref_2169_offset_inst_req_0); -- 
    final_index_ack_10001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_offset_inst_ack_0, ack => cp_elements(801)); -- 
    sum_rename_req_10005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(801), ack => array_obj_ref_2169_root_address_inst_req_0); -- 
    sum_rename_ack_10006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2169_root_address_inst_ack_0, ack => cp_elements(802)); -- 
    final_reg_ack_10011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_2170_final_reg_ack_0, ack => cp_elements(803)); -- 
    base_resize_req_10024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(803), ack => ptr_deref_2174_base_resize_req_0); -- 
    base_resize_ack_10025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_base_resize_ack_0, ack => cp_elements(804)); -- 
    sum_rename_req_10029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(804), ack => ptr_deref_2174_root_address_inst_req_0); -- 
    sum_rename_ack_10030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_root_address_inst_ack_0, ack => cp_elements(805)); -- 
    root_rename_req_10034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(805), ack => ptr_deref_2174_addr_0_req_0); -- 
    root_rename_ack_10035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_addr_0_ack_0, ack => cp_elements(806)); -- 
    rr_10045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_2174_load_0_req_0); -- 
    ra_10046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_load_0_ack_0, ack => cp_elements(807)); -- 
    cr_10056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(807), ack => ptr_deref_2174_load_0_req_1); -- 
    ca_10057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_load_0_ack_1, ack => cp_elements(808)); -- 
    merge_req_10058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => ptr_deref_2174_gather_scatter_req_0); -- 
    merge_ack_10059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2174_gather_scatter_ack_0, ack => cp_elements(809)); -- 
    cpelement_group_810 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(811) & cp_elements(814));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(810),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => binary_2183_inst_req_0); -- 
    cp_elements(811) <= cp_elements(789);
    cpelement_group_812 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(809) & cp_elements(813));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(812),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => type_cast_2179_inst_req_0); -- 
    cp_elements(813) <= cp_elements(789);
    ack_10071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2179_inst_ack_0, ack => cp_elements(814)); -- 
    ra_10076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2183_inst_ack_0, ack => cp_elements(815)); -- 
    cr_10077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => binary_2183_inst_req_1); -- 
    ca_10078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2183_inst_ack_1, ack => cp_elements(816)); -- 
    cp_elements(817) <= cp_elements(816);
    cp_elements(818) <= false;
    cp_elements(819) <= cp_elements(818);
    cp_elements(820) <= cp_elements(816);
    branch_req_10086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(820), ack => if_stmt_2185_branch_req_0); -- 
    cp_elements(821) <= cp_elements(820);
    cp_elements(822) <= cp_elements(821);
    if_choice_transition_10091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2185_branch_ack_1, ack => cp_elements(823)); -- 
    cp_elements(824) <= cp_elements(821);
    else_choice_transition_10095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2185_branch_ack_0, ack => cp_elements(825)); -- 
    cp_elements(826) <= cp_elements(17);
    cpelement_group_827 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(828) & cp_elements(832));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(827),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(827), ack => binary_2198_inst_req_0); -- 
    cp_elements(828) <= cp_elements(826);
    cpelement_group_829 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(830) & cp_elements(831));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(829),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(829), ack => type_cast_2194_inst_req_0); -- 
    cp_elements(830) <= cp_elements(826);
    cp_elements(831) <= cp_elements(826);
    ack_10112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2194_inst_ack_0, ack => cp_elements(832)); -- 
    ra_10117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2198_inst_ack_0, ack => cp_elements(833)); -- 
    cr_10118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(833), ack => binary_2198_inst_req_1); -- 
    ca_10119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2198_inst_ack_1, ack => cp_elements(834)); -- 
    cp_elements(835) <= cp_elements(834);
    cp_elements(836) <= false;
    cp_elements(837) <= cp_elements(836);
    cp_elements(838) <= cp_elements(834);
    branch_req_10127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(838), ack => if_stmt_2200_branch_req_0); -- 
    cp_elements(839) <= cp_elements(838);
    cp_elements(840) <= cp_elements(839);
    if_choice_transition_10132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2200_branch_ack_1, ack => cp_elements(841)); -- 
    cp_elements(842) <= cp_elements(839);
    else_choice_transition_10136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2200_branch_ack_0, ack => cp_elements(843)); -- 
    cp_elements(844) <= cp_elements(18);
    cpelement_group_845 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(846) & cp_elements(847));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(845),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(845), ack => binary_2211_inst_req_0); -- 
    cp_elements(846) <= cp_elements(844);
    cp_elements(847) <= cp_elements(844);
    ra_10151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2211_inst_ack_0, ack => cp_elements(848)); -- 
    cr_10152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(848), ack => binary_2211_inst_req_1); -- 
    ca_10153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2211_inst_ack_1, ack => cp_elements(849)); -- 
    cp_elements(850) <= cp_elements(849);
    cp_elements(851) <= false;
    cp_elements(852) <= cp_elements(851);
    cp_elements(853) <= cp_elements(849);
    branch_req_10161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => if_stmt_2213_branch_req_0); -- 
    cp_elements(854) <= cp_elements(853);
    cp_elements(855) <= cp_elements(854);
    if_choice_transition_10166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2213_branch_ack_1, ack => cp_elements(856)); -- 
    cp_elements(857) <= cp_elements(854);
    else_choice_transition_10170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2213_branch_ack_0, ack => cp_elements(858)); -- 
    cp_elements(859) <= cp_elements(19);
    cpelement_group_860 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(861) & cp_elements(862));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(860),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(860), ack => binary_2224_inst_req_0); -- 
    cp_elements(861) <= cp_elements(859);
    cp_elements(862) <= cp_elements(859);
    ra_10185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2224_inst_ack_0, ack => cp_elements(863)); -- 
    cr_10186_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(863), ack => binary_2224_inst_req_1); -- 
    ca_10187_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2224_inst_ack_1, ack => cp_elements(864)); -- 
    cp_elements(865) <= cp_elements(864);
    cp_elements(866) <= false;
    cp_elements(867) <= cp_elements(866);
    cp_elements(868) <= cp_elements(864);
    branch_req_10195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(868), ack => if_stmt_2226_branch_req_0); -- 
    cp_elements(869) <= cp_elements(868);
    cp_elements(870) <= cp_elements(869);
    if_choice_transition_10200_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2226_branch_ack_1, ack => cp_elements(871)); -- 
    cp_elements(872) <= cp_elements(869);
    else_choice_transition_10204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2226_branch_ack_0, ack => cp_elements(873)); -- 
    cp_elements(874) <= cp_elements(20);
    cpelement_group_875 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(876) & cp_elements(880));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(875),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(875), ack => binary_2239_inst_req_0); -- 
    cp_elements(876) <= cp_elements(874);
    cpelement_group_877 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(878) & cp_elements(879));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(877),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(877), ack => type_cast_2235_inst_req_0); -- 
    cp_elements(878) <= cp_elements(874);
    cp_elements(879) <= cp_elements(874);
    ack_10221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2235_inst_ack_0, ack => cp_elements(880)); -- 
    ra_10226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2239_inst_ack_0, ack => cp_elements(881)); -- 
    cr_10227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(881), ack => binary_2239_inst_req_1); -- 
    ca_10228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2239_inst_ack_1, ack => cp_elements(882)); -- 
    cp_elements(883) <= cp_elements(882);
    cp_elements(884) <= false;
    cp_elements(885) <= cp_elements(884);
    cp_elements(886) <= cp_elements(882);
    branch_req_10236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(886), ack => if_stmt_2241_branch_req_0); -- 
    cp_elements(887) <= cp_elements(886);
    cp_elements(888) <= cp_elements(887);
    if_choice_transition_10241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2241_branch_ack_1, ack => cp_elements(889)); -- 
    cp_elements(890) <= cp_elements(887);
    else_choice_transition_10245_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2241_branch_ack_0, ack => cp_elements(891)); -- 
    cp_elements(892) <= cp_elements(21);
    cpelement_group_893 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(894) & cp_elements(895));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(893),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(893), ack => binary_2252_inst_req_0); -- 
    cp_elements(894) <= cp_elements(892);
    cp_elements(895) <= cp_elements(892);
    ra_10260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2252_inst_ack_0, ack => cp_elements(896)); -- 
    cr_10261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(896), ack => binary_2252_inst_req_1); -- 
    ca_10262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2252_inst_ack_1, ack => cp_elements(897)); -- 
    cp_elements(898) <= cp_elements(897);
    cp_elements(899) <= false;
    cp_elements(900) <= cp_elements(899);
    cp_elements(901) <= cp_elements(897);
    branch_req_10270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(901), ack => if_stmt_2254_branch_req_0); -- 
    cp_elements(902) <= cp_elements(901);
    cp_elements(903) <= cp_elements(902);
    if_choice_transition_10275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2254_branch_ack_1, ack => cp_elements(904)); -- 
    cp_elements(905) <= cp_elements(902);
    else_choice_transition_10279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2254_branch_ack_0, ack => cp_elements(906)); -- 
    cp_elements(907) <= cp_elements(22);
    cpelement_group_908 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(909) & cp_elements(910));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(908),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10293_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(908), ack => binary_2265_inst_req_0); -- 
    cp_elements(909) <= cp_elements(907);
    cp_elements(910) <= cp_elements(907);
    ra_10294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2265_inst_ack_0, ack => cp_elements(911)); -- 
    cr_10295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(911), ack => binary_2265_inst_req_1); -- 
    ca_10296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2265_inst_ack_1, ack => cp_elements(912)); -- 
    cp_elements(913) <= cp_elements(912);
    cp_elements(914) <= false;
    cp_elements(915) <= cp_elements(914);
    cp_elements(916) <= cp_elements(912);
    branch_req_10304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(916), ack => if_stmt_2267_branch_req_0); -- 
    cp_elements(917) <= cp_elements(916);
    cp_elements(918) <= cp_elements(917);
    if_choice_transition_10309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2267_branch_ack_1, ack => cp_elements(919)); -- 
    cp_elements(920) <= cp_elements(917);
    else_choice_transition_10313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_2267_branch_ack_0, ack => cp_elements(921)); -- 
    cp_elements(922) <= cp_elements(23);
    cpelement_group_923 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(924) & cp_elements(925));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(923),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(923), ack => type_cast_2276_inst_req_0); -- 
    cp_elements(924) <= cp_elements(922);
    cp_elements(925) <= cp_elements(922);
    ack_10328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2276_inst_ack_0, ack => cp_elements(926)); -- 
    pipe_wreq_10333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(926), ack => simple_obj_ref_2274_inst_req_0); -- 
    pipe_wack_10334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2274_inst_ack_0, ack => cp_elements(927)); -- 
    cp_elements(928) <= cp_elements(904);
    cpelement_group_929 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(930) & cp_elements(931));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(929),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => type_cast_2282_inst_req_0); -- 
    cp_elements(930) <= cp_elements(928);
    cp_elements(931) <= cp_elements(928);
    ack_10347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2282_inst_ack_0, ack => cp_elements(932)); -- 
    pipe_wreq_10352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => simple_obj_ref_2280_inst_req_0); -- 
    pipe_wack_10353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2280_inst_ack_0, ack => cp_elements(933)); -- 
    cp_elements(934) <= cp_elements(871);
    cpelement_group_935 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(936) & cp_elements(937));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(935),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(935), ack => type_cast_2288_inst_req_0); -- 
    cp_elements(936) <= cp_elements(934);
    cp_elements(937) <= cp_elements(934);
    ack_10366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2288_inst_ack_0, ack => cp_elements(938)); -- 
    pipe_wreq_10371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(938), ack => simple_obj_ref_2286_inst_req_0); -- 
    pipe_wack_10372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2286_inst_ack_0, ack => cp_elements(939)); -- 
    cp_elements(940) <= cp_elements(856);
    cpelement_group_941 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(942) & cp_elements(943));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(941),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(941), ack => type_cast_2294_inst_req_0); -- 
    cp_elements(942) <= cp_elements(940);
    cp_elements(943) <= cp_elements(940);
    ack_10385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2294_inst_ack_0, ack => cp_elements(944)); -- 
    pipe_wreq_10390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => simple_obj_ref_2292_inst_req_0); -- 
    pipe_wack_10391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2292_inst_ack_0, ack => cp_elements(945)); -- 
    cp_elements(946) <= cp_elements(1029);
    cpelement_group_947 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(948) & cp_elements(949));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(947),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(947), ack => type_cast_2300_inst_req_0); -- 
    cp_elements(948) <= cp_elements(946);
    cp_elements(949) <= cp_elements(946);
    ack_10404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2300_inst_ack_0, ack => cp_elements(950)); -- 
    pipe_wreq_10409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(950), ack => simple_obj_ref_2298_inst_req_0); -- 
    pipe_wack_10410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2298_inst_ack_0, ack => cp_elements(951)); -- 
    cp_elements(952) <= false;
    cp_elements(953) <= cp_elements(952);
    ack_10459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1781_inst_ack_0, ack => cp_elements(954)); -- 
    phi_stmt_1778_req_10460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(954), ack => phi_stmt_1778_req_0); -- 
    cp_elements(955) <= OrReduce(cp_elements(77) & cp_elements(954));
    cp_elements(956) <= cp_elements(955);
    phi_stmt_1778_ack_10465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1778_ack_0, ack => cp_elements(957)); -- 
    cp_elements(958) <= false;
    cp_elements(959) <= cp_elements(958);
    cp_elements(960) <= false;
    cp_elements(961) <= cp_elements(960);
    cp_elements(962) <= OrReduce(cp_elements(158) & cp_elements(176));
    cp_elements(963) <= cp_elements(962);
    cp_elements(964) <= false;
    cp_elements(965) <= cp_elements(964);
    cp_elements(966) <= cp_elements(5);
    cp_elements(967) <= cp_elements(966);
    phi_stmt_1845_req_10519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(967), ack => phi_stmt_1845_req_1); -- 
    cp_elements(968) <= cp_elements(966);
    phi_stmt_1852_req_10531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(968), ack => phi_stmt_1852_req_1); -- 
    cpelement_group_969 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(967) & cp_elements(968));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(969),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(970) <= cp_elements(271);
    cp_elements(971) <= cp_elements(970);
    req_10544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(971), ack => type_cast_1848_inst_req_0); -- 
    ack_10545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1848_inst_ack_0, ack => cp_elements(972)); -- 
    phi_stmt_1845_req_10546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(972), ack => phi_stmt_1845_req_0); -- 
    cp_elements(973) <= cp_elements(970);
    req_10556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(973), ack => type_cast_1855_inst_req_0); -- 
    ack_10557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1855_inst_ack_0, ack => cp_elements(974)); -- 
    phi_stmt_1852_req_10558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(974), ack => phi_stmt_1852_req_0); -- 
    cpelement_group_975 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(972) & cp_elements(974));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(975),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(976) <= OrReduce(cp_elements(969) & cp_elements(975));
    cp_elements(977) <= cp_elements(976);
    phi_stmt_1845_ack_10563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1845_ack_0, ack => cp_elements(978)); -- 
    phi_stmt_1852_ack_10564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1852_ack_0, ack => cp_elements(979)); -- 
    cpelement_group_980 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(978) & cp_elements(979));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(980),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(981) <= false;
    cp_elements(982) <= cp_elements(981);
    cp_elements(983) <= cp_elements(240);
    cp_elements(984) <= cp_elements(240);
    req_10594_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(984), ack => type_cast_1898_inst_req_0); -- 
    ack_10595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1898_inst_ack_0, ack => cp_elements(985)); -- 
    cpelement_group_986 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(983) & cp_elements(985));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(986),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1893_req_10596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(986), ack => phi_stmt_1893_req_1); -- 
    cp_elements(987) <= cp_elements(252);
    req_10609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(987), ack => type_cast_1896_inst_req_0); -- 
    ack_10610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1896_inst_ack_0, ack => cp_elements(988)); -- 
    cp_elements(989) <= cp_elements(252);
    cpelement_group_990 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(988) & cp_elements(989));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(990),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    phi_stmt_1893_req_10616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(990), ack => phi_stmt_1893_req_0); -- 
    cp_elements(991) <= OrReduce(cp_elements(986) & cp_elements(990));
    cp_elements(992) <= cp_elements(991);
    phi_stmt_1893_ack_10621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1893_ack_0, ack => cp_elements(993)); -- 
    cp_elements(994) <= false;
    cp_elements(995) <= cp_elements(994);
    cp_elements(996) <= false;
    cp_elements(997) <= cp_elements(996);
    cp_elements(998) <= false;
    cp_elements(999) <= cp_elements(998);
    cp_elements(1000) <= OrReduce(cp_elements(427) & cp_elements(440));
    cp_elements(1001) <= cp_elements(1000);
    cp_elements(1002) <= false;
    cp_elements(1003) <= cp_elements(1002);
    cp_elements(1004) <= false;
    cp_elements(1005) <= cp_elements(1004);
    cp_elements(1006) <= OrReduce(cp_elements(653) & cp_elements(687));
    cp_elements(1007) <= cp_elements(1006);
    cp_elements(1008) <= OrReduce(cp_elements(9) & cp_elements(209) & cp_elements(569) & cp_elements(698));
    cp_elements(1009) <= cp_elements(1008);
    cp_elements(1010) <= false;
    cp_elements(1011) <= cp_elements(1010);
    cp_elements(1012) <= false;
    cp_elements(1013) <= cp_elements(1012);
    cp_elements(1014) <= false;
    cp_elements(1015) <= cp_elements(1014);
    cp_elements(1016) <= false;
    cp_elements(1017) <= cp_elements(1016);
    cp_elements(1018) <= false;
    cp_elements(1019) <= cp_elements(1018);
    cp_elements(1020) <= false;
    cp_elements(1021) <= cp_elements(1020);
    cp_elements(1022) <= false;
    cp_elements(1023) <= cp_elements(1022);
    cp_elements(1024) <= false;
    cp_elements(1025) <= cp_elements(1024);
    cp_elements(1026) <= false;
    cp_elements(1027) <= cp_elements(1026);
    cp_elements(1028) <= OrReduce(cp_elements(754) & cp_elements(788) & cp_elements(858) & cp_elements(873) & cp_elements(906) & cp_elements(921));
    cp_elements(1029) <= cp_elements(1028);
    cp_elements(1030) <= OrReduce(cp_elements(704) & cp_elements(927) & cp_elements(933) & cp_elements(939) & cp_elements(945) & cp_elements(951));
    cp_elements(1031) <= cp_elements(1030);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal Pivot13_2199 : std_logic_vector(0 downto 0);
    signal Pivot15_2184 : std_logic_vector(0 downto 0);
    signal Pivot_2240 : std_logic_vector(0 downto 0);
    signal SwitchLeaf11_2212 : std_logic_vector(0 downto 0);
    signal SwitchLeaf7_2253 : std_logic_vector(0 downto 0);
    signal SwitchLeaf9_2225 : std_logic_vector(0 downto 0);
    signal SwitchLeaf_2266 : std_logic_vector(0 downto 0);
    signal array_obj_ref_1709_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_1709_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1709_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_1727_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_offset_scale_factor_2 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1727_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_offset_scale_factor_2 : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1736_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_1864_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_index_partial_sum_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1864_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_index_partial_sum_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_offset_scale_factor_1 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1888_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1937_constant_part_of_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1937_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1937_offset_scale_factor_0 : std_logic_vector(13 downto 0);
    signal array_obj_ref_1937_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1937_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1947_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1947_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1947_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1961_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1987_final_offset : std_logic_vector(13 downto 0);
    signal array_obj_ref_1987_resized_base_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_1987_root_address : std_logic_vector(13 downto 0);
    signal array_obj_ref_2086_constant_part_of_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_final_offset : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_index_partial_sum_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_offset_scale_factor_0 : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_offset_scale_factor_1 : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_resized_base_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_2086_root_address : std_logic_vector(4 downto 0);
    signal array_obj_ref_2105_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_2105_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_2137_root_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_constant_part_of_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_final_offset : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_index_partial_sum_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_offset_scale_factor_0 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_offset_scale_factor_1 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_offset_scale_factor_2 : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_resized_base_address : std_logic_vector(8 downto 0);
    signal array_obj_ref_2169_root_address : std_logic_vector(8 downto 0);
    signal binary_2077_wire : std_logic_vector(31 downto 0);
    signal elt1x_xi5x_xix_xi_1738 : std_logic_vector(31 downto 0);
    signal eltx_xi3x_xix_xi_1729 : std_logic_vector(31 downto 0);
    signal exitcond_1911 : std_logic_vector(0 downto 0);
    signal expr_2076_wire_constant : std_logic_vector(31 downto 0);
    signal ptr_deref_1717_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1717_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1717_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1717_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1717_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_1717_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_1741_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1741_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1741_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1741_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1741_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1745_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_1745_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1745_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_1745_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1745_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_1869_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1869_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1869_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1869_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1869_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1940_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1940_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1940_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1940_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_1940_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1940_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1954_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1954_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1954_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1954_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1954_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1954_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_1972_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_1972_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_1972_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_1972_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_1972_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_1972_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2003_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2003_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2003_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2003_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2003_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2003_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2011_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2011_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2011_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2011_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2011_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2020_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2020_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2020_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2020_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2020_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2020_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2025_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2025_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2025_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2025_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2025_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2042_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2042_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2042_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2042_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2042_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2046_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2046_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2046_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2046_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2046_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2062_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2062_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2062_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2062_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_address_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_address_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_address_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_offset_1 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_offset_2 : std_logic_vector(13 downto 0);
    signal ptr_deref_2062_word_offset_3 : std_logic_vector(13 downto 0);
    signal ptr_deref_2067_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2067_resized_base_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2067_root_address : std_logic_vector(13 downto 0);
    signal ptr_deref_2067_wire : std_logic_vector(7 downto 0);
    signal ptr_deref_2067_word_address_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2067_word_offset_0 : std_logic_vector(13 downto 0);
    signal ptr_deref_2091_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_2091_resized_base_address : std_logic_vector(4 downto 0);
    signal ptr_deref_2091_root_address : std_logic_vector(4 downto 0);
    signal ptr_deref_2091_word_address_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_2091_word_offset_0 : std_logic_vector(4 downto 0);
    signal ptr_deref_2110_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2110_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2110_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2110_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2110_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2142_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2142_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2142_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2142_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2142_word_offset_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2174_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2174_resized_base_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2174_root_address : std_logic_vector(8 downto 0);
    signal ptr_deref_2174_word_address_0 : std_logic_vector(8 downto 0);
    signal ptr_deref_2174_word_offset_0 : std_logic_vector(8 downto 0);
    signal scevgep1x_xix_xix_xix_xix_xi_1890 : std_logic_vector(31 downto 0);
    signal scevgepx_xix_xix_xix_xix_xi_1866 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1697_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1722_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1722_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1731_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1731_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_1817_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1817_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1825_data_0 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_1825_word_address_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_1861_resized : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1861_scaled : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1885_resized : std_logic_vector(13 downto 0);
    signal simple_obj_ref_1885_scaled : std_logic_vector(13 downto 0);
    signal simple_obj_ref_2083_resized : std_logic_vector(4 downto 0);
    signal simple_obj_ref_2083_scaled : std_logic_vector(4 downto 0);
    signal simple_obj_ref_2104_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_2104_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_2136_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_2136_scaled : std_logic_vector(8 downto 0);
    signal simple_obj_ref_2168_resized : std_logic_vector(8 downto 0);
    signal simple_obj_ref_2168_scaled : std_logic_vector(8 downto 0);
    signal tmp16_1703 : std_logic_vector(31 downto 0);
    signal tmp17_1710 : std_logic_vector(31 downto 0);
    signal tmp18_1714 : std_logic_vector(31 downto 0);
    signal tmp19_1718 : std_logic_vector(31 downto 0);
    signal tmp20_1751 : std_logic_vector(31 downto 0);
    signal tmp21_1756 : std_logic_vector(31 downto 0);
    signal tmp22_1762 : std_logic_vector(0 downto 0);
    signal tmp23_1775 : std_logic_vector(31 downto 0);
    signal tmp24_1778 : std_logic_vector(31 downto 0);
    signal tmp25_1793 : std_logic_vector(0 downto 0);
    signal tmp26_1808 : std_logic_vector(0 downto 0);
    signal tmp27_1818 : std_logic_vector(31 downto 0);
    signal tmp28_1824 : std_logic_vector(31 downto 0);
    signal tmp29_1835 : std_logic_vector(0 downto 0);
    signal tmp35_1845 : std_logic_vector(31 downto 0);
    signal tmp36_1852 : std_logic_vector(31 downto 0);
    signal tmp37_1870 : std_logic_vector(7 downto 0);
    signal tmp38_1876 : std_logic_vector(0 downto 0);
    signal tmp39_1893 : std_logic_vector(31 downto 0);
    signal tmp40_1905 : std_logic_vector(31 downto 0);
    signal tmp41_1924 : std_logic_vector(0 downto 0);
    signal tmp42_1938 : std_logic_vector(31 downto 0);
    signal tmp43_1948 : std_logic_vector(31 downto 0);
    signal tmp44_1952 : std_logic_vector(31 downto 0);
    signal tmp45_1962 : std_logic_vector(31 downto 0);
    signal tmp46_1966 : std_logic_vector(31 downto 0);
    signal tmp47_1970 : std_logic_vector(31 downto 0);
    signal tmp48_1979 : std_logic_vector(31 downto 0);
    signal tmp50_1988 : std_logic_vector(31 downto 0);
    signal tmp51_1994 : std_logic_vector(0 downto 0);
    signal tmp52_2012 : std_logic_vector(31 downto 0);
    signal tmp53_2018 : std_logic_vector(31 downto 0);
    signal tmp54_2026 : std_logic_vector(31 downto 0);
    signal tmp55_2032 : std_logic_vector(0 downto 0);
    signal tmp56_2043 : std_logic_vector(31 downto 0);
    signal tmp57_2047 : std_logic_vector(31 downto 0);
    signal tmp58_2052 : std_logic_vector(0 downto 0);
    signal tmp59_2063 : std_logic_vector(31 downto 0);
    signal tmp60_2088 : std_logic_vector(31 downto 0);
    signal tmp61_2092 : std_logic_vector(31 downto 0);
    signal tmp62_2098 : std_logic_vector(31 downto 0);
    signal tmp63_2107 : std_logic_vector(31 downto 0);
    signal tmp64_2111 : std_logic_vector(7 downto 0);
    signal tmp65_2117 : std_logic_vector(0 downto 0);
    signal tmp66_2139 : std_logic_vector(31 downto 0);
    signal tmp67_2143 : std_logic_vector(7 downto 0);
    signal tmp68_2149 : std_logic_vector(0 downto 0);
    signal tmp69_2171 : std_logic_vector(31 downto 0);
    signal tmp70_2175 : std_logic_vector(7 downto 0);
    signal tmp_1699 : std_logic_vector(31 downto 0);
    signal type_cast_1760_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1773_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1781_wire : std_logic_vector(31 downto 0);
    signal type_cast_1784_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1788_wire : std_logic_vector(31 downto 0);
    signal type_cast_1791_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1803_wire : std_logic_vector(31 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1822_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1830_wire : std_logic_vector(31 downto 0);
    signal type_cast_1833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1848_wire : std_logic_vector(31 downto 0);
    signal type_cast_1851_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1855_wire : std_logic_vector(31 downto 0);
    signal type_cast_1858_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1874_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1896_wire : std_logic_vector(31 downto 0);
    signal type_cast_1898_wire : std_logic_vector(31 downto 0);
    signal type_cast_1903_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1909_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1922_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1942_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_1956_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1974_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1992_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2005_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2016_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2030_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2069_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2096_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2115_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2128_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2147_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2160_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2179_wire : std_logic_vector(7 downto 0);
    signal type_cast_2182_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2194_wire : std_logic_vector(7 downto 0);
    signal type_cast_2197_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2210_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2223_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2235_wire : std_logic_vector(7 downto 0);
    signal type_cast_2238_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2251_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2264_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_2276_wire : std_logic_vector(31 downto 0);
    signal type_cast_2282_wire : std_logic_vector(31 downto 0);
    signal type_cast_2288_wire : std_logic_vector(31 downto 0);
    signal type_cast_2294_wire : std_logic_vector(31 downto 0);
    signal type_cast_2300_wire : std_logic_vector(31 downto 0);
    signal val2x_xi6x_xix_xi_1746 : std_logic_vector(31 downto 0);
    signal valx_xi4x_xix_xi_1742 : std_logic_vector(31 downto 0);
    signal xx_xsum26x_xi_2130 : std_logic_vector(31 downto 0);
    signal xx_xsum27x_xi_2162 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1709_final_offset <= "0000000000011100";
    array_obj_ref_1727_constant_part_of_offset <= "00000";
    array_obj_ref_1727_offset_scale_factor_0 <= "00101";
    array_obj_ref_1727_offset_scale_factor_1 <= "00001";
    array_obj_ref_1727_offset_scale_factor_2 <= "00001";
    array_obj_ref_1727_resized_base_address <= "00000";
    array_obj_ref_1736_constant_part_of_offset <= "00001";
    array_obj_ref_1736_offset_scale_factor_0 <= "00101";
    array_obj_ref_1736_offset_scale_factor_1 <= "00001";
    array_obj_ref_1736_offset_scale_factor_2 <= "00001";
    array_obj_ref_1736_resized_base_address <= "00000";
    array_obj_ref_1864_constant_part_of_offset <= "00000000000000";
    array_obj_ref_1864_offset_scale_factor_0 <= "00000010000000";
    array_obj_ref_1864_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1864_resized_base_address <= "00000000000000";
    array_obj_ref_1888_constant_part_of_offset <= "00000000000001";
    array_obj_ref_1888_offset_scale_factor_0 <= "00000010000000";
    array_obj_ref_1888_offset_scale_factor_1 <= "00000000000001";
    array_obj_ref_1888_resized_base_address <= "00000000000000";
    array_obj_ref_1937_constant_part_of_offset <= "11111111111111";
    array_obj_ref_1937_offset_scale_factor_0 <= "00000000000001";
    array_obj_ref_1947_final_offset <= "00000000000100";
    array_obj_ref_1961_final_offset <= "00000000001000";
    array_obj_ref_1987_final_offset <= "00000000001100";
    array_obj_ref_2086_constant_part_of_offset <= "00011";
    array_obj_ref_2086_offset_scale_factor_0 <= "00101";
    array_obj_ref_2086_offset_scale_factor_1 <= "00001";
    array_obj_ref_2086_resized_base_address <= "00000";
    array_obj_ref_2105_constant_part_of_offset <= "000000000";
    array_obj_ref_2105_offset_scale_factor_0 <= "001001000";
    array_obj_ref_2105_offset_scale_factor_1 <= "001000000";
    array_obj_ref_2105_offset_scale_factor_2 <= "000000001";
    array_obj_ref_2105_resized_base_address <= "000000000";
    array_obj_ref_2137_constant_part_of_offset <= "000000000";
    array_obj_ref_2137_offset_scale_factor_0 <= "001001000";
    array_obj_ref_2137_offset_scale_factor_1 <= "001000000";
    array_obj_ref_2137_offset_scale_factor_2 <= "000000001";
    array_obj_ref_2137_resized_base_address <= "000000000";
    array_obj_ref_2169_constant_part_of_offset <= "000000000";
    array_obj_ref_2169_offset_scale_factor_0 <= "001001000";
    array_obj_ref_2169_offset_scale_factor_1 <= "001000000";
    array_obj_ref_2169_offset_scale_factor_2 <= "000000001";
    array_obj_ref_2169_resized_base_address <= "000000000";
    expr_2076_wire_constant <= "11111111111111111111100000000000";
    ptr_deref_1717_word_offset_0 <= "0000000000000000";
    ptr_deref_1717_word_offset_1 <= "0000000000000001";
    ptr_deref_1717_word_offset_2 <= "0000000000000010";
    ptr_deref_1717_word_offset_3 <= "0000000000000011";
    ptr_deref_1741_word_offset_0 <= "00000";
    ptr_deref_1745_word_offset_0 <= "00000";
    ptr_deref_1869_word_offset_0 <= "00000000000000";
    ptr_deref_1940_word_offset_0 <= "00000000000000";
    ptr_deref_1954_word_offset_0 <= "00000000000000";
    ptr_deref_1954_word_offset_1 <= "00000000000001";
    ptr_deref_1954_word_offset_2 <= "00000000000010";
    ptr_deref_1954_word_offset_3 <= "00000000000011";
    ptr_deref_1972_word_offset_0 <= "00000000000000";
    ptr_deref_1972_word_offset_1 <= "00000000000001";
    ptr_deref_1972_word_offset_2 <= "00000000000010";
    ptr_deref_1972_word_offset_3 <= "00000000000011";
    ptr_deref_2003_word_offset_0 <= "00000000000000";
    ptr_deref_2011_word_offset_0 <= "00000000000000";
    ptr_deref_2011_word_offset_1 <= "00000000000001";
    ptr_deref_2011_word_offset_2 <= "00000000000010";
    ptr_deref_2011_word_offset_3 <= "00000000000011";
    ptr_deref_2020_word_offset_0 <= "00000000000000";
    ptr_deref_2020_word_offset_1 <= "00000000000001";
    ptr_deref_2020_word_offset_2 <= "00000000000010";
    ptr_deref_2020_word_offset_3 <= "00000000000011";
    ptr_deref_2025_word_offset_0 <= "00000000000000";
    ptr_deref_2025_word_offset_1 <= "00000000000001";
    ptr_deref_2025_word_offset_2 <= "00000000000010";
    ptr_deref_2025_word_offset_3 <= "00000000000011";
    ptr_deref_2042_word_offset_0 <= "00000000000000";
    ptr_deref_2042_word_offset_1 <= "00000000000001";
    ptr_deref_2042_word_offset_2 <= "00000000000010";
    ptr_deref_2042_word_offset_3 <= "00000000000011";
    ptr_deref_2046_word_offset_0 <= "00000000000000";
    ptr_deref_2046_word_offset_1 <= "00000000000001";
    ptr_deref_2046_word_offset_2 <= "00000000000010";
    ptr_deref_2046_word_offset_3 <= "00000000000011";
    ptr_deref_2062_word_offset_0 <= "00000000000000";
    ptr_deref_2062_word_offset_1 <= "00000000000001";
    ptr_deref_2062_word_offset_2 <= "00000000000010";
    ptr_deref_2062_word_offset_3 <= "00000000000011";
    ptr_deref_2067_word_offset_0 <= "00000000000000";
    ptr_deref_2091_word_offset_0 <= "00000";
    ptr_deref_2110_word_offset_0 <= "000000000";
    ptr_deref_2142_word_offset_0 <= "000000000";
    ptr_deref_2174_word_offset_0 <= "000000000";
    simple_obj_ref_1817_word_address_0 <= "0";
    simple_obj_ref_1825_word_address_0 <= "0";
    type_cast_1760_wire_constant <= "00000000000000000000000000000000";
    type_cast_1773_wire_constant <= "00000000000000000000000000000001";
    type_cast_1784_wire_constant <= "00000000000000000000000000000000";
    type_cast_1791_wire_constant <= "00000000000000000000000000000100";
    type_cast_1806_wire_constant <= "11111111111111111111111111111111";
    type_cast_1822_wire_constant <= "00000000000000000000000000000001";
    type_cast_1833_wire_constant <= "00000000000000000000000000000110";
    type_cast_1851_wire_constant <= "00000000000000000000000000000000";
    type_cast_1858_wire_constant <= "11111111111111111111111111111111";
    type_cast_1874_wire_constant <= "00000001";
    type_cast_1903_wire_constant <= "00000000000000000000000000000001";
    type_cast_1909_wire_constant <= "00000000000000000000000001000000";
    type_cast_1922_wire_constant <= "11111111111111111111111111111111";
    type_cast_1942_wire_constant <= "00010001";
    type_cast_1956_wire_constant <= "00000000000000000000011111110100";
    type_cast_1974_wire_constant <= "00000000000000000000000000000001";
    type_cast_1992_wire_constant <= "11111111111111111111111111111111";
    type_cast_2005_wire_constant <= "00000000";
    type_cast_2016_wire_constant <= "11111111111111111111111111111111";
    type_cast_2030_wire_constant <= "00000000000000000000000000000000";
    type_cast_2069_wire_constant <= "00000001";
    type_cast_2096_wire_constant <= "00000000000000000000000001001000";
    type_cast_2115_wire_constant <= "01110100";
    type_cast_2128_wire_constant <= "00000000000000000000000000000001";
    type_cast_2147_wire_constant <= "01101111";
    type_cast_2160_wire_constant <= "00000000000000000000000000000010";
    type_cast_2182_wire_constant <= "00110010";
    type_cast_2197_wire_constant <= "00110011";
    type_cast_2210_wire_constant <= "00110011";
    type_cast_2223_wire_constant <= "00110010";
    type_cast_2238_wire_constant <= "00110001";
    type_cast_2251_wire_constant <= "00110001";
    type_cast_2264_wire_constant <= "00110000";
    phi_stmt_1778: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1781_wire & type_cast_1784_wire_constant;
      req <= phi_stmt_1778_req_0 & phi_stmt_1778_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1778_ack_0,
          idata => idata,
          odata => tmp24_1778,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1778
    phi_stmt_1845: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1848_wire & type_cast_1851_wire_constant;
      req <= phi_stmt_1845_req_0 & phi_stmt_1845_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1845_ack_0,
          idata => idata,
          odata => tmp35_1845,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1845
    phi_stmt_1852: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1855_wire & type_cast_1858_wire_constant;
      req <= phi_stmt_1852_req_0 & phi_stmt_1852_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1852_ack_0,
          idata => idata,
          odata => tmp36_1852,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1852
    phi_stmt_1893: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1896_wire & type_cast_1898_wire;
      req <= phi_stmt_1893_req_0 & phi_stmt_1893_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1893_ack_0,
          idata => idata,
          odata => tmp39_1893,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1893
    addr_of_1728_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1727_root_address, dout => eltx_xi3x_xix_xi_1729, req => addr_of_1728_final_reg_req_0, ack => addr_of_1728_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1737_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1736_root_address, dout => elt1x_xi5x_xix_xi_1738, req => addr_of_1737_final_reg_req_0, ack => addr_of_1737_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1865_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1864_root_address, dout => scevgepx_xix_xix_xix_xix_xi_1866, req => addr_of_1865_final_reg_req_0, ack => addr_of_1865_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_1889_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1888_root_address, dout => scevgep1x_xix_xix_xix_xix_xi_1890, req => addr_of_1889_final_reg_req_0, ack => addr_of_1889_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_2087_final_reg: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2086_root_address, dout => tmp60_2088, req => addr_of_2087_final_reg_req_0, ack => addr_of_2087_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_2106_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2105_root_address, dout => tmp63_2107, req => addr_of_2106_final_reg_req_0, ack => addr_of_2106_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_2138_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2137_root_address, dout => tmp66_2139, req => addr_of_2138_final_reg_req_0, ack => addr_of_2138_final_reg_ack_0, clk => clk, reset => reset); -- 
    addr_of_2170_final_reg: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2169_root_address, dout => tmp69_2171, req => addr_of_2170_final_reg_req_0, ack => addr_of_2170_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1709_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_1703, dout => array_obj_ref_1709_resized_base_address, req => array_obj_ref_1709_base_resize_req_0, ack => array_obj_ref_1709_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1709_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1709_root_address, dout => tmp17_1710, req => array_obj_ref_1709_final_reg_req_0, ack => array_obj_ref_1709_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1727_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1778, dout => simple_obj_ref_1722_resized, req => array_obj_ref_1727_index_0_resize_req_0, ack => array_obj_ref_1727_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1727_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_1727_index_partial_sum_1, dout => array_obj_ref_1727_final_offset, req => array_obj_ref_1727_offset_inst_req_0, ack => array_obj_ref_1727_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1736_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1778, dout => simple_obj_ref_1731_resized, req => array_obj_ref_1736_index_0_resize_req_0, ack => array_obj_ref_1736_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1736_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_1736_index_partial_sum_1, dout => array_obj_ref_1736_final_offset, req => array_obj_ref_1736_offset_inst_req_0, ack => array_obj_ref_1736_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp35_1845, dout => simple_obj_ref_1861_resized, req => array_obj_ref_1864_index_0_resize_req_0, ack => array_obj_ref_1864_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1864_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1864_index_partial_sum_1, dout => array_obj_ref_1864_final_offset, req => array_obj_ref_1864_offset_inst_req_0, ack => array_obj_ref_1864_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp35_1845, dout => simple_obj_ref_1885_resized, req => array_obj_ref_1888_index_0_resize_req_0, ack => array_obj_ref_1888_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1888_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1888_index_partial_sum_1, dout => array_obj_ref_1888_final_offset, req => array_obj_ref_1888_offset_inst_req_0, ack => array_obj_ref_1888_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1937_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1893, dout => array_obj_ref_1937_resized_base_address, req => array_obj_ref_1937_base_resize_req_0, ack => array_obj_ref_1937_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1937_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1937_root_address, dout => tmp42_1938, req => array_obj_ref_1937_final_reg_req_0, ack => array_obj_ref_1937_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1937_offset_inst: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 14, flow_through => true ) 
      port map( din => array_obj_ref_1937_constant_part_of_offset, dout => array_obj_ref_1937_final_offset, req => array_obj_ref_1937_offset_inst_req_0, ack => array_obj_ref_1937_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1947_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1893, dout => array_obj_ref_1947_resized_base_address, req => array_obj_ref_1947_base_resize_req_0, ack => array_obj_ref_1947_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1947_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1947_root_address, dout => tmp43_1948, req => array_obj_ref_1947_final_reg_req_0, ack => array_obj_ref_1947_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1961_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp39_1893, dout => array_obj_ref_1961_resized_base_address, req => array_obj_ref_1961_base_resize_req_0, ack => array_obj_ref_1961_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1961_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1961_root_address, dout => tmp45_1962, req => array_obj_ref_1961_final_reg_req_0, ack => array_obj_ref_1961_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1987_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp48_1979, dout => array_obj_ref_1987_resized_base_address, req => array_obj_ref_1987_base_resize_req_0, ack => array_obj_ref_1987_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1987_final_reg: RegisterBase --
      generic map(in_data_width => 14,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_1987_root_address, dout => tmp50_1988, req => array_obj_ref_1987_final_reg_req_0, ack => array_obj_ref_1987_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2086_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp24_1778, dout => simple_obj_ref_2083_resized, req => array_obj_ref_2086_index_0_resize_req_0, ack => array_obj_ref_2086_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2086_offset_inst: RegisterBase --
      generic map(in_data_width => 5,out_data_width => 5, flow_through => true ) 
      port map( din => array_obj_ref_2086_index_partial_sum_1, dout => array_obj_ref_2086_final_offset, req => array_obj_ref_2086_offset_inst_req_0, ack => array_obj_ref_2086_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2105_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp62_2098, dout => simple_obj_ref_2104_resized, req => array_obj_ref_2105_index_2_resize_req_0, ack => array_obj_ref_2105_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2105_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_2105_index_partial_sum_1, dout => array_obj_ref_2105_final_offset, req => array_obj_ref_2105_offset_inst_req_0, ack => array_obj_ref_2105_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2137_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => xx_xsum26x_xi_2130, dout => simple_obj_ref_2136_resized, req => array_obj_ref_2137_index_2_resize_req_0, ack => array_obj_ref_2137_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2137_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_2137_index_partial_sum_1, dout => array_obj_ref_2137_final_offset, req => array_obj_ref_2137_offset_inst_req_0, ack => array_obj_ref_2137_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2169_index_2_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => xx_xsum27x_xi_2162, dout => simple_obj_ref_2168_resized, req => array_obj_ref_2169_index_2_resize_req_0, ack => array_obj_ref_2169_index_2_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2169_offset_inst: RegisterBase --
      generic map(in_data_width => 9,out_data_width => 9, flow_through => true ) 
      port map( din => array_obj_ref_2169_index_partial_sum_1, dout => array_obj_ref_2169_final_offset, req => array_obj_ref_2169_offset_inst_req_0, ack => array_obj_ref_2169_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1717_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp18_1714, dout => ptr_deref_1717_resized_base_address, req => ptr_deref_1717_base_resize_req_0, ack => ptr_deref_1717_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1741_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => eltx_xi3x_xix_xi_1729, dout => ptr_deref_1741_resized_base_address, req => ptr_deref_1741_base_resize_req_0, ack => ptr_deref_1741_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1745_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => elt1x_xi5x_xix_xi_1738, dout => ptr_deref_1745_resized_base_address, req => ptr_deref_1745_base_resize_req_0, ack => ptr_deref_1745_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1869_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => scevgepx_xix_xix_xix_xix_xi_1866, dout => ptr_deref_1869_resized_base_address, req => ptr_deref_1869_base_resize_req_0, ack => ptr_deref_1869_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1940_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp42_1938, dout => ptr_deref_1940_resized_base_address, req => ptr_deref_1940_base_resize_req_0, ack => ptr_deref_1940_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1954_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp44_1952, dout => ptr_deref_1954_resized_base_address, req => ptr_deref_1954_base_resize_req_0, ack => ptr_deref_1954_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_1972_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1970, dout => ptr_deref_1972_resized_base_address, req => ptr_deref_1972_base_resize_req_0, ack => ptr_deref_1972_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2003_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp50_1988, dout => ptr_deref_2003_resized_base_address, req => ptr_deref_2003_base_resize_req_0, ack => ptr_deref_2003_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2011_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1970, dout => ptr_deref_2011_resized_base_address, req => ptr_deref_2011_base_resize_req_0, ack => ptr_deref_2011_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2020_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1970, dout => ptr_deref_2020_resized_base_address, req => ptr_deref_2020_base_resize_req_0, ack => ptr_deref_2020_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2025_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp47_1970, dout => ptr_deref_2025_resized_base_address, req => ptr_deref_2025_base_resize_req_0, ack => ptr_deref_2025_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2042_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp44_1952, dout => ptr_deref_2042_resized_base_address, req => ptr_deref_2042_base_resize_req_0, ack => ptr_deref_2042_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2046_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp46_1966, dout => ptr_deref_2046_resized_base_address, req => ptr_deref_2046_base_resize_req_0, ack => ptr_deref_2046_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2062_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp46_1966, dout => ptr_deref_2062_resized_base_address, req => ptr_deref_2062_base_resize_req_0, ack => ptr_deref_2062_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2067_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 14, flow_through => true ) 
      port map( din => tmp42_1938, dout => ptr_deref_2067_resized_base_address, req => ptr_deref_2067_base_resize_req_0, ack => ptr_deref_2067_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2091_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 5, flow_through => true ) 
      port map( din => tmp60_2088, dout => ptr_deref_2091_resized_base_address, req => ptr_deref_2091_base_resize_req_0, ack => ptr_deref_2091_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2110_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp63_2107, dout => ptr_deref_2110_resized_base_address, req => ptr_deref_2110_base_resize_req_0, ack => ptr_deref_2110_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2142_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp66_2139, dout => ptr_deref_2142_resized_base_address, req => ptr_deref_2142_base_resize_req_0, ack => ptr_deref_2142_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2174_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 9, flow_through => true ) 
      port map( din => tmp69_2171, dout => ptr_deref_2174_resized_base_address, req => ptr_deref_2174_base_resize_req_0, ack => ptr_deref_2174_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_1698_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_1697_wire, dout => tmp_1699, req => type_cast_1698_inst_req_0, ack => type_cast_1698_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1702_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_1699, dout => tmp16_1703, req => type_cast_1702_inst_req_0, ack => type_cast_1702_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1713_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp17_1710, dout => tmp18_1714, req => type_cast_1713_inst_req_0, ack => type_cast_1713_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1781_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp23_1775, dout => type_cast_1781_wire, req => type_cast_1781_inst_req_0, ack => type_cast_1781_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1788_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp24_1778, dout => type_cast_1788_wire, req => type_cast_1788_inst_req_0, ack => type_cast_1788_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1803_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp24_1778, dout => type_cast_1803_wire, req => type_cast_1803_inst_req_0, ack => type_cast_1803_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1830_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp28_1824, dout => type_cast_1830_wire, req => type_cast_1830_inst_req_0, ack => type_cast_1830_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1848_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp40_1905, dout => type_cast_1848_wire, req => type_cast_1848_inst_req_0, ack => type_cast_1848_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1855_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp39_1893, dout => type_cast_1855_wire, req => type_cast_1855_inst_req_0, ack => type_cast_1855_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1896_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => scevgep1x_xix_xix_xix_xix_xi_1890, dout => type_cast_1896_wire, req => type_cast_1896_inst_req_0, ack => type_cast_1896_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1898_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp36_1852, dout => type_cast_1898_wire, req => type_cast_1898_inst_req_0, ack => type_cast_1898_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1951_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp43_1948, dout => tmp44_1952, req => type_cast_1951_inst_req_0, ack => type_cast_1951_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1965_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp45_1962, dout => tmp46_1966, req => type_cast_1965_inst_req_0, ack => type_cast_1965_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1969_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp39_1893, dout => tmp47_1970, req => type_cast_1969_inst_req_0, ack => type_cast_1969_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_1978_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp39_1893, dout => tmp48_1979, req => type_cast_1978_inst_req_0, ack => type_cast_1978_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2179_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_2175, dout => type_cast_2179_wire, req => type_cast_2179_inst_req_0, ack => type_cast_2179_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2194_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_2175, dout => type_cast_2194_wire, req => type_cast_2194_inst_req_0, ack => type_cast_2194_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2235_inst: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 8, flow_through => true ) 
      port map( din => tmp70_2175, dout => type_cast_2235_wire, req => type_cast_2235_inst_req_0, ack => type_cast_2235_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2276_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1699, dout => type_cast_2276_wire, req => type_cast_2276_inst_req_0, ack => type_cast_2276_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2282_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1699, dout => type_cast_2282_wire, req => type_cast_2282_inst_req_0, ack => type_cast_2282_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2288_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1699, dout => type_cast_2288_wire, req => type_cast_2288_inst_req_0, ack => type_cast_2288_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2294_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1699, dout => type_cast_2294_wire, req => type_cast_2294_inst_req_0, ack => type_cast_2294_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2300_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp_1699, dout => type_cast_2300_wire, req => type_cast_2300_inst_req_0, ack => type_cast_2300_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_1727_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_1727_root_address_inst_ack_0 <= array_obj_ref_1727_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1727_final_offset;
      array_obj_ref_1727_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_1736_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_1736_root_address_inst_ack_0 <= array_obj_ref_1736_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1736_final_offset;
      array_obj_ref_1736_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_1864_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      array_obj_ref_1864_root_address_inst_ack_0 <= array_obj_ref_1864_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1864_final_offset;
      array_obj_ref_1864_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    array_obj_ref_1888_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      array_obj_ref_1888_root_address_inst_ack_0 <= array_obj_ref_1888_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_1888_final_offset;
      array_obj_ref_1888_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    array_obj_ref_2086_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      array_obj_ref_2086_root_address_inst_ack_0 <= array_obj_ref_2086_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2086_final_offset;
      array_obj_ref_2086_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    array_obj_ref_2105_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2105_index_2_rename_ack_0 <= array_obj_ref_2105_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_2104_resized;
      simple_obj_ref_2104_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_2105_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2105_root_address_inst_ack_0 <= array_obj_ref_2105_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2105_final_offset;
      array_obj_ref_2105_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_2137_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2137_index_2_rename_ack_0 <= array_obj_ref_2137_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_2136_resized;
      simple_obj_ref_2136_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_2137_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2137_root_address_inst_ack_0 <= array_obj_ref_2137_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2137_final_offset;
      array_obj_ref_2137_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_2169_index_2_rename: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2169_index_2_rename_ack_0 <= array_obj_ref_2169_index_2_rename_req_0;
      aggregated_sig <= simple_obj_ref_2168_resized;
      simple_obj_ref_2168_scaled <= aggregated_sig(8 downto 0);
      --
    end Block;
    array_obj_ref_2169_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      array_obj_ref_2169_root_address_inst_ack_0 <= array_obj_ref_2169_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_2169_final_offset;
      array_obj_ref_2169_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_1717_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1717_gather_scatter_ack_0 <= ptr_deref_1717_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1717_data_3 & ptr_deref_1717_data_2 & ptr_deref_1717_data_1 & ptr_deref_1717_data_0;
      tmp19_1718 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1717_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_1717_root_address_inst_ack_0 <= ptr_deref_1717_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1717_resized_base_address;
      ptr_deref_1717_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_1741_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1741_addr_0_ack_0 <= ptr_deref_1741_addr_0_req_0;
      aggregated_sig <= ptr_deref_1741_root_address;
      ptr_deref_1741_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1741_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1741_gather_scatter_ack_0 <= ptr_deref_1741_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1741_data_0;
      valx_xi4x_xix_xi_1742 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1741_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1741_root_address_inst_ack_0 <= ptr_deref_1741_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1741_resized_base_address;
      ptr_deref_1741_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1745_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1745_addr_0_ack_0 <= ptr_deref_1745_addr_0_req_0;
      aggregated_sig <= ptr_deref_1745_root_address;
      ptr_deref_1745_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1745_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1745_gather_scatter_ack_0 <= ptr_deref_1745_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1745_data_0;
      val2x_xi6x_xix_xi_1746 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_1745_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_1745_root_address_inst_ack_0 <= ptr_deref_1745_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1745_resized_base_address;
      ptr_deref_1745_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_1869_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1869_addr_0_ack_0 <= ptr_deref_1869_addr_0_req_0;
      aggregated_sig <= ptr_deref_1869_root_address;
      ptr_deref_1869_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1869_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1869_gather_scatter_ack_0 <= ptr_deref_1869_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_1869_data_0;
      tmp37_1870 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1869_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1869_root_address_inst_ack_0 <= ptr_deref_1869_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1869_resized_base_address;
      ptr_deref_1869_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1940_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1940_addr_0_ack_0 <= ptr_deref_1940_addr_0_req_0;
      aggregated_sig <= ptr_deref_1940_root_address;
      ptr_deref_1940_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1940_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_1940_gather_scatter_ack_0 <= ptr_deref_1940_gather_scatter_req_0;
      aggregated_sig <= type_cast_1942_wire_constant;
      ptr_deref_1940_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1940_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1940_root_address_inst_ack_0 <= ptr_deref_1940_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1940_resized_base_address;
      ptr_deref_1940_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1954_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1954_gather_scatter_ack_0 <= ptr_deref_1954_gather_scatter_req_0;
      aggregated_sig <= type_cast_1956_wire_constant;
      ptr_deref_1954_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1954_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1954_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1954_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1954_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1954_root_address_inst_ack_0 <= ptr_deref_1954_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1954_resized_base_address;
      ptr_deref_1954_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_1972_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_1972_gather_scatter_ack_0 <= ptr_deref_1972_gather_scatter_req_0;
      aggregated_sig <= type_cast_1974_wire_constant;
      ptr_deref_1972_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_1972_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_1972_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_1972_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_1972_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_1972_root_address_inst_ack_0 <= ptr_deref_1972_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_1972_resized_base_address;
      ptr_deref_1972_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2003_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2003_addr_0_ack_0 <= ptr_deref_2003_addr_0_req_0;
      aggregated_sig <= ptr_deref_2003_root_address;
      ptr_deref_2003_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2003_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2003_gather_scatter_ack_0 <= ptr_deref_2003_gather_scatter_req_0;
      aggregated_sig <= type_cast_2005_wire_constant;
      ptr_deref_2003_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2003_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2003_root_address_inst_ack_0 <= ptr_deref_2003_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2003_resized_base_address;
      ptr_deref_2003_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2011_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2011_gather_scatter_ack_0 <= ptr_deref_2011_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2011_data_3 & ptr_deref_2011_data_2 & ptr_deref_2011_data_1 & ptr_deref_2011_data_0;
      tmp52_2012 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2011_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2011_root_address_inst_ack_0 <= ptr_deref_2011_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2011_resized_base_address;
      ptr_deref_2011_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2020_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2020_gather_scatter_ack_0 <= ptr_deref_2020_gather_scatter_req_0;
      aggregated_sig <= tmp53_2018;
      ptr_deref_2020_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2020_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2020_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2020_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2020_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2020_root_address_inst_ack_0 <= ptr_deref_2020_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2020_resized_base_address;
      ptr_deref_2020_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2025_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2025_gather_scatter_ack_0 <= ptr_deref_2025_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2025_data_3 & ptr_deref_2025_data_2 & ptr_deref_2025_data_1 & ptr_deref_2025_data_0;
      tmp54_2026 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2025_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2025_root_address_inst_ack_0 <= ptr_deref_2025_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2025_resized_base_address;
      ptr_deref_2025_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2042_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2042_gather_scatter_ack_0 <= ptr_deref_2042_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2042_data_3 & ptr_deref_2042_data_2 & ptr_deref_2042_data_1 & ptr_deref_2042_data_0;
      tmp56_2043 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2042_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2042_root_address_inst_ack_0 <= ptr_deref_2042_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2042_resized_base_address;
      ptr_deref_2042_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2046_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2046_gather_scatter_ack_0 <= ptr_deref_2046_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2046_data_3 & ptr_deref_2046_data_2 & ptr_deref_2046_data_1 & ptr_deref_2046_data_0;
      tmp57_2047 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2046_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2046_root_address_inst_ack_0 <= ptr_deref_2046_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2046_resized_base_address;
      ptr_deref_2046_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2062_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2062_gather_scatter_ack_0 <= ptr_deref_2062_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2062_data_3 & ptr_deref_2062_data_2 & ptr_deref_2062_data_1 & ptr_deref_2062_data_0;
      tmp59_2063 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2062_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2062_root_address_inst_ack_0 <= ptr_deref_2062_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2062_resized_base_address;
      ptr_deref_2062_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2067_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2067_addr_0_ack_0 <= ptr_deref_2067_addr_0_req_0;
      aggregated_sig <= ptr_deref_2067_root_address;
      ptr_deref_2067_word_address_0 <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2067_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2067_gather_scatter_ack_0 <= ptr_deref_2067_gather_scatter_req_0;
      aggregated_sig <= type_cast_2069_wire_constant;
      ptr_deref_2067_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2067_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(13 downto 0); --
    begin -- 
      ptr_deref_2067_root_address_inst_ack_0 <= ptr_deref_2067_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2067_resized_base_address;
      ptr_deref_2067_root_address <= aggregated_sig(13 downto 0);
      --
    end Block;
    ptr_deref_2091_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_2091_addr_0_ack_0 <= ptr_deref_2091_addr_0_req_0;
      aggregated_sig <= ptr_deref_2091_root_address;
      ptr_deref_2091_word_address_0 <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_2091_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2091_gather_scatter_ack_0 <= ptr_deref_2091_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2091_data_0;
      tmp61_2092 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2091_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(4 downto 0); --
    begin -- 
      ptr_deref_2091_root_address_inst_ack_0 <= ptr_deref_2091_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2091_resized_base_address;
      ptr_deref_2091_root_address <= aggregated_sig(4 downto 0);
      --
    end Block;
    ptr_deref_2110_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2110_addr_0_ack_0 <= ptr_deref_2110_addr_0_req_0;
      aggregated_sig <= ptr_deref_2110_root_address;
      ptr_deref_2110_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2110_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2110_gather_scatter_ack_0 <= ptr_deref_2110_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2110_data_0;
      tmp64_2111 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2110_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2110_root_address_inst_ack_0 <= ptr_deref_2110_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2110_resized_base_address;
      ptr_deref_2110_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2142_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2142_addr_0_ack_0 <= ptr_deref_2142_addr_0_req_0;
      aggregated_sig <= ptr_deref_2142_root_address;
      ptr_deref_2142_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2142_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2142_gather_scatter_ack_0 <= ptr_deref_2142_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2142_data_0;
      tmp67_2143 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2142_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2142_root_address_inst_ack_0 <= ptr_deref_2142_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2142_resized_base_address;
      ptr_deref_2142_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2174_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2174_addr_0_ack_0 <= ptr_deref_2174_addr_0_req_0;
      aggregated_sig <= ptr_deref_2174_root_address;
      ptr_deref_2174_word_address_0 <= aggregated_sig(8 downto 0);
      --
    end Block;
    ptr_deref_2174_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(7 downto 0); --
    begin -- 
      ptr_deref_2174_gather_scatter_ack_0 <= ptr_deref_2174_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2174_data_0;
      tmp70_2175 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2174_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(8 downto 0); --
    begin -- 
      ptr_deref_2174_root_address_inst_ack_0 <= ptr_deref_2174_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2174_resized_base_address;
      ptr_deref_2174_root_address <= aggregated_sig(8 downto 0);
      --
    end Block;
    simple_obj_ref_1817_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1817_gather_scatter_ack_0 <= simple_obj_ref_1817_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_1817_data_0;
      tmp27_1818 <= aggregated_sig(31 downto 0);
      --
    end Block;
    simple_obj_ref_1825_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      simple_obj_ref_1825_gather_scatter_ack_0 <= simple_obj_ref_1825_gather_scatter_req_0;
      aggregated_sig <= tmp28_1824;
      simple_obj_ref_1825_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    if_stmt_1763_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp22_1762;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1763_branch_req_0,
          ack0 => if_stmt_1763_branch_ack_0,
          ack1 => if_stmt_1763_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1794_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp25_1793;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1794_branch_req_0,
          ack0 => if_stmt_1794_branch_ack_0,
          ack1 => if_stmt_1794_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1809_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp26_1808;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1809_branch_req_0,
          ack0 => if_stmt_1809_branch_ack_0,
          ack1 => if_stmt_1809_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1836_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp29_1835;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1836_branch_req_0,
          ack0 => if_stmt_1836_branch_ack_0,
          ack1 => if_stmt_1836_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1877_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp38_1876;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1877_branch_req_0,
          ack0 => if_stmt_1877_branch_ack_0,
          ack1 => if_stmt_1877_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1912_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond_1911;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1912_branch_req_0,
          ack0 => if_stmt_1912_branch_ack_0,
          ack1 => if_stmt_1912_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1925_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp41_1924;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1925_branch_req_0,
          ack0 => if_stmt_1925_branch_ack_0,
          ack1 => if_stmt_1925_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1995_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp51_1994;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1995_branch_req_0,
          ack0 => if_stmt_1995_branch_ack_0,
          ack1 => if_stmt_1995_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2033_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp55_2032;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2033_branch_req_0,
          ack0 => if_stmt_2033_branch_ack_0,
          ack1 => if_stmt_2033_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2053_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp58_2052;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2053_branch_req_0,
          ack0 => if_stmt_2053_branch_ack_0,
          ack1 => if_stmt_2053_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2118_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp65_2117;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2118_branch_req_0,
          ack0 => if_stmt_2118_branch_ack_0,
          ack1 => if_stmt_2118_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2150_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= tmp68_2149;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2150_branch_req_0,
          ack0 => if_stmt_2150_branch_ack_0,
          ack1 => if_stmt_2150_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2185_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot15_2184;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2185_branch_req_0,
          ack0 => if_stmt_2185_branch_ack_0,
          ack1 => if_stmt_2185_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2200_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot13_2199;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2200_branch_req_0,
          ack0 => if_stmt_2200_branch_ack_0,
          ack1 => if_stmt_2200_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2213_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf11_2212;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2213_branch_req_0,
          ack0 => if_stmt_2213_branch_ack_0,
          ack1 => if_stmt_2213_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2226_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf9_2225;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2226_branch_req_0,
          ack0 => if_stmt_2226_branch_ack_0,
          ack1 => if_stmt_2226_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2241_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= Pivot_2240;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2241_branch_req_0,
          ack0 => if_stmt_2241_branch_ack_0,
          ack1 => if_stmt_2241_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2254_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf7_2253;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2254_branch_req_0,
          ack0 => if_stmt_2254_branch_ack_0,
          ack1 => if_stmt_2254_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_2267_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= SwitchLeaf_2266;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_2267_branch_req_0,
          ack0 => if_stmt_2267_branch_ack_0,
          ack1 => if_stmt_2267_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_1709_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1709_resized_base_address;
      array_obj_ref_1709_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000011100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1709_root_address_inst_req_0,
          ackL => array_obj_ref_1709_root_address_inst_ack_0,
          reqR => array_obj_ref_1709_root_address_inst_req_1,
          ackR => array_obj_ref_1709_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_1727_index_0_scale array_obj_ref_1736_index_0_scale array_obj_ref_2086_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(14 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1722_resized & simple_obj_ref_1731_resized & simple_obj_ref_2083_resized;
      simple_obj_ref_1722_scaled <= data_out(14 downto 10);
      simple_obj_ref_1731_scaled <= data_out(9 downto 5);
      simple_obj_ref_2083_scaled <= data_out(4 downto 0);
      reqL(2) <= array_obj_ref_1727_index_0_scale_req_0;
      reqL(1) <= array_obj_ref_1736_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_2086_index_0_scale_req_0;
      array_obj_ref_1727_index_0_scale_ack_0 <= ackL(2);
      array_obj_ref_1736_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_2086_index_0_scale_ack_0 <= ackL(0);
      reqR(2) <= array_obj_ref_1727_index_0_scale_req_1;
      reqR(1) <= array_obj_ref_1736_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_2086_index_0_scale_req_1;
      array_obj_ref_1727_index_0_scale_ack_1 <= ackR(2);
      array_obj_ref_1736_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_2086_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00101",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 3--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_1727_index_sum_1 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1722_scaled;
      array_obj_ref_1727_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00000",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1727_index_sum_1_req_0,
          ackL => array_obj_ref_1727_index_sum_1_ack_0,
          reqR => array_obj_ref_1727_index_sum_1_req_1,
          ackR => array_obj_ref_1727_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_1736_index_sum_1 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1731_scaled;
      array_obj_ref_1736_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00001",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1736_index_sum_1_req_0,
          ackL => array_obj_ref_1736_index_sum_1_ack_0,
          reqR => array_obj_ref_1736_index_sum_1_req_1,
          ackR => array_obj_ref_1736_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_1864_index_0_scale array_obj_ref_1888_index_0_scale 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(27 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1861_resized & simple_obj_ref_1885_resized;
      simple_obj_ref_1861_scaled <= data_out(27 downto 14);
      simple_obj_ref_1885_scaled <= data_out(13 downto 0);
      reqL(1) <= array_obj_ref_1864_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_1888_index_0_scale_req_0;
      array_obj_ref_1864_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_1888_index_0_scale_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_1864_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_1888_index_0_scale_req_1;
      array_obj_ref_1864_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_1888_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000010000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_1864_index_sum_1 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1861_scaled;
      array_obj_ref_1864_index_partial_sum_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1864_index_sum_1_req_0,
          ackL => array_obj_ref_1864_index_sum_1_ack_0,
          reqR => array_obj_ref_1864_index_sum_1_req_1,
          ackR => array_obj_ref_1864_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : array_obj_ref_1888_index_sum_1 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_1885_scaled;
      array_obj_ref_1888_index_partial_sum_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1888_index_sum_1_req_0,
          ackL => array_obj_ref_1888_index_sum_1_ack_0,
          reqR => array_obj_ref_1888_index_sum_1_req_1,
          ackR => array_obj_ref_1888_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : array_obj_ref_1937_root_address_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1937_final_offset & array_obj_ref_1937_resized_base_address;
      array_obj_ref_1937_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 14, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1937_root_address_inst_req_0,
          ackL => array_obj_ref_1937_root_address_inst_ack_0,
          reqR => array_obj_ref_1937_root_address_inst_req_1,
          ackR => array_obj_ref_1937_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : array_obj_ref_1947_root_address_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1947_resized_base_address;
      array_obj_ref_1947_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000100",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1947_root_address_inst_req_0,
          ackL => array_obj_ref_1947_root_address_inst_ack_0,
          reqR => array_obj_ref_1947_root_address_inst_req_1,
          ackR => array_obj_ref_1947_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : array_obj_ref_1961_root_address_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1961_resized_base_address;
      array_obj_ref_1961_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000001000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1961_root_address_inst_req_0,
          ackL => array_obj_ref_1961_root_address_inst_ack_0,
          reqR => array_obj_ref_1961_root_address_inst_req_1,
          ackR => array_obj_ref_1961_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : array_obj_ref_1987_root_address_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_1987_resized_base_address;
      array_obj_ref_1987_root_address <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000001100",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_1987_root_address_inst_req_0,
          ackL => array_obj_ref_1987_root_address_inst_ack_0,
          reqR => array_obj_ref_1987_root_address_inst_req_1,
          ackR => array_obj_ref_1987_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : array_obj_ref_2086_index_sum_1 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(4 downto 0);
      signal data_out: std_logic_vector(4 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2083_scaled;
      array_obj_ref_2086_index_partial_sum_1 <= data_out(4 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 5,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 5,
          constant_operand => "00011",
          constant_width => 5,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2086_index_sum_1_req_0,
          ackL => array_obj_ref_2086_index_sum_1_ack_0,
          reqR => array_obj_ref_2086_index_sum_1_req_1,
          ackR => array_obj_ref_2086_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : array_obj_ref_2105_index_sum_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2104_scaled;
      array_obj_ref_2105_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2105_index_sum_1_req_0,
          ackL => array_obj_ref_2105_index_sum_1_ack_0,
          reqR => array_obj_ref_2105_index_sum_1_req_1,
          ackR => array_obj_ref_2105_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : array_obj_ref_2137_index_sum_1 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2136_scaled;
      array_obj_ref_2137_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2137_index_sum_1_req_0,
          ackL => array_obj_ref_2137_index_sum_1_ack_0,
          reqR => array_obj_ref_2137_index_sum_1_req_1,
          ackR => array_obj_ref_2137_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : array_obj_ref_2169_index_sum_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(8 downto 0);
      signal data_out: std_logic_vector(8 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_2168_scaled;
      array_obj_ref_2169_index_partial_sum_1 <= data_out(8 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 9,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 9,
          constant_operand => "000000000",
          constant_width => 9,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2169_index_sum_1_req_0,
          ackL => array_obj_ref_2169_index_sum_1_ack_0,
          reqR => array_obj_ref_2169_index_sum_1_req_1,
          ackR => array_obj_ref_2169_index_sum_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_1750_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= valx_xi4x_xix_xi_1742 & tmp19_1718;
      tmp20_1751 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntXor",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1750_inst_req_0,
          ackL => binary_1750_inst_ack_0,
          reqR => binary_1750_inst_req_1,
          ackR => binary_1750_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_1755_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp20_1751 & val2x_xi6x_xix_xi_1746;
      tmp21_1756 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1755_inst_req_0,
          ackL => binary_1755_inst_ack_0,
          reqR => binary_1755_inst_req_1,
          ackR => binary_1755_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_1761_inst binary_2031_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp21_1756 & tmp54_2026;
      tmp22_1762 <= data_out(1 downto 1);
      tmp55_2032 <= data_out(0 downto 0);
      reqL(1) <= binary_1761_inst_req_0;
      reqL(0) <= binary_2031_inst_req_0;
      binary_1761_inst_ack_0 <= ackL(1);
      binary_2031_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1761_inst_req_1;
      reqR(0) <= binary_2031_inst_req_1;
      binary_1761_inst_ack_1 <= ackR(1);
      binary_2031_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_1774_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp24_1778;
      tmp23_1775 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1774_inst_req_0,
          ackL => binary_1774_inst_ack_0,
          reqR => binary_1774_inst_req_1,
          ackR => binary_1774_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_1792_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1788_wire;
      tmp25_1793 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1792_inst_req_0,
          ackL => binary_1792_inst_ack_0,
          reqR => binary_1792_inst_req_1,
          ackR => binary_1792_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_1807_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1803_wire;
      tmp26_1808 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1807_inst_req_0,
          ackL => binary_1807_inst_ack_0,
          reqR => binary_1807_inst_req_1,
          ackR => binary_1807_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_1823_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp27_1818;
      tmp28_1824 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1823_inst_req_0,
          ackL => binary_1823_inst_ack_0,
          reqR => binary_1823_inst_req_1,
          ackR => binary_1823_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_1834_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_1830_wire;
      tmp29_1835 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1834_inst_req_0,
          ackL => binary_1834_inst_ack_0,
          reqR => binary_1834_inst_req_1,
          ackR => binary_1834_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_1875_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp37_1870;
      tmp38_1876 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1875_inst_req_0,
          ackL => binary_1875_inst_ack_0,
          reqR => binary_1875_inst_req_1,
          ackR => binary_1875_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_1904_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp35_1845;
      tmp40_1905 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1904_inst_req_0,
          ackL => binary_1904_inst_ack_0,
          reqR => binary_1904_inst_req_1,
          ackR => binary_1904_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_1910_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp40_1905;
      exitcond_1911 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_1910_inst_req_0,
          ackL => binary_1910_inst_ack_0,
          reqR => binary_1910_inst_req_1,
          ackR => binary_1910_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_1923_inst binary_1993_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= tmp39_1893 & tmp50_1988;
      tmp41_1924 <= data_out(1 downto 1);
      tmp51_1994 <= data_out(0 downto 0);
      reqL(1) <= binary_1923_inst_req_0;
      reqL(0) <= binary_1993_inst_req_0;
      binary_1923_inst_ack_0 <= ackL(1);
      binary_1993_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_1923_inst_req_1;
      reqR(0) <= binary_1993_inst_req_1;
      binary_1923_inst_ack_1 <= ackR(1);
      binary_1993_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : binary_2017_inst 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp52_2012;
      tmp53_2018 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2017_inst_req_0,
          ackL => binary_2017_inst_ack_0,
          reqR => binary_2017_inst_req_1,
          ackR => binary_2017_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : binary_2051_inst 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp56_2043 & tmp57_2047;
      tmp58_2052 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2051_inst_req_0,
          ackL => binary_2051_inst_ack_0,
          reqR => binary_2051_inst_req_1,
          ackR => binary_2051_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : binary_2077_inst 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_1699;
      binary_2077_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_2077_inst_req_0,
          ackL => binary_2077_inst_ack_0,
          reqR => binary_2077_inst_req_1,
          ackR => binary_2077_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : binary_2097_inst 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp61_2092;
      tmp62_2098 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000001001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2097_inst_req_0,
          ackL => binary_2097_inst_ack_0,
          reqR => binary_2097_inst_req_1,
          ackR => binary_2097_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : binary_2116_inst 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp64_2111;
      tmp65_2117 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01110100",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2116_inst_req_0,
          ackL => binary_2116_inst_ack_0,
          reqR => binary_2116_inst_req_1,
          ackR => binary_2116_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : binary_2129_inst 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp62_2098;
      xx_xsum26x_xi_2130 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2129_inst_req_0,
          ackL => binary_2129_inst_ack_0,
          reqR => binary_2129_inst_req_1,
          ackR => binary_2129_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : binary_2148_inst 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp67_2143;
      tmp68_2149 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "01101111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2148_inst_req_0,
          ackL => binary_2148_inst_ack_0,
          reqR => binary_2148_inst_req_1,
          ackR => binary_2148_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : binary_2161_inst 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp62_2098;
      xx_xsum27x_xi_2162 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2161_inst_req_0,
          ackL => binary_2161_inst_ack_0,
          reqR => binary_2161_inst_req_1,
          ackR => binary_2161_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared split operator group (35) : binary_2183_inst 
    SplitOperatorGroup35: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2179_wire;
      Pivot15_2184 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2183_inst_req_0,
          ackL => binary_2183_inst_ack_0,
          reqR => binary_2183_inst_req_1,
          ackR => binary_2183_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 35
    -- shared split operator group (36) : binary_2198_inst 
    SplitOperatorGroup36: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2194_wire;
      Pivot13_2199 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2198_inst_req_0,
          ackL => binary_2198_inst_ack_0,
          reqR => binary_2198_inst_req_1,
          ackR => binary_2198_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 36
    -- shared split operator group (37) : binary_2211_inst 
    SplitOperatorGroup37: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_2175;
      SwitchLeaf11_2212 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110011",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2211_inst_req_0,
          ackL => binary_2211_inst_ack_0,
          reqR => binary_2211_inst_req_1,
          ackR => binary_2211_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 37
    -- shared split operator group (38) : binary_2224_inst 
    SplitOperatorGroup38: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_2175;
      SwitchLeaf9_2225 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110010",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2224_inst_req_0,
          ackL => binary_2224_inst_ack_0,
          reqR => binary_2224_inst_req_1,
          ackR => binary_2224_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 38
    -- shared split operator group (39) : binary_2239_inst 
    SplitOperatorGroup39: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2235_wire;
      Pivot_2240 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2239_inst_req_0,
          ackL => binary_2239_inst_ack_0,
          reqR => binary_2239_inst_req_1,
          ackR => binary_2239_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 39
    -- shared split operator group (40) : binary_2252_inst 
    SplitOperatorGroup40: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_2175;
      SwitchLeaf7_2253 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2252_inst_req_0,
          ackL => binary_2252_inst_ack_0,
          reqR => binary_2252_inst_req_1,
          ackR => binary_2252_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 40
    -- shared split operator group (41) : binary_2265_inst 
    SplitOperatorGroup41: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp70_2175;
      SwitchLeaf_2266 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00110000",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2265_inst_req_0,
          ackL => binary_2265_inst_ack_0,
          reqR => binary_2265_inst_req_1,
          ackR => binary_2265_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 41
    -- shared split operator group (42) : ptr_deref_1717_addr_0 
    SplitOperatorGroup42: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1717_root_address;
      ptr_deref_1717_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1717_addr_0_req_0,
          ackL => ptr_deref_1717_addr_0_ack_0,
          reqR => ptr_deref_1717_addr_0_req_1,
          ackR => ptr_deref_1717_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 42
    -- shared split operator group (43) : ptr_deref_1717_addr_1 
    SplitOperatorGroup43: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1717_root_address;
      ptr_deref_1717_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1717_addr_1_req_0,
          ackL => ptr_deref_1717_addr_1_ack_0,
          reqR => ptr_deref_1717_addr_1_req_1,
          ackR => ptr_deref_1717_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 43
    -- shared split operator group (44) : ptr_deref_1717_addr_2 
    SplitOperatorGroup44: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1717_root_address;
      ptr_deref_1717_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1717_addr_2_req_0,
          ackL => ptr_deref_1717_addr_2_ack_0,
          reqR => ptr_deref_1717_addr_2_req_1,
          ackR => ptr_deref_1717_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- shared split operator group (45) : ptr_deref_1717_addr_3 
    SplitOperatorGroup45: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1717_root_address;
      ptr_deref_1717_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1717_addr_3_req_0,
          ackL => ptr_deref_1717_addr_3_ack_0,
          reqR => ptr_deref_1717_addr_3_req_1,
          ackR => ptr_deref_1717_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 45
    -- shared split operator group (46) : ptr_deref_1954_addr_0 
    SplitOperatorGroup46: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1954_root_address;
      ptr_deref_1954_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1954_addr_0_req_0,
          ackL => ptr_deref_1954_addr_0_ack_0,
          reqR => ptr_deref_1954_addr_0_req_1,
          ackR => ptr_deref_1954_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 46
    -- shared split operator group (47) : ptr_deref_1954_addr_1 
    SplitOperatorGroup47: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1954_root_address;
      ptr_deref_1954_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1954_addr_1_req_0,
          ackL => ptr_deref_1954_addr_1_ack_0,
          reqR => ptr_deref_1954_addr_1_req_1,
          ackR => ptr_deref_1954_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 47
    -- shared split operator group (48) : ptr_deref_1954_addr_2 
    SplitOperatorGroup48: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1954_root_address;
      ptr_deref_1954_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1954_addr_2_req_0,
          ackL => ptr_deref_1954_addr_2_ack_0,
          reqR => ptr_deref_1954_addr_2_req_1,
          ackR => ptr_deref_1954_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 48
    -- shared split operator group (49) : ptr_deref_1954_addr_3 
    SplitOperatorGroup49: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1954_root_address;
      ptr_deref_1954_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1954_addr_3_req_0,
          ackL => ptr_deref_1954_addr_3_ack_0,
          reqR => ptr_deref_1954_addr_3_req_1,
          ackR => ptr_deref_1954_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 49
    -- shared split operator group (50) : ptr_deref_1972_addr_0 
    SplitOperatorGroup50: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1972_root_address;
      ptr_deref_1972_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1972_addr_0_req_0,
          ackL => ptr_deref_1972_addr_0_ack_0,
          reqR => ptr_deref_1972_addr_0_req_1,
          ackR => ptr_deref_1972_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 50
    -- shared split operator group (51) : ptr_deref_1972_addr_1 
    SplitOperatorGroup51: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1972_root_address;
      ptr_deref_1972_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1972_addr_1_req_0,
          ackL => ptr_deref_1972_addr_1_ack_0,
          reqR => ptr_deref_1972_addr_1_req_1,
          ackR => ptr_deref_1972_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 51
    -- shared split operator group (52) : ptr_deref_1972_addr_2 
    SplitOperatorGroup52: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1972_root_address;
      ptr_deref_1972_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1972_addr_2_req_0,
          ackL => ptr_deref_1972_addr_2_ack_0,
          reqR => ptr_deref_1972_addr_2_req_1,
          ackR => ptr_deref_1972_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 52
    -- shared split operator group (53) : ptr_deref_1972_addr_3 
    SplitOperatorGroup53: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_1972_root_address;
      ptr_deref_1972_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_1972_addr_3_req_0,
          ackL => ptr_deref_1972_addr_3_ack_0,
          reqR => ptr_deref_1972_addr_3_req_1,
          ackR => ptr_deref_1972_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 53
    -- shared split operator group (54) : ptr_deref_2011_addr_0 
    SplitOperatorGroup54: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2011_root_address;
      ptr_deref_2011_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2011_addr_0_req_0,
          ackL => ptr_deref_2011_addr_0_ack_0,
          reqR => ptr_deref_2011_addr_0_req_1,
          ackR => ptr_deref_2011_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 54
    -- shared split operator group (55) : ptr_deref_2011_addr_1 
    SplitOperatorGroup55: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2011_root_address;
      ptr_deref_2011_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2011_addr_1_req_0,
          ackL => ptr_deref_2011_addr_1_ack_0,
          reqR => ptr_deref_2011_addr_1_req_1,
          ackR => ptr_deref_2011_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 55
    -- shared split operator group (56) : ptr_deref_2011_addr_2 
    SplitOperatorGroup56: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2011_root_address;
      ptr_deref_2011_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2011_addr_2_req_0,
          ackL => ptr_deref_2011_addr_2_ack_0,
          reqR => ptr_deref_2011_addr_2_req_1,
          ackR => ptr_deref_2011_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 56
    -- shared split operator group (57) : ptr_deref_2011_addr_3 
    SplitOperatorGroup57: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2011_root_address;
      ptr_deref_2011_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2011_addr_3_req_0,
          ackL => ptr_deref_2011_addr_3_ack_0,
          reqR => ptr_deref_2011_addr_3_req_1,
          ackR => ptr_deref_2011_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 57
    -- shared split operator group (58) : ptr_deref_2020_addr_0 
    SplitOperatorGroup58: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2020_root_address;
      ptr_deref_2020_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2020_addr_0_req_0,
          ackL => ptr_deref_2020_addr_0_ack_0,
          reqR => ptr_deref_2020_addr_0_req_1,
          ackR => ptr_deref_2020_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 58
    -- shared split operator group (59) : ptr_deref_2020_addr_1 
    SplitOperatorGroup59: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2020_root_address;
      ptr_deref_2020_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2020_addr_1_req_0,
          ackL => ptr_deref_2020_addr_1_ack_0,
          reqR => ptr_deref_2020_addr_1_req_1,
          ackR => ptr_deref_2020_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 59
    -- shared split operator group (60) : ptr_deref_2020_addr_2 
    SplitOperatorGroup60: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2020_root_address;
      ptr_deref_2020_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2020_addr_2_req_0,
          ackL => ptr_deref_2020_addr_2_ack_0,
          reqR => ptr_deref_2020_addr_2_req_1,
          ackR => ptr_deref_2020_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 60
    -- shared split operator group (61) : ptr_deref_2020_addr_3 
    SplitOperatorGroup61: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2020_root_address;
      ptr_deref_2020_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2020_addr_3_req_0,
          ackL => ptr_deref_2020_addr_3_ack_0,
          reqR => ptr_deref_2020_addr_3_req_1,
          ackR => ptr_deref_2020_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 61
    -- shared split operator group (62) : ptr_deref_2025_addr_0 
    SplitOperatorGroup62: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2025_root_address;
      ptr_deref_2025_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2025_addr_0_req_0,
          ackL => ptr_deref_2025_addr_0_ack_0,
          reqR => ptr_deref_2025_addr_0_req_1,
          ackR => ptr_deref_2025_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 62
    -- shared split operator group (63) : ptr_deref_2025_addr_1 
    SplitOperatorGroup63: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2025_root_address;
      ptr_deref_2025_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2025_addr_1_req_0,
          ackL => ptr_deref_2025_addr_1_ack_0,
          reqR => ptr_deref_2025_addr_1_req_1,
          ackR => ptr_deref_2025_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 63
    -- shared split operator group (64) : ptr_deref_2025_addr_2 
    SplitOperatorGroup64: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2025_root_address;
      ptr_deref_2025_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2025_addr_2_req_0,
          ackL => ptr_deref_2025_addr_2_ack_0,
          reqR => ptr_deref_2025_addr_2_req_1,
          ackR => ptr_deref_2025_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 64
    -- shared split operator group (65) : ptr_deref_2025_addr_3 
    SplitOperatorGroup65: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2025_root_address;
      ptr_deref_2025_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2025_addr_3_req_0,
          ackL => ptr_deref_2025_addr_3_ack_0,
          reqR => ptr_deref_2025_addr_3_req_1,
          ackR => ptr_deref_2025_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 65
    -- shared split operator group (66) : ptr_deref_2042_addr_0 
    SplitOperatorGroup66: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2042_root_address;
      ptr_deref_2042_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2042_addr_0_req_0,
          ackL => ptr_deref_2042_addr_0_ack_0,
          reqR => ptr_deref_2042_addr_0_req_1,
          ackR => ptr_deref_2042_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 66
    -- shared split operator group (67) : ptr_deref_2042_addr_1 
    SplitOperatorGroup67: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2042_root_address;
      ptr_deref_2042_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2042_addr_1_req_0,
          ackL => ptr_deref_2042_addr_1_ack_0,
          reqR => ptr_deref_2042_addr_1_req_1,
          ackR => ptr_deref_2042_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 67
    -- shared split operator group (68) : ptr_deref_2042_addr_2 
    SplitOperatorGroup68: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2042_root_address;
      ptr_deref_2042_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2042_addr_2_req_0,
          ackL => ptr_deref_2042_addr_2_ack_0,
          reqR => ptr_deref_2042_addr_2_req_1,
          ackR => ptr_deref_2042_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 68
    -- shared split operator group (69) : ptr_deref_2042_addr_3 
    SplitOperatorGroup69: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2042_root_address;
      ptr_deref_2042_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2042_addr_3_req_0,
          ackL => ptr_deref_2042_addr_3_ack_0,
          reqR => ptr_deref_2042_addr_3_req_1,
          ackR => ptr_deref_2042_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 69
    -- shared split operator group (70) : ptr_deref_2046_addr_0 
    SplitOperatorGroup70: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2046_root_address;
      ptr_deref_2046_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2046_addr_0_req_0,
          ackL => ptr_deref_2046_addr_0_ack_0,
          reqR => ptr_deref_2046_addr_0_req_1,
          ackR => ptr_deref_2046_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 70
    -- shared split operator group (71) : ptr_deref_2046_addr_1 
    SplitOperatorGroup71: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2046_root_address;
      ptr_deref_2046_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2046_addr_1_req_0,
          ackL => ptr_deref_2046_addr_1_ack_0,
          reqR => ptr_deref_2046_addr_1_req_1,
          ackR => ptr_deref_2046_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 71
    -- shared split operator group (72) : ptr_deref_2046_addr_2 
    SplitOperatorGroup72: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2046_root_address;
      ptr_deref_2046_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2046_addr_2_req_0,
          ackL => ptr_deref_2046_addr_2_ack_0,
          reqR => ptr_deref_2046_addr_2_req_1,
          ackR => ptr_deref_2046_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 72
    -- shared split operator group (73) : ptr_deref_2046_addr_3 
    SplitOperatorGroup73: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2046_root_address;
      ptr_deref_2046_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2046_addr_3_req_0,
          ackL => ptr_deref_2046_addr_3_ack_0,
          reqR => ptr_deref_2046_addr_3_req_1,
          ackR => ptr_deref_2046_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 73
    -- shared split operator group (74) : ptr_deref_2062_addr_0 
    SplitOperatorGroup74: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2062_root_address;
      ptr_deref_2062_word_address_0 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000000",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2062_addr_0_req_0,
          ackL => ptr_deref_2062_addr_0_ack_0,
          reqR => ptr_deref_2062_addr_0_req_1,
          ackR => ptr_deref_2062_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 74
    -- shared split operator group (75) : ptr_deref_2062_addr_1 
    SplitOperatorGroup75: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2062_root_address;
      ptr_deref_2062_word_address_1 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000001",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2062_addr_1_req_0,
          ackL => ptr_deref_2062_addr_1_ack_0,
          reqR => ptr_deref_2062_addr_1_req_1,
          ackR => ptr_deref_2062_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 75
    -- shared split operator group (76) : ptr_deref_2062_addr_2 
    SplitOperatorGroup76: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2062_root_address;
      ptr_deref_2062_word_address_2 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000010",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2062_addr_2_req_0,
          ackL => ptr_deref_2062_addr_2_ack_0,
          reqR => ptr_deref_2062_addr_2_req_1,
          ackR => ptr_deref_2062_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 76
    -- shared split operator group (77) : ptr_deref_2062_addr_3 
    SplitOperatorGroup77: Block -- 
      signal data_in: std_logic_vector(13 downto 0);
      signal data_out: std_logic_vector(13 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2062_root_address;
      ptr_deref_2062_word_address_3 <= data_out(13 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 14,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 14,
          constant_operand => "00000000000011",
          constant_width => 14,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2062_addr_3_req_0,
          ackL => ptr_deref_2062_addr_3_ack_0,
          reqR => ptr_deref_2062_addr_3_req_1,
          ackR => ptr_deref_2062_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 77
    -- shared load operator group (0) : ptr_deref_1717_load_0 ptr_deref_1717_load_1 ptr_deref_1717_load_2 ptr_deref_1717_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1717_load_0_req_0,
        ptr_deref_1717_load_0_ack_0,
        ptr_deref_1717_load_0_req_1,
        ptr_deref_1717_load_0_ack_1,
        "ptr_deref_1717_load_0",
        "memory_space_5" ,
        ptr_deref_1717_data_0,
        ptr_deref_1717_word_address_0,
        "ptr_deref_1717_data_0",
        "ptr_deref_1717_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1717_load_1_req_0,
        ptr_deref_1717_load_1_ack_0,
        ptr_deref_1717_load_1_req_1,
        ptr_deref_1717_load_1_ack_1,
        "ptr_deref_1717_load_1",
        "memory_space_5" ,
        ptr_deref_1717_data_1,
        ptr_deref_1717_word_address_1,
        "ptr_deref_1717_data_1",
        "ptr_deref_1717_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1717_load_2_req_0,
        ptr_deref_1717_load_2_ack_0,
        ptr_deref_1717_load_2_req_1,
        ptr_deref_1717_load_2_ack_1,
        "ptr_deref_1717_load_2",
        "memory_space_5" ,
        ptr_deref_1717_data_2,
        ptr_deref_1717_word_address_2,
        "ptr_deref_1717_data_2",
        "ptr_deref_1717_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1717_load_3_req_0,
        ptr_deref_1717_load_3_ack_0,
        ptr_deref_1717_load_3_req_1,
        ptr_deref_1717_load_3_ack_1,
        "ptr_deref_1717_load_3",
        "memory_space_5" ,
        ptr_deref_1717_data_3,
        ptr_deref_1717_word_address_3,
        "ptr_deref_1717_data_3",
        "ptr_deref_1717_word_address_3" -- 
      );
      reqL(3) <= ptr_deref_1717_load_0_req_0;
      reqL(2) <= ptr_deref_1717_load_1_req_0;
      reqL(1) <= ptr_deref_1717_load_2_req_0;
      reqL(0) <= ptr_deref_1717_load_3_req_0;
      ptr_deref_1717_load_0_ack_0 <= ackL(3);
      ptr_deref_1717_load_1_ack_0 <= ackL(2);
      ptr_deref_1717_load_2_ack_0 <= ackL(1);
      ptr_deref_1717_load_3_ack_0 <= ackL(0);
      reqR(3) <= ptr_deref_1717_load_0_req_1;
      reqR(2) <= ptr_deref_1717_load_1_req_1;
      reqR(1) <= ptr_deref_1717_load_2_req_1;
      reqR(0) <= ptr_deref_1717_load_3_req_1;
      ptr_deref_1717_load_0_ack_1 <= ackR(3);
      ptr_deref_1717_load_1_ack_1 <= ackR(2);
      ptr_deref_1717_load_2_ack_1 <= ackR(1);
      ptr_deref_1717_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_1717_word_address_0 & ptr_deref_1717_word_address_1 & ptr_deref_1717_word_address_2 & ptr_deref_1717_word_address_3;
      ptr_deref_1717_data_0 <= data_out(31 downto 24);
      ptr_deref_1717_data_1 <= data_out(23 downto 16);
      ptr_deref_1717_data_2 <= data_out(15 downto 8);
      ptr_deref_1717_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 4,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 4,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_1741_load_0 ptr_deref_1745_load_0 ptr_deref_2091_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(14 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1741_load_0_req_0,
        ptr_deref_1741_load_0_ack_0,
        ptr_deref_1741_load_0_req_1,
        ptr_deref_1741_load_0_ack_1,
        "ptr_deref_1741_load_0",
        "memory_space_2" ,
        ptr_deref_1741_data_0,
        ptr_deref_1741_word_address_0,
        "ptr_deref_1741_data_0",
        "ptr_deref_1741_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_1745_load_0_req_0,
        ptr_deref_1745_load_0_ack_0,
        ptr_deref_1745_load_0_req_1,
        ptr_deref_1745_load_0_ack_1,
        "ptr_deref_1745_load_0",
        "memory_space_2" ,
        ptr_deref_1745_data_0,
        ptr_deref_1745_word_address_0,
        "ptr_deref_1745_data_0",
        "ptr_deref_1745_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2091_load_0_req_0,
        ptr_deref_2091_load_0_ack_0,
        ptr_deref_2091_load_0_req_1,
        ptr_deref_2091_load_0_ack_1,
        "ptr_deref_2091_load_0",
        "memory_space_2" ,
        ptr_deref_2091_data_0,
        ptr_deref_2091_word_address_0,
        "ptr_deref_2091_data_0",
        "ptr_deref_2091_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_1741_load_0_req_0;
      reqL(1) <= ptr_deref_1745_load_0_req_0;
      reqL(0) <= ptr_deref_2091_load_0_req_0;
      ptr_deref_1741_load_0_ack_0 <= ackL(2);
      ptr_deref_1745_load_0_ack_0 <= ackL(1);
      ptr_deref_2091_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_1741_load_0_req_1;
      reqR(1) <= ptr_deref_1745_load_0_req_1;
      reqR(0) <= ptr_deref_2091_load_0_req_1;
      ptr_deref_1741_load_0_ack_1 <= ackR(2);
      ptr_deref_1745_load_0_ack_1 <= ackR(1);
      ptr_deref_2091_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_1741_word_address_0 & ptr_deref_1745_word_address_0 & ptr_deref_2091_word_address_0;
      ptr_deref_1741_data_0 <= data_out(95 downto 64);
      ptr_deref_1745_data_0 <= data_out(63 downto 32);
      ptr_deref_2091_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 5,
        num_reqs => 3,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(4 downto 0),
          mtag => memory_space_2_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- shared load operator group (2) : ptr_deref_1869_load_0 ptr_deref_2011_load_0 ptr_deref_2011_load_1 ptr_deref_2011_load_2 ptr_deref_2011_load_3 ptr_deref_2025_load_0 ptr_deref_2025_load_1 ptr_deref_2025_load_2 ptr_deref_2025_load_3 ptr_deref_2042_load_0 ptr_deref_2042_load_1 ptr_deref_2042_load_2 ptr_deref_2042_load_3 ptr_deref_2046_load_0 ptr_deref_2046_load_1 ptr_deref_2046_load_2 ptr_deref_2046_load_3 ptr_deref_2062_load_0 ptr_deref_2062_load_1 ptr_deref_2062_load_2 ptr_deref_2062_load_3 
    LoadGroup2: Block -- 
      signal data_in: std_logic_vector(293 downto 0);
      signal data_out: std_logic_vector(167 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 20 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_1869_load_0_req_0,
        ptr_deref_1869_load_0_ack_0,
        ptr_deref_1869_load_0_req_1,
        ptr_deref_1869_load_0_ack_1,
        "ptr_deref_1869_load_0",
        "memory_space_3" ,
        ptr_deref_1869_data_0,
        ptr_deref_1869_word_address_0,
        "ptr_deref_1869_data_0",
        "ptr_deref_1869_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2011_load_0_req_0,
        ptr_deref_2011_load_0_ack_0,
        ptr_deref_2011_load_0_req_1,
        ptr_deref_2011_load_0_ack_1,
        "ptr_deref_2011_load_0",
        "memory_space_3" ,
        ptr_deref_2011_data_0,
        ptr_deref_2011_word_address_0,
        "ptr_deref_2011_data_0",
        "ptr_deref_2011_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2011_load_1_req_0,
        ptr_deref_2011_load_1_ack_0,
        ptr_deref_2011_load_1_req_1,
        ptr_deref_2011_load_1_ack_1,
        "ptr_deref_2011_load_1",
        "memory_space_3" ,
        ptr_deref_2011_data_1,
        ptr_deref_2011_word_address_1,
        "ptr_deref_2011_data_1",
        "ptr_deref_2011_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2011_load_2_req_0,
        ptr_deref_2011_load_2_ack_0,
        ptr_deref_2011_load_2_req_1,
        ptr_deref_2011_load_2_ack_1,
        "ptr_deref_2011_load_2",
        "memory_space_3" ,
        ptr_deref_2011_data_2,
        ptr_deref_2011_word_address_2,
        "ptr_deref_2011_data_2",
        "ptr_deref_2011_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2011_load_3_req_0,
        ptr_deref_2011_load_3_ack_0,
        ptr_deref_2011_load_3_req_1,
        ptr_deref_2011_load_3_ack_1,
        "ptr_deref_2011_load_3",
        "memory_space_3" ,
        ptr_deref_2011_data_3,
        ptr_deref_2011_word_address_3,
        "ptr_deref_2011_data_3",
        "ptr_deref_2011_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2025_load_0_req_0,
        ptr_deref_2025_load_0_ack_0,
        ptr_deref_2025_load_0_req_1,
        ptr_deref_2025_load_0_ack_1,
        "ptr_deref_2025_load_0",
        "memory_space_3" ,
        ptr_deref_2025_data_0,
        ptr_deref_2025_word_address_0,
        "ptr_deref_2025_data_0",
        "ptr_deref_2025_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2025_load_1_req_0,
        ptr_deref_2025_load_1_ack_0,
        ptr_deref_2025_load_1_req_1,
        ptr_deref_2025_load_1_ack_1,
        "ptr_deref_2025_load_1",
        "memory_space_3" ,
        ptr_deref_2025_data_1,
        ptr_deref_2025_word_address_1,
        "ptr_deref_2025_data_1",
        "ptr_deref_2025_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2025_load_2_req_0,
        ptr_deref_2025_load_2_ack_0,
        ptr_deref_2025_load_2_req_1,
        ptr_deref_2025_load_2_ack_1,
        "ptr_deref_2025_load_2",
        "memory_space_3" ,
        ptr_deref_2025_data_2,
        ptr_deref_2025_word_address_2,
        "ptr_deref_2025_data_2",
        "ptr_deref_2025_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2025_load_3_req_0,
        ptr_deref_2025_load_3_ack_0,
        ptr_deref_2025_load_3_req_1,
        ptr_deref_2025_load_3_ack_1,
        "ptr_deref_2025_load_3",
        "memory_space_3" ,
        ptr_deref_2025_data_3,
        ptr_deref_2025_word_address_3,
        "ptr_deref_2025_data_3",
        "ptr_deref_2025_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2042_load_0_req_0,
        ptr_deref_2042_load_0_ack_0,
        ptr_deref_2042_load_0_req_1,
        ptr_deref_2042_load_0_ack_1,
        "ptr_deref_2042_load_0",
        "memory_space_3" ,
        ptr_deref_2042_data_0,
        ptr_deref_2042_word_address_0,
        "ptr_deref_2042_data_0",
        "ptr_deref_2042_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2042_load_1_req_0,
        ptr_deref_2042_load_1_ack_0,
        ptr_deref_2042_load_1_req_1,
        ptr_deref_2042_load_1_ack_1,
        "ptr_deref_2042_load_1",
        "memory_space_3" ,
        ptr_deref_2042_data_1,
        ptr_deref_2042_word_address_1,
        "ptr_deref_2042_data_1",
        "ptr_deref_2042_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2042_load_2_req_0,
        ptr_deref_2042_load_2_ack_0,
        ptr_deref_2042_load_2_req_1,
        ptr_deref_2042_load_2_ack_1,
        "ptr_deref_2042_load_2",
        "memory_space_3" ,
        ptr_deref_2042_data_2,
        ptr_deref_2042_word_address_2,
        "ptr_deref_2042_data_2",
        "ptr_deref_2042_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2042_load_3_req_0,
        ptr_deref_2042_load_3_ack_0,
        ptr_deref_2042_load_3_req_1,
        ptr_deref_2042_load_3_ack_1,
        "ptr_deref_2042_load_3",
        "memory_space_3" ,
        ptr_deref_2042_data_3,
        ptr_deref_2042_word_address_3,
        "ptr_deref_2042_data_3",
        "ptr_deref_2042_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2046_load_0_req_0,
        ptr_deref_2046_load_0_ack_0,
        ptr_deref_2046_load_0_req_1,
        ptr_deref_2046_load_0_ack_1,
        "ptr_deref_2046_load_0",
        "memory_space_3" ,
        ptr_deref_2046_data_0,
        ptr_deref_2046_word_address_0,
        "ptr_deref_2046_data_0",
        "ptr_deref_2046_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2046_load_1_req_0,
        ptr_deref_2046_load_1_ack_0,
        ptr_deref_2046_load_1_req_1,
        ptr_deref_2046_load_1_ack_1,
        "ptr_deref_2046_load_1",
        "memory_space_3" ,
        ptr_deref_2046_data_1,
        ptr_deref_2046_word_address_1,
        "ptr_deref_2046_data_1",
        "ptr_deref_2046_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2046_load_2_req_0,
        ptr_deref_2046_load_2_ack_0,
        ptr_deref_2046_load_2_req_1,
        ptr_deref_2046_load_2_ack_1,
        "ptr_deref_2046_load_2",
        "memory_space_3" ,
        ptr_deref_2046_data_2,
        ptr_deref_2046_word_address_2,
        "ptr_deref_2046_data_2",
        "ptr_deref_2046_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2046_load_3_req_0,
        ptr_deref_2046_load_3_ack_0,
        ptr_deref_2046_load_3_req_1,
        ptr_deref_2046_load_3_ack_1,
        "ptr_deref_2046_load_3",
        "memory_space_3" ,
        ptr_deref_2046_data_3,
        ptr_deref_2046_word_address_3,
        "ptr_deref_2046_data_3",
        "ptr_deref_2046_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2062_load_0_req_0,
        ptr_deref_2062_load_0_ack_0,
        ptr_deref_2062_load_0_req_1,
        ptr_deref_2062_load_0_ack_1,
        "ptr_deref_2062_load_0",
        "memory_space_3" ,
        ptr_deref_2062_data_0,
        ptr_deref_2062_word_address_0,
        "ptr_deref_2062_data_0",
        "ptr_deref_2062_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2062_load_1_req_0,
        ptr_deref_2062_load_1_ack_0,
        ptr_deref_2062_load_1_req_1,
        ptr_deref_2062_load_1_ack_1,
        "ptr_deref_2062_load_1",
        "memory_space_3" ,
        ptr_deref_2062_data_1,
        ptr_deref_2062_word_address_1,
        "ptr_deref_2062_data_1",
        "ptr_deref_2062_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2062_load_2_req_0,
        ptr_deref_2062_load_2_ack_0,
        ptr_deref_2062_load_2_req_1,
        ptr_deref_2062_load_2_ack_1,
        "ptr_deref_2062_load_2",
        "memory_space_3" ,
        ptr_deref_2062_data_2,
        ptr_deref_2062_word_address_2,
        "ptr_deref_2062_data_2",
        "ptr_deref_2062_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2062_load_3_req_0,
        ptr_deref_2062_load_3_ack_0,
        ptr_deref_2062_load_3_req_1,
        ptr_deref_2062_load_3_ack_1,
        "ptr_deref_2062_load_3",
        "memory_space_3" ,
        ptr_deref_2062_data_3,
        ptr_deref_2062_word_address_3,
        "ptr_deref_2062_data_3",
        "ptr_deref_2062_word_address_3" -- 
      );
      reqL(20) <= ptr_deref_1869_load_0_req_0;
      reqL(19) <= ptr_deref_2011_load_0_req_0;
      reqL(18) <= ptr_deref_2011_load_1_req_0;
      reqL(17) <= ptr_deref_2011_load_2_req_0;
      reqL(16) <= ptr_deref_2011_load_3_req_0;
      reqL(15) <= ptr_deref_2025_load_0_req_0;
      reqL(14) <= ptr_deref_2025_load_1_req_0;
      reqL(13) <= ptr_deref_2025_load_2_req_0;
      reqL(12) <= ptr_deref_2025_load_3_req_0;
      reqL(11) <= ptr_deref_2042_load_0_req_0;
      reqL(10) <= ptr_deref_2042_load_1_req_0;
      reqL(9) <= ptr_deref_2042_load_2_req_0;
      reqL(8) <= ptr_deref_2042_load_3_req_0;
      reqL(7) <= ptr_deref_2046_load_0_req_0;
      reqL(6) <= ptr_deref_2046_load_1_req_0;
      reqL(5) <= ptr_deref_2046_load_2_req_0;
      reqL(4) <= ptr_deref_2046_load_3_req_0;
      reqL(3) <= ptr_deref_2062_load_0_req_0;
      reqL(2) <= ptr_deref_2062_load_1_req_0;
      reqL(1) <= ptr_deref_2062_load_2_req_0;
      reqL(0) <= ptr_deref_2062_load_3_req_0;
      ptr_deref_1869_load_0_ack_0 <= ackL(20);
      ptr_deref_2011_load_0_ack_0 <= ackL(19);
      ptr_deref_2011_load_1_ack_0 <= ackL(18);
      ptr_deref_2011_load_2_ack_0 <= ackL(17);
      ptr_deref_2011_load_3_ack_0 <= ackL(16);
      ptr_deref_2025_load_0_ack_0 <= ackL(15);
      ptr_deref_2025_load_1_ack_0 <= ackL(14);
      ptr_deref_2025_load_2_ack_0 <= ackL(13);
      ptr_deref_2025_load_3_ack_0 <= ackL(12);
      ptr_deref_2042_load_0_ack_0 <= ackL(11);
      ptr_deref_2042_load_1_ack_0 <= ackL(10);
      ptr_deref_2042_load_2_ack_0 <= ackL(9);
      ptr_deref_2042_load_3_ack_0 <= ackL(8);
      ptr_deref_2046_load_0_ack_0 <= ackL(7);
      ptr_deref_2046_load_1_ack_0 <= ackL(6);
      ptr_deref_2046_load_2_ack_0 <= ackL(5);
      ptr_deref_2046_load_3_ack_0 <= ackL(4);
      ptr_deref_2062_load_0_ack_0 <= ackL(3);
      ptr_deref_2062_load_1_ack_0 <= ackL(2);
      ptr_deref_2062_load_2_ack_0 <= ackL(1);
      ptr_deref_2062_load_3_ack_0 <= ackL(0);
      reqR(20) <= ptr_deref_1869_load_0_req_1;
      reqR(19) <= ptr_deref_2011_load_0_req_1;
      reqR(18) <= ptr_deref_2011_load_1_req_1;
      reqR(17) <= ptr_deref_2011_load_2_req_1;
      reqR(16) <= ptr_deref_2011_load_3_req_1;
      reqR(15) <= ptr_deref_2025_load_0_req_1;
      reqR(14) <= ptr_deref_2025_load_1_req_1;
      reqR(13) <= ptr_deref_2025_load_2_req_1;
      reqR(12) <= ptr_deref_2025_load_3_req_1;
      reqR(11) <= ptr_deref_2042_load_0_req_1;
      reqR(10) <= ptr_deref_2042_load_1_req_1;
      reqR(9) <= ptr_deref_2042_load_2_req_1;
      reqR(8) <= ptr_deref_2042_load_3_req_1;
      reqR(7) <= ptr_deref_2046_load_0_req_1;
      reqR(6) <= ptr_deref_2046_load_1_req_1;
      reqR(5) <= ptr_deref_2046_load_2_req_1;
      reqR(4) <= ptr_deref_2046_load_3_req_1;
      reqR(3) <= ptr_deref_2062_load_0_req_1;
      reqR(2) <= ptr_deref_2062_load_1_req_1;
      reqR(1) <= ptr_deref_2062_load_2_req_1;
      reqR(0) <= ptr_deref_2062_load_3_req_1;
      ptr_deref_1869_load_0_ack_1 <= ackR(20);
      ptr_deref_2011_load_0_ack_1 <= ackR(19);
      ptr_deref_2011_load_1_ack_1 <= ackR(18);
      ptr_deref_2011_load_2_ack_1 <= ackR(17);
      ptr_deref_2011_load_3_ack_1 <= ackR(16);
      ptr_deref_2025_load_0_ack_1 <= ackR(15);
      ptr_deref_2025_load_1_ack_1 <= ackR(14);
      ptr_deref_2025_load_2_ack_1 <= ackR(13);
      ptr_deref_2025_load_3_ack_1 <= ackR(12);
      ptr_deref_2042_load_0_ack_1 <= ackR(11);
      ptr_deref_2042_load_1_ack_1 <= ackR(10);
      ptr_deref_2042_load_2_ack_1 <= ackR(9);
      ptr_deref_2042_load_3_ack_1 <= ackR(8);
      ptr_deref_2046_load_0_ack_1 <= ackR(7);
      ptr_deref_2046_load_1_ack_1 <= ackR(6);
      ptr_deref_2046_load_2_ack_1 <= ackR(5);
      ptr_deref_2046_load_3_ack_1 <= ackR(4);
      ptr_deref_2062_load_0_ack_1 <= ackR(3);
      ptr_deref_2062_load_1_ack_1 <= ackR(2);
      ptr_deref_2062_load_2_ack_1 <= ackR(1);
      ptr_deref_2062_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_1869_word_address_0 & ptr_deref_2011_word_address_0 & ptr_deref_2011_word_address_1 & ptr_deref_2011_word_address_2 & ptr_deref_2011_word_address_3 & ptr_deref_2025_word_address_0 & ptr_deref_2025_word_address_1 & ptr_deref_2025_word_address_2 & ptr_deref_2025_word_address_3 & ptr_deref_2042_word_address_0 & ptr_deref_2042_word_address_1 & ptr_deref_2042_word_address_2 & ptr_deref_2042_word_address_3 & ptr_deref_2046_word_address_0 & ptr_deref_2046_word_address_1 & ptr_deref_2046_word_address_2 & ptr_deref_2046_word_address_3 & ptr_deref_2062_word_address_0 & ptr_deref_2062_word_address_1 & ptr_deref_2062_word_address_2 & ptr_deref_2062_word_address_3;
      ptr_deref_1869_data_0 <= data_out(167 downto 160);
      ptr_deref_2011_data_0 <= data_out(159 downto 152);
      ptr_deref_2011_data_1 <= data_out(151 downto 144);
      ptr_deref_2011_data_2 <= data_out(143 downto 136);
      ptr_deref_2011_data_3 <= data_out(135 downto 128);
      ptr_deref_2025_data_0 <= data_out(127 downto 120);
      ptr_deref_2025_data_1 <= data_out(119 downto 112);
      ptr_deref_2025_data_2 <= data_out(111 downto 104);
      ptr_deref_2025_data_3 <= data_out(103 downto 96);
      ptr_deref_2042_data_0 <= data_out(95 downto 88);
      ptr_deref_2042_data_1 <= data_out(87 downto 80);
      ptr_deref_2042_data_2 <= data_out(79 downto 72);
      ptr_deref_2042_data_3 <= data_out(71 downto 64);
      ptr_deref_2046_data_0 <= data_out(63 downto 56);
      ptr_deref_2046_data_1 <= data_out(55 downto 48);
      ptr_deref_2046_data_2 <= data_out(47 downto 40);
      ptr_deref_2046_data_3 <= data_out(39 downto 32);
      ptr_deref_2062_data_0 <= data_out(31 downto 24);
      ptr_deref_2062_data_1 <= data_out(23 downto 16);
      ptr_deref_2062_data_2 <= data_out(15 downto 8);
      ptr_deref_2062_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 14,
        num_reqs => 21,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_3_lr_req(0),
          mack => memory_space_3_lr_ack(0),
          maddr => memory_space_3_lr_addr(13 downto 0),
          mtag => memory_space_3_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 21,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_3_lc_req(0),
          mack => memory_space_3_lc_ack(0),
          mdata => memory_space_3_lc_data(7 downto 0),
          mtag => memory_space_3_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 2
    -- shared load operator group (3) : ptr_deref_2110_load_0 ptr_deref_2142_load_0 ptr_deref_2174_load_0 
    LoadGroup3: Block -- 
      signal data_in: std_logic_vector(26 downto 0);
      signal data_out: std_logic_vector(23 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2110_load_0_req_0,
        ptr_deref_2110_load_0_ack_0,
        ptr_deref_2110_load_0_req_1,
        ptr_deref_2110_load_0_ack_1,
        "ptr_deref_2110_load_0",
        "memory_space_1" ,
        ptr_deref_2110_data_0,
        ptr_deref_2110_word_address_0,
        "ptr_deref_2110_data_0",
        "ptr_deref_2110_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2142_load_0_req_0,
        ptr_deref_2142_load_0_ack_0,
        ptr_deref_2142_load_0_req_1,
        ptr_deref_2142_load_0_ack_1,
        "ptr_deref_2142_load_0",
        "memory_space_1" ,
        ptr_deref_2142_data_0,
        ptr_deref_2142_word_address_0,
        "ptr_deref_2142_data_0",
        "ptr_deref_2142_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2174_load_0_req_0,
        ptr_deref_2174_load_0_ack_0,
        ptr_deref_2174_load_0_req_1,
        ptr_deref_2174_load_0_ack_1,
        "ptr_deref_2174_load_0",
        "memory_space_1" ,
        ptr_deref_2174_data_0,
        ptr_deref_2174_word_address_0,
        "ptr_deref_2174_data_0",
        "ptr_deref_2174_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_2110_load_0_req_0;
      reqL(1) <= ptr_deref_2142_load_0_req_0;
      reqL(0) <= ptr_deref_2174_load_0_req_0;
      ptr_deref_2110_load_0_ack_0 <= ackL(2);
      ptr_deref_2142_load_0_ack_0 <= ackL(1);
      ptr_deref_2174_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_2110_load_0_req_1;
      reqR(1) <= ptr_deref_2142_load_0_req_1;
      reqR(0) <= ptr_deref_2174_load_0_req_1;
      ptr_deref_2110_load_0_ack_1 <= ackR(2);
      ptr_deref_2142_load_0_ack_1 <= ackR(1);
      ptr_deref_2174_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2110_word_address_0 & ptr_deref_2142_word_address_0 & ptr_deref_2174_word_address_0;
      ptr_deref_2110_data_0 <= data_out(23 downto 16);
      ptr_deref_2142_data_0 <= data_out(15 downto 8);
      ptr_deref_2174_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 9,
        num_reqs => 3,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(8 downto 0),
          mtag => memory_space_1_lr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 3,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(7 downto 0),
          mtag => memory_space_1_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 3
    -- shared load operator group (4) : simple_obj_ref_1817_load_0 
    LoadGroup4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        simple_obj_ref_1817_load_0_req_0,
        simple_obj_ref_1817_load_0_ack_0,
        simple_obj_ref_1817_load_0_req_1,
        simple_obj_ref_1817_load_0_ack_1,
        "simple_obj_ref_1817_load_0",
        "memory_space_4" ,
        simple_obj_ref_1817_data_0,
        simple_obj_ref_1817_word_address_0,
        "simple_obj_ref_1817_data_0",
        "simple_obj_ref_1817_word_address_0" -- 
      );
      reqL(0) <= simple_obj_ref_1817_load_0_req_0;
      simple_obj_ref_1817_load_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1817_load_0_req_1;
      simple_obj_ref_1817_load_0_ack_1 <= ackR(0);
      data_in <= simple_obj_ref_1817_word_address_0;
      simple_obj_ref_1817_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_4_lr_req(0),
          mack => memory_space_4_lr_ack(0),
          maddr => memory_space_4_lr_addr(0 downto 0),
          mtag => memory_space_4_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_4_lc_req(0),
          mack => memory_space_4_lc_ack(0),
          mdata => memory_space_4_lc_data(31 downto 0),
          mtag => memory_space_4_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_1940_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1940_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1940_word_address_0) &  " data ptr_deref_1940_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1940_data_0) severity note; --
        end if;
        if ptr_deref_1954_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1954_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1954_word_address_0) &  " data ptr_deref_1954_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1954_data_0) severity note; --
        end if;
        if ptr_deref_1954_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1954_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1954_word_address_1) &  " data ptr_deref_1954_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1954_data_1) severity note; --
        end if;
        if ptr_deref_1954_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1954_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1954_word_address_2) &  " data ptr_deref_1954_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1954_data_2) severity note; --
        end if;
        if ptr_deref_1954_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1954_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1954_word_address_3) &  " data ptr_deref_1954_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1954_data_3) severity note; --
        end if;
        if ptr_deref_1972_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1972_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_1972_word_address_0) &  " data ptr_deref_1972_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_1972_data_0) severity note; --
        end if;
        if ptr_deref_1972_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1972_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_1972_word_address_1) &  " data ptr_deref_1972_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_1972_data_1) severity note; --
        end if;
        if ptr_deref_1972_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1972_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_1972_word_address_2) &  " data ptr_deref_1972_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_1972_data_2) severity note; --
        end if;
        if ptr_deref_1972_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_1972_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_1972_word_address_3) &  " data ptr_deref_1972_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_1972_data_3) severity note; --
        end if;
        if ptr_deref_2003_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2003_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2003_word_address_0) &  " data ptr_deref_2003_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2003_data_0) severity note; --
        end if;
        if ptr_deref_2020_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2020_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2020_word_address_0) &  " data ptr_deref_2020_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2020_data_0) severity note; --
        end if;
        if ptr_deref_2020_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2020_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2020_word_address_1) &  " data ptr_deref_2020_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2020_data_1) severity note; --
        end if;
        if ptr_deref_2020_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2020_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2020_word_address_2) &  " data ptr_deref_2020_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2020_data_2) severity note; --
        end if;
        if ptr_deref_2020_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2020_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2020_word_address_3) &  " data ptr_deref_2020_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2020_data_3) severity note; --
        end if;
        if ptr_deref_2067_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_3 address ptr_deref_2067_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2067_word_address_0) &  " data ptr_deref_2067_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2067_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_1940_store_0 ptr_deref_1954_store_0 ptr_deref_1954_store_1 ptr_deref_1954_store_2 ptr_deref_1954_store_3 ptr_deref_1972_store_0 ptr_deref_1972_store_1 ptr_deref_1972_store_2 ptr_deref_1972_store_3 ptr_deref_2003_store_0 ptr_deref_2020_store_0 ptr_deref_2020_store_1 ptr_deref_2020_store_2 ptr_deref_2020_store_3 ptr_deref_2067_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(209 downto 0);
      signal data_in: std_logic_vector(119 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 14 downto 0);
      -- 
    begin -- 
      reqL(14) <= ptr_deref_1940_store_0_req_0;
      reqL(13) <= ptr_deref_1954_store_0_req_0;
      reqL(12) <= ptr_deref_1954_store_1_req_0;
      reqL(11) <= ptr_deref_1954_store_2_req_0;
      reqL(10) <= ptr_deref_1954_store_3_req_0;
      reqL(9) <= ptr_deref_1972_store_0_req_0;
      reqL(8) <= ptr_deref_1972_store_1_req_0;
      reqL(7) <= ptr_deref_1972_store_2_req_0;
      reqL(6) <= ptr_deref_1972_store_3_req_0;
      reqL(5) <= ptr_deref_2003_store_0_req_0;
      reqL(4) <= ptr_deref_2020_store_0_req_0;
      reqL(3) <= ptr_deref_2020_store_1_req_0;
      reqL(2) <= ptr_deref_2020_store_2_req_0;
      reqL(1) <= ptr_deref_2020_store_3_req_0;
      reqL(0) <= ptr_deref_2067_store_0_req_0;
      ptr_deref_1940_store_0_ack_0 <= ackL(14);
      ptr_deref_1954_store_0_ack_0 <= ackL(13);
      ptr_deref_1954_store_1_ack_0 <= ackL(12);
      ptr_deref_1954_store_2_ack_0 <= ackL(11);
      ptr_deref_1954_store_3_ack_0 <= ackL(10);
      ptr_deref_1972_store_0_ack_0 <= ackL(9);
      ptr_deref_1972_store_1_ack_0 <= ackL(8);
      ptr_deref_1972_store_2_ack_0 <= ackL(7);
      ptr_deref_1972_store_3_ack_0 <= ackL(6);
      ptr_deref_2003_store_0_ack_0 <= ackL(5);
      ptr_deref_2020_store_0_ack_0 <= ackL(4);
      ptr_deref_2020_store_1_ack_0 <= ackL(3);
      ptr_deref_2020_store_2_ack_0 <= ackL(2);
      ptr_deref_2020_store_3_ack_0 <= ackL(1);
      ptr_deref_2067_store_0_ack_0 <= ackL(0);
      reqR(14) <= ptr_deref_1940_store_0_req_1;
      reqR(13) <= ptr_deref_1954_store_0_req_1;
      reqR(12) <= ptr_deref_1954_store_1_req_1;
      reqR(11) <= ptr_deref_1954_store_2_req_1;
      reqR(10) <= ptr_deref_1954_store_3_req_1;
      reqR(9) <= ptr_deref_1972_store_0_req_1;
      reqR(8) <= ptr_deref_1972_store_1_req_1;
      reqR(7) <= ptr_deref_1972_store_2_req_1;
      reqR(6) <= ptr_deref_1972_store_3_req_1;
      reqR(5) <= ptr_deref_2003_store_0_req_1;
      reqR(4) <= ptr_deref_2020_store_0_req_1;
      reqR(3) <= ptr_deref_2020_store_1_req_1;
      reqR(2) <= ptr_deref_2020_store_2_req_1;
      reqR(1) <= ptr_deref_2020_store_3_req_1;
      reqR(0) <= ptr_deref_2067_store_0_req_1;
      ptr_deref_1940_store_0_ack_1 <= ackR(14);
      ptr_deref_1954_store_0_ack_1 <= ackR(13);
      ptr_deref_1954_store_1_ack_1 <= ackR(12);
      ptr_deref_1954_store_2_ack_1 <= ackR(11);
      ptr_deref_1954_store_3_ack_1 <= ackR(10);
      ptr_deref_1972_store_0_ack_1 <= ackR(9);
      ptr_deref_1972_store_1_ack_1 <= ackR(8);
      ptr_deref_1972_store_2_ack_1 <= ackR(7);
      ptr_deref_1972_store_3_ack_1 <= ackR(6);
      ptr_deref_2003_store_0_ack_1 <= ackR(5);
      ptr_deref_2020_store_0_ack_1 <= ackR(4);
      ptr_deref_2020_store_1_ack_1 <= ackR(3);
      ptr_deref_2020_store_2_ack_1 <= ackR(2);
      ptr_deref_2020_store_3_ack_1 <= ackR(1);
      ptr_deref_2067_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_1940_word_address_0 & ptr_deref_1954_word_address_0 & ptr_deref_1954_word_address_1 & ptr_deref_1954_word_address_2 & ptr_deref_1954_word_address_3 & ptr_deref_1972_word_address_0 & ptr_deref_1972_word_address_1 & ptr_deref_1972_word_address_2 & ptr_deref_1972_word_address_3 & ptr_deref_2003_word_address_0 & ptr_deref_2020_word_address_0 & ptr_deref_2020_word_address_1 & ptr_deref_2020_word_address_2 & ptr_deref_2020_word_address_3 & ptr_deref_2067_word_address_0;
      data_in <= ptr_deref_1940_data_0 & ptr_deref_1954_data_0 & ptr_deref_1954_data_1 & ptr_deref_1954_data_2 & ptr_deref_1954_data_3 & ptr_deref_1972_data_0 & ptr_deref_1972_data_1 & ptr_deref_1972_data_2 & ptr_deref_1972_data_3 & ptr_deref_2003_data_0 & ptr_deref_2020_data_0 & ptr_deref_2020_data_1 & ptr_deref_2020_data_2 & ptr_deref_2020_data_3 & ptr_deref_2067_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 14,
        data_width => 8,
        num_reqs => 15,
        tag_length => 5,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_3_sr_req(0),
          mack => memory_space_3_sr_ack(0),
          maddr => memory_space_3_sr_addr(13 downto 0),
          mdata => memory_space_3_sr_data(7 downto 0),
          mtag => memory_space_3_sr_tag(7 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 15,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_3_sc_req(0),
          mack => memory_space_3_sc_ack(0),
          mtag => memory_space_3_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_1825_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_4 address simple_obj_ref_1825_word_address_0 ="  &  convert_slv_to_hex_string(simple_obj_ref_1825_word_address_0) &  " data simple_obj_ref_1825_data_0 ="  &  convert_slv_to_hex_string(simple_obj_ref_1825_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (1) : simple_obj_ref_1825_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= simple_obj_ref_1825_store_0_req_0;
      simple_obj_ref_1825_store_0_ack_0 <= ackL(0);
      reqR(0) <= simple_obj_ref_1825_store_0_req_1;
      simple_obj_ref_1825_store_0_ack_1 <= ackR(0);
      addr_in <= simple_obj_ref_1825_word_address_0;
      data_in <= simple_obj_ref_1825_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_4_sr_req(0),
          mack => memory_space_4_sr_ack(0),
          maddr => memory_space_4_sr_addr(0 downto 0),
          mdata => memory_space_4_sr_data(31 downto 0),
          mtag => memory_space_4_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_4_sc_req(0),
          mack => memory_space_4_sc_ack(0),
          mtag => memory_space_4_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_1697_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_1697_inst_ack_0 then -- 
            assert false report " ReadPipe rtt_in0 to wire simple_obj_ref_1697_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_1697_inst_req_0;
      simple_obj_ref_1697_inst_ack_0 <= ack(0);
      simple_obj_ref_1697_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => rtt_in0_pipe_read_req(0),
          oack => rtt_in0_pipe_read_ack(0),
          odata => rtt_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2074_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_2077_wire value="  &  convert_slv_to_hex_string(binary_2077_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2074_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2074_inst_req_0;
      simple_obj_ref_2074_inst_ack_0 <= ack(0);
      data_in <= binary_2077_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2274_inst_ack_0 then -- 
          assert false report " WritePipe to0_in0 from wire type_cast_2276_wire value="  &  convert_slv_to_hex_string(type_cast_2276_wire) severity note; --
        end if;
        if simple_obj_ref_2298_inst_ack_0 then -- 
          assert false report " WritePipe to0_in0 from wire type_cast_2300_wire value="  &  convert_slv_to_hex_string(type_cast_2300_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2274_inst simple_obj_ref_2298_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_2274_inst_req_0;
      req(0) <= simple_obj_ref_2298_inst_req_0;
      simple_obj_ref_2274_inst_ack_0 <= ack(1);
      simple_obj_ref_2298_inst_ack_0 <= ack(0);
      data_in <= type_cast_2276_wire & type_cast_2300_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to0_in0_pipe_write_req(0),
          oack => to0_in0_pipe_write_ack(0),
          odata => to0_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2280_inst_ack_0 then -- 
          assert false report " WritePipe to1_in0 from wire type_cast_2282_wire value="  &  convert_slv_to_hex_string(type_cast_2282_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_2280_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2280_inst_req_0;
      simple_obj_ref_2280_inst_ack_0 <= ack(0);
      data_in <= type_cast_2282_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to1_in0_pipe_write_req(0),
          oack => to1_in0_pipe_write_ack(0),
          odata => to1_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2286_inst_ack_0 then -- 
          assert false report " WritePipe to2_in0 from wire type_cast_2288_wire value="  &  convert_slv_to_hex_string(type_cast_2288_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_2286_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2286_inst_req_0;
      simple_obj_ref_2286_inst_ack_0 <= ack(0);
      data_in <= type_cast_2288_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to2_in0_pipe_write_req(0),
          oack => to2_in0_pipe_write_ack(0),
          odata => to2_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2292_inst_ack_0 then -- 
          assert false report " WritePipe to3_in0 from wire type_cast_2294_wire value="  &  convert_slv_to_hex_string(type_cast_2294_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (4) : simple_obj_ref_2292_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2292_inst_req_0;
      simple_obj_ref_2292_inst_ack_0 <= ack(0);
      data_in <= type_cast_2294_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => to3_in0_pipe_write_req(0),
          oack => to3_in0_pipe_write_ack(0),
          odata => to3_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_src is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    src_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    src_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    src_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    chk_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    chk_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    chk_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_src;
architecture Default of ahir_glue_src is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_src_CP_10923_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_2365_base_resize_req_0 : boolean;
  signal array_obj_ref_2365_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2365_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2365_root_address_inst_req_0 : boolean;
  signal binary_2354_inst_ack_1 : boolean;
  signal type_cast_2358_inst_req_0 : boolean;
  signal binary_2354_inst_req_1 : boolean;
  signal binary_2354_inst_ack_0 : boolean;
  signal type_cast_2358_inst_ack_0 : boolean;
  signal binary_2354_inst_req_0 : boolean;
  signal ptr_deref_2368_addr_0_ack_1 : boolean;
  signal ptr_deref_2368_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2368_root_address_inst_req_0 : boolean;
  signal ptr_deref_2368_base_resize_ack_0 : boolean;
  signal ptr_deref_2368_base_resize_req_0 : boolean;
  signal array_obj_ref_2365_base_resize_ack_0 : boolean;
  signal ptr_deref_2383_addr_0_ack_0 : boolean;
  signal ptr_deref_2383_addr_0_req_1 : boolean;
  signal ptr_deref_2383_addr_0_ack_1 : boolean;
  signal array_obj_ref_2394_index_0_resize_req_0 : boolean;
  signal array_obj_ref_2365_root_address_inst_ack_1 : boolean;
  signal call_stmt_2387_call_req_0 : boolean;
  signal call_stmt_2387_call_ack_0 : boolean;
  signal call_stmt_2387_call_req_1 : boolean;
  signal call_stmt_2387_call_ack_1 : boolean;
  signal binary_2375_inst_req_1 : boolean;
  signal binary_2375_inst_ack_1 : boolean;
  signal array_obj_ref_2394_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_2394_index_0_rename_req_0 : boolean;
  signal array_obj_ref_2394_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_2394_offset_inst_req_0 : boolean;
  signal array_obj_ref_2394_offset_inst_ack_0 : boolean;
  signal binary_2375_inst_req_0 : boolean;
  signal binary_2375_inst_ack_0 : boolean;
  signal type_cast_2390_inst_req_0 : boolean;
  signal type_cast_2390_inst_ack_0 : boolean;
  signal array_obj_ref_2365_final_reg_req_0 : boolean;
  signal ptr_deref_2368_addr_0_ack_0 : boolean;
  signal ptr_deref_2368_store_0_req_0 : boolean;
  signal ptr_deref_2368_store_0_ack_0 : boolean;
  signal type_cast_2379_inst_req_0 : boolean;
  signal type_cast_2379_inst_ack_0 : boolean;
  signal ptr_deref_2368_addr_3_req_0 : boolean;
  signal ptr_deref_2368_store_1_req_0 : boolean;
  signal ptr_deref_2368_store_1_ack_0 : boolean;
  signal ptr_deref_2383_base_resize_req_0 : boolean;
  signal ptr_deref_2368_store_0_req_1 : boolean;
  signal ptr_deref_2368_store_0_ack_1 : boolean;
  signal ptr_deref_2368_addr_2_req_0 : boolean;
  signal ptr_deref_2368_addr_2_ack_0 : boolean;
  signal ptr_deref_2368_addr_1_req_1 : boolean;
  signal ptr_deref_2368_addr_1_ack_1 : boolean;
  signal ptr_deref_2368_store_2_req_1 : boolean;
  signal ptr_deref_2368_store_1_req_1 : boolean;
  signal ptr_deref_2383_load_0_req_0 : boolean;
  signal ptr_deref_2368_store_2_req_0 : boolean;
  signal ptr_deref_2368_store_2_ack_0 : boolean;
  signal ptr_deref_2368_addr_3_ack_0 : boolean;
  signal ptr_deref_2368_addr_3_req_1 : boolean;
  signal ptr_deref_2368_addr_1_req_0 : boolean;
  signal ptr_deref_2368_addr_1_ack_0 : boolean;
  signal ptr_deref_2368_store_2_ack_1 : boolean;
  signal ptr_deref_2383_load_0_req_1 : boolean;
  signal ptr_deref_2383_load_0_ack_1 : boolean;
  signal ptr_deref_2383_load_1_req_1 : boolean;
  signal ptr_deref_2368_store_1_ack_1 : boolean;
  signal ptr_deref_2368_addr_3_ack_1 : boolean;
  signal ptr_deref_2368_store_3_req_0 : boolean;
  signal ptr_deref_2368_store_3_ack_0 : boolean;
  signal ptr_deref_2383_root_address_inst_req_0 : boolean;
  signal ptr_deref_2383_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2383_addr_1_ack_1 : boolean;
  signal ptr_deref_2368_store_3_req_1 : boolean;
  signal ptr_deref_2368_store_3_ack_1 : boolean;
  signal ptr_deref_2368_addr_2_req_1 : boolean;
  signal ptr_deref_2368_addr_2_ack_1 : boolean;
  signal ptr_deref_2383_addr_0_req_0 : boolean;
  signal ptr_deref_2383_load_1_ack_1 : boolean;
  signal ptr_deref_2383_gather_scatter_req_0 : boolean;
  signal ptr_deref_2383_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2368_addr_0_req_1 : boolean;
  signal ptr_deref_2383_base_resize_ack_0 : boolean;
  signal array_obj_ref_2365_final_reg_ack_0 : boolean;
  signal ptr_deref_2383_load_0_ack_0 : boolean;
  signal ptr_deref_2383_load_1_req_0 : boolean;
  signal ptr_deref_2383_load_1_ack_0 : boolean;
  signal ptr_deref_2368_addr_0_req_0 : boolean;
  signal ptr_deref_2383_addr_1_req_0 : boolean;
  signal ptr_deref_2383_addr_1_ack_0 : boolean;
  signal ptr_deref_2383_addr_1_req_1 : boolean;
  signal simple_obj_ref_2311_inst_req_0 : boolean;
  signal simple_obj_ref_2311_inst_ack_0 : boolean;
  signal type_cast_2312_inst_req_0 : boolean;
  signal type_cast_2312_inst_ack_0 : boolean;
  signal binary_2318_inst_req_0 : boolean;
  signal binary_2318_inst_ack_0 : boolean;
  signal binary_2318_inst_req_1 : boolean;
  signal binary_2318_inst_ack_1 : boolean;
  signal binary_2324_inst_req_0 : boolean;
  signal binary_2324_inst_ack_0 : boolean;
  signal binary_2324_inst_req_1 : boolean;
  signal binary_2324_inst_ack_1 : boolean;
  signal type_cast_2328_inst_req_0 : boolean;
  signal type_cast_2328_inst_ack_0 : boolean;
  signal type_cast_2332_inst_req_0 : boolean;
  signal type_cast_2332_inst_ack_0 : boolean;
  signal array_obj_ref_2337_base_resize_req_0 : boolean;
  signal array_obj_ref_2337_base_resize_ack_0 : boolean;
  signal ptr_deref_2368_gather_scatter_req_0 : boolean;
  signal ptr_deref_2368_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2337_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2337_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2337_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2337_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2337_final_reg_req_0 : boolean;
  signal array_obj_ref_2337_final_reg_ack_0 : boolean;
  signal array_obj_ref_2344_base_resize_req_0 : boolean;
  signal array_obj_ref_2344_base_resize_ack_0 : boolean;
  signal array_obj_ref_2344_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2344_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2344_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2344_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2344_final_reg_req_0 : boolean;
  signal array_obj_ref_2344_final_reg_ack_0 : boolean;
  signal ptr_deref_2347_base_resize_req_0 : boolean;
  signal ptr_deref_2347_base_resize_ack_0 : boolean;
  signal ptr_deref_2347_root_address_inst_req_0 : boolean;
  signal ptr_deref_2347_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2347_addr_0_req_0 : boolean;
  signal ptr_deref_2347_addr_0_ack_0 : boolean;
  signal ptr_deref_2347_addr_0_req_1 : boolean;
  signal ptr_deref_2347_addr_0_ack_1 : boolean;
  signal ptr_deref_2347_addr_1_req_0 : boolean;
  signal ptr_deref_2347_addr_1_ack_0 : boolean;
  signal ptr_deref_2347_addr_1_req_1 : boolean;
  signal ptr_deref_2347_addr_1_ack_1 : boolean;
  signal ptr_deref_2347_addr_2_req_0 : boolean;
  signal ptr_deref_2347_addr_2_ack_0 : boolean;
  signal ptr_deref_2347_addr_2_req_1 : boolean;
  signal ptr_deref_2347_addr_2_ack_1 : boolean;
  signal ptr_deref_2347_addr_3_req_0 : boolean;
  signal ptr_deref_2347_addr_3_ack_0 : boolean;
  signal ptr_deref_2347_addr_3_req_1 : boolean;
  signal ptr_deref_2347_addr_3_ack_1 : boolean;
  signal ptr_deref_2347_gather_scatter_req_0 : boolean;
  signal ptr_deref_2347_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2347_store_0_req_0 : boolean;
  signal ptr_deref_2347_store_0_ack_0 : boolean;
  signal ptr_deref_2347_store_1_req_0 : boolean;
  signal ptr_deref_2347_store_1_ack_0 : boolean;
  signal ptr_deref_2347_store_2_req_0 : boolean;
  signal ptr_deref_2347_store_2_ack_0 : boolean;
  signal ptr_deref_2347_store_3_req_0 : boolean;
  signal ptr_deref_2347_store_3_ack_0 : boolean;
  signal ptr_deref_2347_store_0_req_1 : boolean;
  signal ptr_deref_2347_store_0_ack_1 : boolean;
  signal ptr_deref_2347_store_1_req_1 : boolean;
  signal ptr_deref_2347_store_1_ack_1 : boolean;
  signal ptr_deref_2347_store_2_req_1 : boolean;
  signal ptr_deref_2347_store_2_ack_1 : boolean;
  signal ptr_deref_2347_store_3_req_1 : boolean;
  signal ptr_deref_2347_store_3_ack_1 : boolean;
  signal array_obj_ref_2394_base_resize_req_0 : boolean;
  signal array_obj_ref_2394_base_resize_ack_0 : boolean;
  signal array_obj_ref_2394_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2394_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2394_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2394_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2394_final_reg_req_0 : boolean;
  signal array_obj_ref_2394_final_reg_ack_0 : boolean;
  signal array_obj_ref_2401_base_resize_req_0 : boolean;
  signal array_obj_ref_2401_base_resize_ack_0 : boolean;
  signal array_obj_ref_2401_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2401_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2401_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2401_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2401_final_reg_req_0 : boolean;
  signal array_obj_ref_2401_final_reg_ack_0 : boolean;
  signal ptr_deref_2404_base_resize_req_0 : boolean;
  signal ptr_deref_2404_base_resize_ack_0 : boolean;
  signal ptr_deref_2404_root_address_inst_req_0 : boolean;
  signal ptr_deref_2404_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2404_addr_0_req_0 : boolean;
  signal ptr_deref_2404_addr_0_ack_0 : boolean;
  signal ptr_deref_2404_addr_0_req_1 : boolean;
  signal ptr_deref_2404_addr_0_ack_1 : boolean;
  signal ptr_deref_2404_addr_1_req_0 : boolean;
  signal ptr_deref_2404_addr_1_ack_0 : boolean;
  signal ptr_deref_2404_addr_1_req_1 : boolean;
  signal ptr_deref_2404_addr_1_ack_1 : boolean;
  signal ptr_deref_2404_addr_2_req_0 : boolean;
  signal ptr_deref_2404_addr_2_ack_0 : boolean;
  signal ptr_deref_2404_addr_2_req_1 : boolean;
  signal ptr_deref_2404_addr_2_ack_1 : boolean;
  signal ptr_deref_2404_addr_3_req_0 : boolean;
  signal ptr_deref_2404_addr_3_ack_0 : boolean;
  signal ptr_deref_2404_addr_3_req_1 : boolean;
  signal ptr_deref_2404_addr_3_ack_1 : boolean;
  signal ptr_deref_2404_gather_scatter_req_0 : boolean;
  signal ptr_deref_2404_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2404_store_0_req_0 : boolean;
  signal ptr_deref_2404_store_0_ack_0 : boolean;
  signal ptr_deref_2404_store_1_req_0 : boolean;
  signal ptr_deref_2404_store_1_ack_0 : boolean;
  signal ptr_deref_2404_store_2_req_0 : boolean;
  signal ptr_deref_2404_store_2_ack_0 : boolean;
  signal ptr_deref_2404_store_3_req_0 : boolean;
  signal ptr_deref_2404_store_3_ack_0 : boolean;
  signal ptr_deref_2404_store_0_req_1 : boolean;
  signal ptr_deref_2404_store_0_ack_1 : boolean;
  signal ptr_deref_2404_store_1_req_1 : boolean;
  signal ptr_deref_2404_store_1_ack_1 : boolean;
  signal ptr_deref_2404_store_2_req_1 : boolean;
  signal ptr_deref_2404_store_2_ack_1 : boolean;
  signal ptr_deref_2404_store_3_req_1 : boolean;
  signal ptr_deref_2404_store_3_ack_1 : boolean;
  signal binary_2411_inst_req_0 : boolean;
  signal binary_2411_inst_ack_0 : boolean;
  signal binary_2411_inst_req_1 : boolean;
  signal binary_2411_inst_ack_1 : boolean;
  signal binary_2417_inst_req_0 : boolean;
  signal binary_2417_inst_ack_0 : boolean;
  signal binary_2417_inst_req_1 : boolean;
  signal binary_2417_inst_ack_1 : boolean;
  signal type_cast_2421_inst_req_0 : boolean;
  signal type_cast_2421_inst_ack_0 : boolean;
  signal array_obj_ref_2428_base_resize_req_0 : boolean;
  signal array_obj_ref_2428_base_resize_ack_0 : boolean;
  signal array_obj_ref_2428_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2428_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2428_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2428_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2428_final_reg_req_0 : boolean;
  signal array_obj_ref_2428_final_reg_ack_0 : boolean;
  signal ptr_deref_2431_base_resize_req_0 : boolean;
  signal ptr_deref_2431_base_resize_ack_0 : boolean;
  signal ptr_deref_2431_root_address_inst_req_0 : boolean;
  signal ptr_deref_2431_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2431_addr_0_req_0 : boolean;
  signal ptr_deref_2431_addr_0_ack_0 : boolean;
  signal ptr_deref_2431_addr_0_req_1 : boolean;
  signal ptr_deref_2431_addr_0_ack_1 : boolean;
  signal ptr_deref_2431_addr_1_req_0 : boolean;
  signal ptr_deref_2431_addr_1_ack_0 : boolean;
  signal ptr_deref_2431_addr_1_req_1 : boolean;
  signal ptr_deref_2431_addr_1_ack_1 : boolean;
  signal ptr_deref_2431_addr_2_req_0 : boolean;
  signal ptr_deref_2431_addr_2_ack_0 : boolean;
  signal ptr_deref_2431_addr_2_req_1 : boolean;
  signal ptr_deref_2431_addr_2_ack_1 : boolean;
  signal ptr_deref_2431_addr_3_req_0 : boolean;
  signal ptr_deref_2431_addr_3_ack_0 : boolean;
  signal ptr_deref_2431_addr_3_req_1 : boolean;
  signal ptr_deref_2431_addr_3_ack_1 : boolean;
  signal ptr_deref_2431_gather_scatter_req_0 : boolean;
  signal ptr_deref_2431_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2431_store_0_req_0 : boolean;
  signal ptr_deref_2431_store_0_ack_0 : boolean;
  signal ptr_deref_2431_store_1_req_0 : boolean;
  signal ptr_deref_2431_store_1_ack_0 : boolean;
  signal ptr_deref_2431_store_2_req_0 : boolean;
  signal ptr_deref_2431_store_2_ack_0 : boolean;
  signal ptr_deref_2431_store_3_req_0 : boolean;
  signal ptr_deref_2431_store_3_ack_0 : boolean;
  signal ptr_deref_2431_store_0_req_1 : boolean;
  signal ptr_deref_2431_store_0_ack_1 : boolean;
  signal ptr_deref_2431_store_1_req_1 : boolean;
  signal ptr_deref_2431_store_1_ack_1 : boolean;
  signal ptr_deref_2431_store_2_req_1 : boolean;
  signal ptr_deref_2431_store_2_ack_1 : boolean;
  signal ptr_deref_2431_store_3_req_1 : boolean;
  signal ptr_deref_2431_store_3_ack_1 : boolean;
  signal type_cast_2436_inst_req_0 : boolean;
  signal type_cast_2436_inst_ack_0 : boolean;
  signal simple_obj_ref_2434_inst_req_0 : boolean;
  signal simple_obj_ref_2434_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_src_CP_10923: Block -- control-path 
    signal cp_elements: BooleanArray(283 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(283);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(283), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(159);
    crr_11416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2387_call_req_0); -- 
    cp_elements(2) <= cp_elements(277);
    cp_elements(3) <= cp_elements(0);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(5) & cp_elements(7));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10959_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => type_cast_2312_inst_req_0); -- 
    cp_elements(5) <= cp_elements(3);
    cp_elements(6) <= cp_elements(3);
    req_10954_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => simple_obj_ref_2311_inst_req_0); -- 
    ack_10955_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2311_inst_ack_0, ack => cp_elements(7)); -- 
    ack_10960_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2312_inst_ack_0, ack => cp_elements(8)); -- 
    cp_elements(9) <= cp_elements(8);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(12));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_2318_inst_req_0); -- 
    cp_elements(11) <= cp_elements(9);
    cp_elements(12) <= cp_elements(9);
    ra_10973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2318_inst_ack_0, ack => cp_elements(13)); -- 
    cr_10974_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => binary_2318_inst_req_1); -- 
    cp_elements(14) <= binary_2318_inst_ack_1;
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_10984_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2324_inst_req_0); -- 
    cp_elements(16) <= cp_elements(9);
    cp_elements(17) <= cp_elements(14);
    ra_10985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2324_inst_ack_0, ack => cp_elements(18)); -- 
    cr_10986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2324_inst_req_1); -- 
    cp_elements(19) <= binary_2324_inst_ack_1;
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(21) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_10996_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2328_inst_req_0); -- 
    cp_elements(21) <= cp_elements(9);
    cp_elements(22) <= cp_elements(19);
    cp_elements(23) <= type_cast_2328_inst_ack_0;
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(25) & cp_elements(26));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => type_cast_2332_inst_req_0); -- 
    cp_elements(25) <= cp_elements(9);
    cp_elements(26) <= cp_elements(19);
    ack_11007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2332_inst_ack_0, ack => cp_elements(27)); -- 
    base_resize_req_11018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => array_obj_ref_2337_base_resize_req_0); -- 
    cp_elements(28) <= cp_elements(9);
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(28) & cp_elements(32));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => array_obj_ref_2337_final_reg_req_0); -- 
    base_resize_ack_11019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2337_base_resize_ack_0, ack => cp_elements(30)); -- 
    plus_base_rr_11024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => array_obj_ref_2337_root_address_inst_req_0); -- 
    plus_base_ra_11025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2337_root_address_inst_ack_0, ack => cp_elements(31)); -- 
    plus_base_cr_11026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => array_obj_ref_2337_root_address_inst_req_1); -- 
    plus_base_ca_11027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2337_root_address_inst_ack_1, ack => cp_elements(32)); -- 
    final_reg_ack_11032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2337_final_reg_ack_0, ack => cp_elements(33)); -- 
    cp_elements(34) <= cp_elements(9);
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => array_obj_ref_2344_final_reg_req_0); -- 
    cp_elements(36) <= cp_elements(23);
    base_resize_req_11043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => array_obj_ref_2344_base_resize_req_0); -- 
    base_resize_ack_11044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2344_base_resize_ack_0, ack => cp_elements(37)); -- 
    plus_base_rr_11049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => array_obj_ref_2344_root_address_inst_req_0); -- 
    plus_base_ra_11050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2344_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    plus_base_cr_11051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => array_obj_ref_2344_root_address_inst_req_1); -- 
    plus_base_ca_11052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2344_root_address_inst_ack_1, ack => cp_elements(39)); -- 
    final_reg_ack_11057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2344_final_reg_ack_0, ack => cp_elements(40)); -- 
    base_resize_req_11071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_2347_base_resize_req_0); -- 
    cpelement_group_41 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(33) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(41),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11112_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2347_gather_scatter_req_0); -- 
    base_resize_ack_11072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_base_resize_ack_0, ack => cp_elements(42)); -- 
    sum_rename_req_11076_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_2347_root_address_inst_req_0); -- 
    cp_elements(43) <= ptr_deref_2347_root_address_inst_ack_0;
    cp_elements(44) <= cp_elements(43);
    rr_11084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_2347_addr_0_req_0); -- 
    ra_11085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_0_ack_0, ack => cp_elements(45)); -- 
    cr_11086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => ptr_deref_2347_addr_0_req_1); -- 
    ca_11087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_0_ack_1, ack => cp_elements(46)); -- 
    cp_elements(47) <= cp_elements(43);
    rr_11091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2347_addr_1_req_0); -- 
    ra_11092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_1_ack_0, ack => cp_elements(48)); -- 
    cr_11093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => ptr_deref_2347_addr_1_req_1); -- 
    ca_11094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_1_ack_1, ack => cp_elements(49)); -- 
    cp_elements(50) <= cp_elements(43);
    rr_11098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => ptr_deref_2347_addr_2_req_0); -- 
    ra_11099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_2_ack_0, ack => cp_elements(51)); -- 
    cr_11100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => ptr_deref_2347_addr_2_req_1); -- 
    ca_11101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_2_ack_1, ack => cp_elements(52)); -- 
    cp_elements(53) <= cp_elements(43);
    rr_11105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => ptr_deref_2347_addr_3_req_0); -- 
    ra_11106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_3_ack_0, ack => cp_elements(54)); -- 
    cr_11107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => ptr_deref_2347_addr_3_req_1); -- 
    ca_11108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_addr_3_ack_1, ack => cp_elements(55)); -- 
    cpelement_group_56 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(46) & cp_elements(49) & cp_elements(52) & cp_elements(55));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(56),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(57) <= ptr_deref_2347_gather_scatter_ack_0;
    cp_elements(58) <= cp_elements(57);
    rr_11120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_2347_store_0_req_0); -- 
    ra_11121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_0_ack_0, ack => cp_elements(59)); -- 
    cp_elements(60) <= cp_elements(57);
    rr_11125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => ptr_deref_2347_store_1_req_0); -- 
    ra_11126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_1_ack_0, ack => cp_elements(61)); -- 
    cp_elements(62) <= cp_elements(57);
    rr_11130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_2347_store_2_req_0); -- 
    ra_11131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_2_ack_0, ack => cp_elements(63)); -- 
    cp_elements(64) <= cp_elements(57);
    rr_11135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_2347_store_3_req_0); -- 
    ra_11136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_3_ack_0, ack => cp_elements(65)); -- 
    cpelement_group_66 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(59) & cp_elements(61) & cp_elements(63) & cp_elements(65));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(66),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(67) <= cp_elements(66);
    cp_elements(68) <= cp_elements(67);
    cr_11146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_2347_store_0_req_1); -- 
    ca_11147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_0_ack_1, ack => cp_elements(69)); -- 
    cp_elements(70) <= cp_elements(67);
    cr_11151_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_2347_store_1_req_1); -- 
    ca_11152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_1_ack_1, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(67);
    cr_11156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_2347_store_2_req_1); -- 
    ca_11157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_2_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= cp_elements(67);
    cr_11161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_2347_store_3_req_1); -- 
    ca_11162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2347_store_3_ack_1, ack => cp_elements(75)); -- 
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(69) & cp_elements(71) & cp_elements(73) & cp_elements(75));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(79));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => binary_2354_inst_req_0); -- 
    cp_elements(78) <= cp_elements(9);
    cp_elements(79) <= cp_elements(14);
    ra_11172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2354_inst_ack_0, ack => cp_elements(80)); -- 
    cr_11173_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => binary_2354_inst_req_1); -- 
    ca_11174_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2354_inst_ack_1, ack => cp_elements(81)); -- 
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(83));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11183_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => type_cast_2358_inst_req_0); -- 
    cp_elements(83) <= cp_elements(9);
    ack_11184_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2358_inst_ack_0, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(9);
    cpelement_group_86 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(85) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(86),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => array_obj_ref_2365_final_reg_req_0); -- 
    cp_elements(87) <= cp_elements(23);
    base_resize_req_11195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => array_obj_ref_2365_base_resize_req_0); -- 
    base_resize_ack_11196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2365_base_resize_ack_0, ack => cp_elements(88)); -- 
    plus_base_rr_11201_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => array_obj_ref_2365_root_address_inst_req_0); -- 
    plus_base_ra_11202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2365_root_address_inst_ack_0, ack => cp_elements(89)); -- 
    plus_base_cr_11203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => array_obj_ref_2365_root_address_inst_req_1); -- 
    plus_base_ca_11204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2365_root_address_inst_ack_1, ack => cp_elements(90)); -- 
    cp_elements(91) <= array_obj_ref_2365_final_reg_ack_0;
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(84) & cp_elements(91) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2368_gather_scatter_req_0); -- 
    cp_elements(93) <= cp_elements(91);
    base_resize_req_11223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => ptr_deref_2368_base_resize_req_0); -- 
    base_resize_ack_11224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_base_resize_ack_0, ack => cp_elements(94)); -- 
    sum_rename_req_11228_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2368_root_address_inst_req_0); -- 
    cp_elements(95) <= ptr_deref_2368_root_address_inst_ack_0;
    cp_elements(96) <= cp_elements(95);
    rr_11236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2368_addr_0_req_0); -- 
    ra_11237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_0_ack_0, ack => cp_elements(97)); -- 
    cr_11238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => ptr_deref_2368_addr_0_req_1); -- 
    ca_11239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_0_ack_1, ack => cp_elements(98)); -- 
    cp_elements(99) <= cp_elements(95);
    rr_11243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => ptr_deref_2368_addr_1_req_0); -- 
    ra_11244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_1_ack_0, ack => cp_elements(100)); -- 
    cr_11245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => ptr_deref_2368_addr_1_req_1); -- 
    ca_11246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_1_ack_1, ack => cp_elements(101)); -- 
    cp_elements(102) <= cp_elements(95);
    rr_11250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => ptr_deref_2368_addr_2_req_0); -- 
    ra_11251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_2_ack_0, ack => cp_elements(103)); -- 
    cr_11252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2368_addr_2_req_1); -- 
    ca_11253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_2_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(95);
    rr_11257_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2368_addr_3_req_0); -- 
    ra_11258_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_3_ack_0, ack => cp_elements(106)); -- 
    cr_11259_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => ptr_deref_2368_addr_3_req_1); -- 
    ca_11260_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_addr_3_ack_1, ack => cp_elements(107)); -- 
    cpelement_group_108 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(98) & cp_elements(101) & cp_elements(104) & cp_elements(107));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(108),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(109) <= ptr_deref_2368_gather_scatter_ack_0;
    cp_elements(110) <= cp_elements(109);
    rr_11272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_2368_store_0_req_0); -- 
    ra_11273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_0_ack_0, ack => cp_elements(111)); -- 
    cp_elements(112) <= cp_elements(109);
    rr_11277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => ptr_deref_2368_store_1_req_0); -- 
    ra_11278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_1_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(109);
    rr_11282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_2368_store_2_req_0); -- 
    ra_11283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_2_ack_0, ack => cp_elements(115)); -- 
    cp_elements(116) <= cp_elements(109);
    rr_11287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => ptr_deref_2368_store_3_req_0); -- 
    ra_11288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_3_ack_0, ack => cp_elements(117)); -- 
    cpelement_group_118 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(111) & cp_elements(113) & cp_elements(115) & cp_elements(117));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(118),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(119) <= cp_elements(118);
    cp_elements(120) <= cp_elements(119);
    cr_11298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => ptr_deref_2368_store_0_req_1); -- 
    ca_11299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_0_ack_1, ack => cp_elements(121)); -- 
    cp_elements(122) <= cp_elements(119);
    cr_11303_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2368_store_1_req_1); -- 
    ca_11304_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_1_ack_1, ack => cp_elements(123)); -- 
    cp_elements(124) <= cp_elements(119);
    cr_11308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => ptr_deref_2368_store_2_req_1); -- 
    ca_11309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_2_ack_1, ack => cp_elements(125)); -- 
    cp_elements(126) <= cp_elements(119);
    cr_11313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2368_store_3_req_1); -- 
    ca_11314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2368_store_3_ack_1, ack => cp_elements(127)); -- 
    cpelement_group_128 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(121) & cp_elements(123) & cp_elements(125) & cp_elements(127));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(128),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(130) & cp_elements(131));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => binary_2375_inst_req_0); -- 
    cp_elements(130) <= cp_elements(9);
    cp_elements(131) <= cp_elements(14);
    ra_11324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2375_inst_ack_0, ack => cp_elements(132)); -- 
    cr_11325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => binary_2375_inst_req_1); -- 
    ca_11326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2375_inst_ack_1, ack => cp_elements(133)); -- 
    cpelement_group_134 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(133) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(134),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => type_cast_2379_inst_req_0); -- 
    cp_elements(135) <= cp_elements(9);
    cp_elements(136) <= type_cast_2379_inst_ack_0;
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(118) & cp_elements(136) & cp_elements(147));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(136);
    base_resize_req_11349_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2383_base_resize_req_0); -- 
    base_resize_ack_11350_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_base_resize_ack_0, ack => cp_elements(139)); -- 
    sum_rename_req_11354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => ptr_deref_2383_root_address_inst_req_0); -- 
    cp_elements(140) <= ptr_deref_2383_root_address_inst_ack_0;
    cp_elements(141) <= cp_elements(140);
    rr_11362_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(141), ack => ptr_deref_2383_addr_0_req_0); -- 
    ra_11363_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_addr_0_ack_0, ack => cp_elements(142)); -- 
    cr_11364_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2383_addr_0_req_1); -- 
    ca_11365_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_addr_0_ack_1, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(140);
    rr_11369_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2383_addr_1_req_0); -- 
    ra_11370_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_addr_1_ack_0, ack => cp_elements(145)); -- 
    cr_11371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => ptr_deref_2383_addr_1_req_1); -- 
    ca_11372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_addr_1_ack_1, ack => cp_elements(146)); -- 
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(146));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(148) <= cp_elements(137);
    rr_11382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => ptr_deref_2383_load_0_req_0); -- 
    ra_11383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_load_0_ack_0, ack => cp_elements(149)); -- 
    cp_elements(150) <= cp_elements(137);
    rr_11387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => ptr_deref_2383_load_1_req_0); -- 
    ra_11388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_load_1_ack_0, ack => cp_elements(151)); -- 
    cpelement_group_152 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(151));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(152),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(153) <= cp_elements(152);
    cr_11398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2383_load_0_req_1); -- 
    ca_11399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_load_0_ack_1, ack => cp_elements(154)); -- 
    cp_elements(155) <= cp_elements(152);
    cr_11403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2383_load_1_req_1); -- 
    ca_11404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_load_1_ack_1, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(154) & cp_elements(156));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_11405_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => ptr_deref_2383_gather_scatter_req_0); -- 
    merge_ack_11406_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2383_gather_scatter_ack_0, ack => cp_elements(158)); -- 
    cpelement_group_159 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(128) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(159),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_11417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2387_call_ack_0, ack => cp_elements(160)); -- 
    ccr_11421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => call_stmt_2387_call_req_1); -- 
    cca_11422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2387_call_ack_1, ack => cp_elements(161)); -- 
    cp_elements(162) <= cp_elements(161);
    cpelement_group_163 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(164) & cp_elements(165));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(163),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => type_cast_2390_inst_req_0); -- 
    cp_elements(164) <= cp_elements(162);
    cp_elements(165) <= cp_elements(162);
    ack_11437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2390_inst_ack_0, ack => cp_elements(166)); -- 
    index_resize_req_11452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => array_obj_ref_2394_index_0_resize_req_0); -- 
    cp_elements(167) <= cp_elements(162);
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(167) & cp_elements(176));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => array_obj_ref_2394_final_reg_req_0); -- 
    cp_elements(169) <= cp_elements(162);
    base_resize_req_11468_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => array_obj_ref_2394_base_resize_req_0); -- 
    index_resize_ack_11453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_index_0_resize_ack_0, ack => cp_elements(170)); -- 
    scale_rename_req_11457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => array_obj_ref_2394_index_0_rename_req_0); -- 
    scale_rename_ack_11458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_index_0_rename_ack_0, ack => cp_elements(171)); -- 
    final_index_req_11462_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => array_obj_ref_2394_offset_inst_req_0); -- 
    final_index_ack_11463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_offset_inst_ack_0, ack => cp_elements(172)); -- 
    base_resize_ack_11469_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_base_resize_ack_0, ack => cp_elements(173)); -- 
    cpelement_group_174 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(173));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(174),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_11474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(174), ack => array_obj_ref_2394_root_address_inst_req_0); -- 
    plus_base_ra_11475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_root_address_inst_ack_0, ack => cp_elements(175)); -- 
    plus_base_cr_11476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => array_obj_ref_2394_root_address_inst_req_1); -- 
    plus_base_ca_11477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_root_address_inst_ack_1, ack => cp_elements(176)); -- 
    final_reg_ack_11482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2394_final_reg_ack_0, ack => cp_elements(177)); -- 
    cp_elements(178) <= cp_elements(162);
    cpelement_group_179 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(178) & cp_elements(183));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(179),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => array_obj_ref_2401_final_reg_req_0); -- 
    cp_elements(180) <= cp_elements(162);
    base_resize_req_11493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => array_obj_ref_2401_base_resize_req_0); -- 
    base_resize_ack_11494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2401_base_resize_ack_0, ack => cp_elements(181)); -- 
    plus_base_rr_11499_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => array_obj_ref_2401_root_address_inst_req_0); -- 
    plus_base_ra_11500_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2401_root_address_inst_ack_0, ack => cp_elements(182)); -- 
    plus_base_cr_11501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(182), ack => array_obj_ref_2401_root_address_inst_req_1); -- 
    plus_base_ca_11502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2401_root_address_inst_ack_1, ack => cp_elements(183)); -- 
    cp_elements(184) <= array_obj_ref_2401_final_reg_ack_0;
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(177) & cp_elements(184) & cp_elements(201));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => ptr_deref_2404_gather_scatter_req_0); -- 
    cp_elements(186) <= cp_elements(184);
    base_resize_req_11521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => ptr_deref_2404_base_resize_req_0); -- 
    base_resize_ack_11522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_base_resize_ack_0, ack => cp_elements(187)); -- 
    sum_rename_req_11526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => ptr_deref_2404_root_address_inst_req_0); -- 
    cp_elements(188) <= ptr_deref_2404_root_address_inst_ack_0;
    cp_elements(189) <= cp_elements(188);
    rr_11534_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => ptr_deref_2404_addr_0_req_0); -- 
    ra_11535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_0_ack_0, ack => cp_elements(190)); -- 
    cr_11536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_2404_addr_0_req_1); -- 
    ca_11537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_0_ack_1, ack => cp_elements(191)); -- 
    cp_elements(192) <= cp_elements(188);
    rr_11541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => ptr_deref_2404_addr_1_req_0); -- 
    ra_11542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_1_ack_0, ack => cp_elements(193)); -- 
    cr_11543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => ptr_deref_2404_addr_1_req_1); -- 
    ca_11544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_1_ack_1, ack => cp_elements(194)); -- 
    cp_elements(195) <= cp_elements(188);
    rr_11548_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => ptr_deref_2404_addr_2_req_0); -- 
    ra_11549_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_2_ack_0, ack => cp_elements(196)); -- 
    cr_11550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ptr_deref_2404_addr_2_req_1); -- 
    ca_11551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_2_ack_1, ack => cp_elements(197)); -- 
    cp_elements(198) <= cp_elements(188);
    rr_11555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => ptr_deref_2404_addr_3_req_0); -- 
    ra_11556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_3_ack_0, ack => cp_elements(199)); -- 
    cr_11557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => ptr_deref_2404_addr_3_req_1); -- 
    ca_11558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_addr_3_ack_1, ack => cp_elements(200)); -- 
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(194) & cp_elements(197) & cp_elements(200));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(202) <= ptr_deref_2404_gather_scatter_ack_0;
    cp_elements(203) <= cp_elements(202);
    rr_11570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => ptr_deref_2404_store_0_req_0); -- 
    ra_11571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_0_ack_0, ack => cp_elements(204)); -- 
    cp_elements(205) <= cp_elements(202);
    rr_11575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => ptr_deref_2404_store_1_req_0); -- 
    ra_11576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_1_ack_0, ack => cp_elements(206)); -- 
    cp_elements(207) <= cp_elements(202);
    rr_11580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2404_store_2_req_0); -- 
    ra_11581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_2_ack_0, ack => cp_elements(208)); -- 
    cp_elements(209) <= cp_elements(202);
    rr_11585_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2404_store_3_req_0); -- 
    ra_11586_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_3_ack_0, ack => cp_elements(210)); -- 
    cpelement_group_211 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(204) & cp_elements(206) & cp_elements(208) & cp_elements(210));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(211),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(212) <= cp_elements(211);
    cp_elements(213) <= cp_elements(212);
    cr_11596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2404_store_0_req_1); -- 
    ca_11597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_0_ack_1, ack => cp_elements(214)); -- 
    cp_elements(215) <= cp_elements(212);
    cr_11601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => ptr_deref_2404_store_1_req_1); -- 
    ca_11602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_1_ack_1, ack => cp_elements(216)); -- 
    cp_elements(217) <= cp_elements(212);
    cr_11606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2404_store_2_req_1); -- 
    ca_11607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_2_ack_1, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(212);
    cr_11611_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2404_store_3_req_1); -- 
    ca_11612_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2404_store_3_ack_1, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(214) & cp_elements(216) & cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_222 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(224));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(222),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => binary_2411_inst_req_0); -- 
    cp_elements(223) <= cp_elements(162);
    cp_elements(224) <= cp_elements(162);
    ra_11622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2411_inst_ack_0, ack => cp_elements(225)); -- 
    cr_11623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => binary_2411_inst_req_1); -- 
    ca_11624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2411_inst_ack_1, ack => cp_elements(226)); -- 
    cpelement_group_227 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(226) & cp_elements(228));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(227),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => binary_2417_inst_req_0); -- 
    cp_elements(228) <= cp_elements(162);
    ra_11634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2417_inst_ack_0, ack => cp_elements(229)); -- 
    cr_11635_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => binary_2417_inst_req_1); -- 
    ca_11636_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2417_inst_ack_1, ack => cp_elements(230)); -- 
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11645_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => type_cast_2421_inst_req_0); -- 
    cp_elements(232) <= cp_elements(162);
    ack_11646_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2421_inst_ack_0, ack => cp_elements(233)); -- 
    cp_elements(234) <= cp_elements(162);
    cpelement_group_235 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(234) & cp_elements(239));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(235),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_11670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(235), ack => array_obj_ref_2428_final_reg_req_0); -- 
    cp_elements(236) <= cp_elements(162);
    base_resize_req_11657_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => array_obj_ref_2428_base_resize_req_0); -- 
    base_resize_ack_11658_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2428_base_resize_ack_0, ack => cp_elements(237)); -- 
    plus_base_rr_11663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => array_obj_ref_2428_root_address_inst_req_0); -- 
    plus_base_ra_11664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2428_root_address_inst_ack_0, ack => cp_elements(238)); -- 
    plus_base_cr_11665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => array_obj_ref_2428_root_address_inst_req_1); -- 
    plus_base_ca_11666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2428_root_address_inst_ack_1, ack => cp_elements(239)); -- 
    cp_elements(240) <= array_obj_ref_2428_final_reg_ack_0;
    cpelement_group_241 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(233) & cp_elements(240) & cp_elements(257));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(241),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11726_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(241), ack => ptr_deref_2431_gather_scatter_req_0); -- 
    cp_elements(242) <= cp_elements(240);
    base_resize_req_11685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => ptr_deref_2431_base_resize_req_0); -- 
    base_resize_ack_11686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_base_resize_ack_0, ack => cp_elements(243)); -- 
    sum_rename_req_11690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(243), ack => ptr_deref_2431_root_address_inst_req_0); -- 
    cp_elements(244) <= ptr_deref_2431_root_address_inst_ack_0;
    cp_elements(245) <= cp_elements(244);
    rr_11698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(245), ack => ptr_deref_2431_addr_0_req_0); -- 
    ra_11699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_0_ack_0, ack => cp_elements(246)); -- 
    cr_11700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2431_addr_0_req_1); -- 
    ca_11701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_0_ack_1, ack => cp_elements(247)); -- 
    cp_elements(248) <= cp_elements(244);
    rr_11705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => ptr_deref_2431_addr_1_req_0); -- 
    ra_11706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_1_ack_0, ack => cp_elements(249)); -- 
    cr_11707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => ptr_deref_2431_addr_1_req_1); -- 
    ca_11708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_1_ack_1, ack => cp_elements(250)); -- 
    cp_elements(251) <= cp_elements(244);
    rr_11712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => ptr_deref_2431_addr_2_req_0); -- 
    ra_11713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_2_ack_0, ack => cp_elements(252)); -- 
    cr_11714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2431_addr_2_req_1); -- 
    ca_11715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_2_ack_1, ack => cp_elements(253)); -- 
    cp_elements(254) <= cp_elements(244);
    rr_11719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => ptr_deref_2431_addr_3_req_0); -- 
    ra_11720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_3_ack_0, ack => cp_elements(255)); -- 
    cr_11721_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => ptr_deref_2431_addr_3_req_1); -- 
    ca_11722_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_addr_3_ack_1, ack => cp_elements(256)); -- 
    cpelement_group_257 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(247) & cp_elements(250) & cp_elements(253) & cp_elements(256));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(257),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(258) <= ptr_deref_2431_gather_scatter_ack_0;
    cp_elements(259) <= cp_elements(258);
    rr_11734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(259), ack => ptr_deref_2431_store_0_req_0); -- 
    ra_11735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_0_ack_0, ack => cp_elements(260)); -- 
    cp_elements(261) <= cp_elements(258);
    rr_11739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2431_store_1_req_0); -- 
    ra_11740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_1_ack_0, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(258);
    rr_11744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2431_store_2_req_0); -- 
    ra_11745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_2_ack_0, ack => cp_elements(264)); -- 
    cp_elements(265) <= cp_elements(258);
    rr_11749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => ptr_deref_2431_store_3_req_0); -- 
    ra_11750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_3_ack_0, ack => cp_elements(266)); -- 
    cpelement_group_267 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(260) & cp_elements(262) & cp_elements(264) & cp_elements(266));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(267),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(268) <= cp_elements(267);
    cr_11760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => ptr_deref_2431_store_0_req_1); -- 
    ca_11761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_0_ack_1, ack => cp_elements(269)); -- 
    cp_elements(270) <= cp_elements(267);
    cr_11765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2431_store_1_req_1); -- 
    ca_11766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_1_ack_1, ack => cp_elements(271)); -- 
    cp_elements(272) <= cp_elements(267);
    cr_11770_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(272), ack => ptr_deref_2431_store_2_req_1); -- 
    ca_11771_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_2_ack_1, ack => cp_elements(273)); -- 
    cp_elements(274) <= cp_elements(267);
    cr_11775_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => ptr_deref_2431_store_3_req_1); -- 
    ca_11776_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2431_store_3_ack_1, ack => cp_elements(275)); -- 
    cpelement_group_276 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(269) & cp_elements(271) & cp_elements(273) & cp_elements(275));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(276),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(221) & cp_elements(276));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(278) <= cp_elements(2);
    cpelement_group_279 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(280) & cp_elements(281));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(279),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => type_cast_2436_inst_req_0); -- 
    cp_elements(280) <= cp_elements(278);
    cp_elements(281) <= cp_elements(278);
    ack_11789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2436_inst_ack_0, ack => cp_elements(282)); -- 
    pipe_wreq_11794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => simple_obj_ref_2434_inst_req_0); -- 
    pipe_wack_11795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2434_inst_ack_0, ack => cp_elements(283)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2337_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2337_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2337_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2344_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2344_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2344_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2365_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2365_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2365_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2394_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2394_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_2394_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2394_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2401_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2401_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2401_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2428_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2428_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2428_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2347_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2347_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2347_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2347_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2347_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2347_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2368_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2368_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2368_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2368_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2368_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2368_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2383_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2383_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2383_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2404_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2404_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2404_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2404_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2404_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2404_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2431_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2431_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2431_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2431_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_2431_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2431_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2311_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_2393_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2393_scaled : std_logic_vector(15 downto 0);
    signal tmp10_2376 : std_logic_vector(31 downto 0);
    signal tmp11_2380 : std_logic_vector(31 downto 0);
    signal tmp12_2384 : std_logic_vector(15 downto 0);
    signal tmp13_2387 : std_logic_vector(15 downto 0);
    signal tmp14_2391 : std_logic_vector(31 downto 0);
    signal tmp15_2395 : std_logic_vector(31 downto 0);
    signal tmp16_2402 : std_logic_vector(31 downto 0);
    signal tmp17_2412 : std_logic_vector(31 downto 0);
    signal tmp18_2418 : std_logic_vector(31 downto 0);
    signal tmp19_2422 : std_logic_vector(31 downto 0);
    signal tmp1_2319 : std_logic_vector(31 downto 0);
    signal tmp20_2429 : std_logic_vector(31 downto 0);
    signal tmp2_2325 : std_logic_vector(31 downto 0);
    signal tmp3_2329 : std_logic_vector(31 downto 0);
    signal tmp4_2333 : std_logic_vector(31 downto 0);
    signal tmp5_2338 : std_logic_vector(31 downto 0);
    signal tmp6_2345 : std_logic_vector(31 downto 0);
    signal tmp7_2355 : std_logic_vector(31 downto 0);
    signal tmp8_2359 : std_logic_vector(31 downto 0);
    signal tmp9_2366 : std_logic_vector(31 downto 0);
    signal tmp_2313 : std_logic_vector(31 downto 0);
    signal type_cast_2317_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2323_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2353_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2374_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2410_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2416_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2436_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_2337_final_offset <= "0000000001101100";
    array_obj_ref_2344_final_offset <= "0000000000001000";
    array_obj_ref_2365_final_offset <= "0000000000001100";
    array_obj_ref_2394_offset_scale_factor_0 <= "0000000000000001";
    array_obj_ref_2401_final_offset <= "0000000000010000";
    array_obj_ref_2428_final_offset <= "0000000000010100";
    ptr_deref_2347_word_offset_0 <= "0000000000000000";
    ptr_deref_2347_word_offset_1 <= "0000000000000001";
    ptr_deref_2347_word_offset_2 <= "0000000000000010";
    ptr_deref_2347_word_offset_3 <= "0000000000000011";
    ptr_deref_2368_word_offset_0 <= "0000000000000000";
    ptr_deref_2368_word_offset_1 <= "0000000000000001";
    ptr_deref_2368_word_offset_2 <= "0000000000000010";
    ptr_deref_2368_word_offset_3 <= "0000000000000011";
    ptr_deref_2383_word_offset_0 <= "0000000000000000";
    ptr_deref_2383_word_offset_1 <= "0000000000000001";
    ptr_deref_2404_word_offset_0 <= "0000000000000000";
    ptr_deref_2404_word_offset_1 <= "0000000000000001";
    ptr_deref_2404_word_offset_2 <= "0000000000000010";
    ptr_deref_2404_word_offset_3 <= "0000000000000011";
    ptr_deref_2431_word_offset_0 <= "0000000000000000";
    ptr_deref_2431_word_offset_1 <= "0000000000000001";
    ptr_deref_2431_word_offset_2 <= "0000000000000010";
    ptr_deref_2431_word_offset_3 <= "0000000000000011";
    type_cast_2317_wire_constant <= "11111111111111111111100000000000";
    type_cast_2323_wire_constant <= "00000000000000000000000000001000";
    type_cast_2353_wire_constant <= "00000000000000000000000010110100";
    type_cast_2374_wire_constant <= "00000000000000000000000000000110";
    type_cast_2410_wire_constant <= "00000000000000000000011111111111";
    type_cast_2416_wire_constant <= "11111111111111111111111111111000";
    array_obj_ref_2337_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp4_2333, dout => array_obj_ref_2337_resized_base_address, req => array_obj_ref_2337_base_resize_req_0, ack => array_obj_ref_2337_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2337_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2337_root_address, dout => tmp5_2338, req => array_obj_ref_2337_final_reg_req_0, ack => array_obj_ref_2337_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2344_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2329, dout => array_obj_ref_2344_resized_base_address, req => array_obj_ref_2344_base_resize_req_0, ack => array_obj_ref_2344_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2344_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2344_root_address, dout => tmp6_2345, req => array_obj_ref_2344_final_reg_req_0, ack => array_obj_ref_2344_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2365_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2329, dout => array_obj_ref_2365_resized_base_address, req => array_obj_ref_2365_base_resize_req_0, ack => array_obj_ref_2365_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2365_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2365_root_address, dout => tmp9_2366, req => array_obj_ref_2365_final_reg_req_0, ack => array_obj_ref_2365_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2394_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2359, dout => array_obj_ref_2394_resized_base_address, req => array_obj_ref_2394_base_resize_req_0, ack => array_obj_ref_2394_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2394_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2394_root_address, dout => tmp15_2395, req => array_obj_ref_2394_final_reg_req_0, ack => array_obj_ref_2394_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2394_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp14_2391, dout => simple_obj_ref_2393_resized, req => array_obj_ref_2394_index_0_resize_req_0, ack => array_obj_ref_2394_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2394_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_2393_scaled, dout => array_obj_ref_2394_final_offset, req => array_obj_ref_2394_offset_inst_req_0, ack => array_obj_ref_2394_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2401_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2329, dout => array_obj_ref_2401_resized_base_address, req => array_obj_ref_2401_base_resize_req_0, ack => array_obj_ref_2401_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2401_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2401_root_address, dout => tmp16_2402, req => array_obj_ref_2401_final_reg_req_0, ack => array_obj_ref_2401_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2428_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2329, dout => array_obj_ref_2428_resized_base_address, req => array_obj_ref_2428_base_resize_req_0, ack => array_obj_ref_2428_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2428_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2428_root_address, dout => tmp20_2429, req => array_obj_ref_2428_final_reg_req_0, ack => array_obj_ref_2428_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2347_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2345, dout => ptr_deref_2347_resized_base_address, req => ptr_deref_2347_base_resize_req_0, ack => ptr_deref_2347_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2368_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2366, dout => ptr_deref_2368_resized_base_address, req => ptr_deref_2368_base_resize_req_0, ack => ptr_deref_2368_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2383_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp11_2380, dout => ptr_deref_2383_resized_base_address, req => ptr_deref_2383_base_resize_req_0, ack => ptr_deref_2383_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2404_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp16_2402, dout => ptr_deref_2404_resized_base_address, req => ptr_deref_2404_base_resize_req_0, ack => ptr_deref_2404_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2431_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp20_2429, dout => ptr_deref_2431_resized_base_address, req => ptr_deref_2431_base_resize_req_0, ack => ptr_deref_2431_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2312_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2311_wire, dout => tmp_2313, req => type_cast_2312_inst_req_0, ack => type_cast_2312_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2328_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2325, dout => tmp3_2329, req => type_cast_2328_inst_req_0, ack => type_cast_2328_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2332_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2325, dout => tmp4_2333, req => type_cast_2332_inst_req_0, ack => type_cast_2332_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2358_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2355, dout => tmp8_2359, req => type_cast_2358_inst_req_0, ack => type_cast_2358_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2379_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2376, dout => tmp11_2380, req => type_cast_2379_inst_req_0, ack => type_cast_2379_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2390_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2387, dout => tmp14_2391, req => type_cast_2390_inst_req_0, ack => type_cast_2390_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2421_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp18_2418, dout => tmp19_2422, req => type_cast_2421_inst_req_0, ack => type_cast_2421_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2436_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp2_2325, dout => type_cast_2436_wire, req => type_cast_2436_inst_req_0, ack => type_cast_2436_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2394_index_0_rename: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_2394_index_0_rename_ack_0 <= array_obj_ref_2394_index_0_rename_req_0;
      aggregated_sig <= simple_obj_ref_2393_resized;
      simple_obj_ref_2393_scaled <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2347_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2347_gather_scatter_ack_0 <= ptr_deref_2347_gather_scatter_req_0;
      aggregated_sig <= tmp5_2338;
      ptr_deref_2347_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2347_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2347_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2347_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2347_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2347_root_address_inst_ack_0 <= ptr_deref_2347_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2347_resized_base_address;
      ptr_deref_2347_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2368_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2368_gather_scatter_ack_0 <= ptr_deref_2368_gather_scatter_req_0;
      aggregated_sig <= tmp8_2359;
      ptr_deref_2368_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2368_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2368_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2368_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2368_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2368_root_address_inst_ack_0 <= ptr_deref_2368_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2368_resized_base_address;
      ptr_deref_2368_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2383_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2383_gather_scatter_ack_0 <= ptr_deref_2383_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2383_data_1 & ptr_deref_2383_data_0;
      tmp12_2384 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2383_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2383_root_address_inst_ack_0 <= ptr_deref_2383_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2383_resized_base_address;
      ptr_deref_2383_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2404_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2404_gather_scatter_ack_0 <= ptr_deref_2404_gather_scatter_req_0;
      aggregated_sig <= tmp15_2395;
      ptr_deref_2404_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2404_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2404_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2404_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2404_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2404_root_address_inst_ack_0 <= ptr_deref_2404_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2404_resized_base_address;
      ptr_deref_2404_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2431_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2431_gather_scatter_ack_0 <= ptr_deref_2431_gather_scatter_req_0;
      aggregated_sig <= tmp19_2422;
      ptr_deref_2431_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_2431_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_2431_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2431_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2431_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2431_root_address_inst_ack_0 <= ptr_deref_2431_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2431_resized_base_address;
      ptr_deref_2431_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2337_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2337_resized_base_address;
      array_obj_ref_2337_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000001101100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2337_root_address_inst_req_0,
          ackL => array_obj_ref_2337_root_address_inst_ack_0,
          reqR => array_obj_ref_2337_root_address_inst_req_1,
          ackR => array_obj_ref_2337_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2344_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2344_resized_base_address;
      array_obj_ref_2344_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2344_root_address_inst_req_0,
          ackL => array_obj_ref_2344_root_address_inst_ack_0,
          reqR => array_obj_ref_2344_root_address_inst_req_1,
          ackR => array_obj_ref_2344_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_2365_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2365_resized_base_address;
      array_obj_ref_2365_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2365_root_address_inst_req_0,
          ackL => array_obj_ref_2365_root_address_inst_ack_0,
          reqR => array_obj_ref_2365_root_address_inst_req_1,
          ackR => array_obj_ref_2365_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_2394_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2394_final_offset & array_obj_ref_2394_resized_base_address;
      array_obj_ref_2394_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2394_root_address_inst_req_0,
          ackL => array_obj_ref_2394_root_address_inst_ack_0,
          reqR => array_obj_ref_2394_root_address_inst_req_1,
          ackR => array_obj_ref_2394_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : array_obj_ref_2401_root_address_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2401_resized_base_address;
      array_obj_ref_2401_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2401_root_address_inst_req_0,
          ackL => array_obj_ref_2401_root_address_inst_ack_0,
          reqR => array_obj_ref_2401_root_address_inst_req_1,
          ackR => array_obj_ref_2401_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : array_obj_ref_2428_root_address_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2428_resized_base_address;
      array_obj_ref_2428_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2428_root_address_inst_req_0,
          ackL => array_obj_ref_2428_root_address_inst_ack_0,
          reqR => array_obj_ref_2428_root_address_inst_req_1,
          ackR => array_obj_ref_2428_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2318_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2313;
      tmp1_2319 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2318_inst_req_0,
          ackL => binary_2318_inst_ack_0,
          reqR => binary_2318_inst_req_1,
          ackR => binary_2318_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2324_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_2319;
      tmp2_2325 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2324_inst_req_0,
          ackL => binary_2324_inst_ack_0,
          reqR => binary_2324_inst_req_1,
          ackR => binary_2324_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2354_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_2319;
      tmp7_2355 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000010110100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2354_inst_req_0,
          ackL => binary_2354_inst_ack_0,
          reqR => binary_2354_inst_req_1,
          ackR => binary_2354_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2375_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp1_2319;
      tmp10_2376 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2375_inst_req_0,
          ackL => binary_2375_inst_ack_0,
          reqR => binary_2375_inst_req_1,
          ackR => binary_2375_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2411_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2313;
      tmp17_2412 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000011111111111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2411_inst_req_0,
          ackL => binary_2411_inst_ack_0,
          reqR => binary_2411_inst_req_1,
          ackR => binary_2411_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_2417_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp17_2412;
      tmp18_2418 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111111111111000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2417_inst_req_0,
          ackL => binary_2417_inst_ack_0,
          reqR => binary_2417_inst_req_1,
          ackR => binary_2417_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2347_addr_0 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2347_root_address;
      ptr_deref_2347_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2347_addr_0_req_0,
          ackL => ptr_deref_2347_addr_0_ack_0,
          reqR => ptr_deref_2347_addr_0_req_1,
          ackR => ptr_deref_2347_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2347_addr_1 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2347_root_address;
      ptr_deref_2347_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2347_addr_1_req_0,
          ackL => ptr_deref_2347_addr_1_ack_0,
          reqR => ptr_deref_2347_addr_1_req_1,
          ackR => ptr_deref_2347_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2347_addr_2 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2347_root_address;
      ptr_deref_2347_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2347_addr_2_req_0,
          ackL => ptr_deref_2347_addr_2_ack_0,
          reqR => ptr_deref_2347_addr_2_req_1,
          ackR => ptr_deref_2347_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2347_addr_3 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2347_root_address;
      ptr_deref_2347_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2347_addr_3_req_0,
          ackL => ptr_deref_2347_addr_3_ack_0,
          reqR => ptr_deref_2347_addr_3_req_1,
          ackR => ptr_deref_2347_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2368_addr_0 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2368_root_address;
      ptr_deref_2368_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2368_addr_0_req_0,
          ackL => ptr_deref_2368_addr_0_ack_0,
          reqR => ptr_deref_2368_addr_0_req_1,
          ackR => ptr_deref_2368_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2368_addr_1 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2368_root_address;
      ptr_deref_2368_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2368_addr_1_req_0,
          ackL => ptr_deref_2368_addr_1_ack_0,
          reqR => ptr_deref_2368_addr_1_req_1,
          ackR => ptr_deref_2368_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2368_addr_2 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2368_root_address;
      ptr_deref_2368_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2368_addr_2_req_0,
          ackL => ptr_deref_2368_addr_2_ack_0,
          reqR => ptr_deref_2368_addr_2_req_1,
          ackR => ptr_deref_2368_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2368_addr_3 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2368_root_address;
      ptr_deref_2368_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2368_addr_3_req_0,
          ackL => ptr_deref_2368_addr_3_ack_0,
          reqR => ptr_deref_2368_addr_3_req_1,
          ackR => ptr_deref_2368_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2383_addr_0 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2383_root_address;
      ptr_deref_2383_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2383_addr_0_req_0,
          ackL => ptr_deref_2383_addr_0_ack_0,
          reqR => ptr_deref_2383_addr_0_req_1,
          ackR => ptr_deref_2383_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2383_addr_1 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2383_root_address;
      ptr_deref_2383_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2383_addr_1_req_0,
          ackL => ptr_deref_2383_addr_1_ack_0,
          reqR => ptr_deref_2383_addr_1_req_1,
          ackR => ptr_deref_2383_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2404_addr_0 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2404_root_address;
      ptr_deref_2404_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2404_addr_0_req_0,
          ackL => ptr_deref_2404_addr_0_ack_0,
          reqR => ptr_deref_2404_addr_0_req_1,
          ackR => ptr_deref_2404_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2404_addr_1 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2404_root_address;
      ptr_deref_2404_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2404_addr_1_req_0,
          ackL => ptr_deref_2404_addr_1_ack_0,
          reqR => ptr_deref_2404_addr_1_req_1,
          ackR => ptr_deref_2404_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2404_addr_2 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2404_root_address;
      ptr_deref_2404_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2404_addr_2_req_0,
          ackL => ptr_deref_2404_addr_2_ack_0,
          reqR => ptr_deref_2404_addr_2_req_1,
          ackR => ptr_deref_2404_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2404_addr_3 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2404_root_address;
      ptr_deref_2404_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2404_addr_3_req_0,
          ackL => ptr_deref_2404_addr_3_ack_0,
          reqR => ptr_deref_2404_addr_3_req_1,
          ackR => ptr_deref_2404_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2431_addr_0 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2431_root_address;
      ptr_deref_2431_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2431_addr_0_req_0,
          ackL => ptr_deref_2431_addr_0_ack_0,
          reqR => ptr_deref_2431_addr_0_req_1,
          ackR => ptr_deref_2431_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2431_addr_1 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2431_root_address;
      ptr_deref_2431_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2431_addr_1_req_0,
          ackL => ptr_deref_2431_addr_1_ack_0,
          reqR => ptr_deref_2431_addr_1_req_1,
          ackR => ptr_deref_2431_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2431_addr_2 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2431_root_address;
      ptr_deref_2431_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2431_addr_2_req_0,
          ackL => ptr_deref_2431_addr_2_ack_0,
          reqR => ptr_deref_2431_addr_2_req_1,
          ackR => ptr_deref_2431_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : ptr_deref_2431_addr_3 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2431_root_address;
      ptr_deref_2431_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2431_addr_3_req_0,
          ackL => ptr_deref_2431_addr_3_ack_0,
          reqR => ptr_deref_2431_addr_3_req_1,
          ackR => ptr_deref_2431_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared load operator group (0) : ptr_deref_2383_load_0 ptr_deref_2383_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2383_load_0_req_0,
        ptr_deref_2383_load_0_ack_0,
        ptr_deref_2383_load_0_req_1,
        ptr_deref_2383_load_0_ack_1,
        "ptr_deref_2383_load_0",
        "memory_space_5" ,
        ptr_deref_2383_data_0,
        ptr_deref_2383_word_address_0,
        "ptr_deref_2383_data_0",
        "ptr_deref_2383_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2383_load_1_req_0,
        ptr_deref_2383_load_1_ack_0,
        ptr_deref_2383_load_1_req_1,
        ptr_deref_2383_load_1_ack_1,
        "ptr_deref_2383_load_1",
        "memory_space_5" ,
        ptr_deref_2383_data_1,
        ptr_deref_2383_word_address_1,
        "ptr_deref_2383_data_1",
        "ptr_deref_2383_word_address_1" -- 
      );
      reqL(1) <= ptr_deref_2383_load_0_req_0;
      reqL(0) <= ptr_deref_2383_load_1_req_0;
      ptr_deref_2383_load_0_ack_0 <= ackL(1);
      ptr_deref_2383_load_1_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_2383_load_0_req_1;
      reqR(0) <= ptr_deref_2383_load_1_req_1;
      ptr_deref_2383_load_0_ack_1 <= ackR(1);
      ptr_deref_2383_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_2383_word_address_0 & ptr_deref_2383_word_address_1;
      ptr_deref_2383_data_0 <= data_out(15 downto 8);
      ptr_deref_2383_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 2,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 2,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2404_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2404_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2404_word_address_1) &  " data ptr_deref_2404_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2404_data_1) severity note; --
        end if;
        if ptr_deref_2404_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2404_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2404_word_address_2) &  " data ptr_deref_2404_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2404_data_2) severity note; --
        end if;
        if ptr_deref_2431_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2431_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2431_word_address_2) &  " data ptr_deref_2431_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2431_data_2) severity note; --
        end if;
        if ptr_deref_2431_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2431_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2431_word_address_0) &  " data ptr_deref_2431_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2431_data_0) severity note; --
        end if;
        if ptr_deref_2404_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2404_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2404_word_address_0) &  " data ptr_deref_2404_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2404_data_0) severity note; --
        end if;
        if ptr_deref_2404_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2404_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2404_word_address_3) &  " data ptr_deref_2404_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2404_data_3) severity note; --
        end if;
        if ptr_deref_2431_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2431_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2431_word_address_1) &  " data ptr_deref_2431_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2431_data_1) severity note; --
        end if;
        if ptr_deref_2431_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2431_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2431_word_address_3) &  " data ptr_deref_2431_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2431_data_3) severity note; --
        end if;
        if ptr_deref_2347_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2347_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2347_word_address_0) &  " data ptr_deref_2347_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2347_data_0) severity note; --
        end if;
        if ptr_deref_2347_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2347_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2347_word_address_1) &  " data ptr_deref_2347_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2347_data_1) severity note; --
        end if;
        if ptr_deref_2347_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2347_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2347_word_address_2) &  " data ptr_deref_2347_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2347_data_2) severity note; --
        end if;
        if ptr_deref_2347_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2347_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2347_word_address_3) &  " data ptr_deref_2347_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2347_data_3) severity note; --
        end if;
        if ptr_deref_2368_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2368_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2368_word_address_0) &  " data ptr_deref_2368_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2368_data_0) severity note; --
        end if;
        if ptr_deref_2368_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2368_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_2368_word_address_3) &  " data ptr_deref_2368_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_2368_data_3) severity note; --
        end if;
        if ptr_deref_2368_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2368_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2368_word_address_1) &  " data ptr_deref_2368_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2368_data_1) severity note; --
        end if;
        if ptr_deref_2368_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2368_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_2368_word_address_2) &  " data ptr_deref_2368_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_2368_data_2) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2404_store_1 ptr_deref_2404_store_2 ptr_deref_2431_store_2 ptr_deref_2431_store_0 ptr_deref_2404_store_0 ptr_deref_2404_store_3 ptr_deref_2431_store_1 ptr_deref_2431_store_3 ptr_deref_2347_store_0 ptr_deref_2347_store_1 ptr_deref_2347_store_2 ptr_deref_2347_store_3 ptr_deref_2368_store_0 ptr_deref_2368_store_3 ptr_deref_2368_store_1 ptr_deref_2368_store_2 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(255 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 15 downto 0);
      -- 
    begin -- 
      reqL(15) <= ptr_deref_2404_store_1_req_0;
      reqL(14) <= ptr_deref_2404_store_2_req_0;
      reqL(13) <= ptr_deref_2431_store_2_req_0;
      reqL(12) <= ptr_deref_2431_store_0_req_0;
      reqL(11) <= ptr_deref_2404_store_0_req_0;
      reqL(10) <= ptr_deref_2404_store_3_req_0;
      reqL(9) <= ptr_deref_2431_store_1_req_0;
      reqL(8) <= ptr_deref_2431_store_3_req_0;
      reqL(7) <= ptr_deref_2347_store_0_req_0;
      reqL(6) <= ptr_deref_2347_store_1_req_0;
      reqL(5) <= ptr_deref_2347_store_2_req_0;
      reqL(4) <= ptr_deref_2347_store_3_req_0;
      reqL(3) <= ptr_deref_2368_store_0_req_0;
      reqL(2) <= ptr_deref_2368_store_3_req_0;
      reqL(1) <= ptr_deref_2368_store_1_req_0;
      reqL(0) <= ptr_deref_2368_store_2_req_0;
      ptr_deref_2404_store_1_ack_0 <= ackL(15);
      ptr_deref_2404_store_2_ack_0 <= ackL(14);
      ptr_deref_2431_store_2_ack_0 <= ackL(13);
      ptr_deref_2431_store_0_ack_0 <= ackL(12);
      ptr_deref_2404_store_0_ack_0 <= ackL(11);
      ptr_deref_2404_store_3_ack_0 <= ackL(10);
      ptr_deref_2431_store_1_ack_0 <= ackL(9);
      ptr_deref_2431_store_3_ack_0 <= ackL(8);
      ptr_deref_2347_store_0_ack_0 <= ackL(7);
      ptr_deref_2347_store_1_ack_0 <= ackL(6);
      ptr_deref_2347_store_2_ack_0 <= ackL(5);
      ptr_deref_2347_store_3_ack_0 <= ackL(4);
      ptr_deref_2368_store_0_ack_0 <= ackL(3);
      ptr_deref_2368_store_3_ack_0 <= ackL(2);
      ptr_deref_2368_store_1_ack_0 <= ackL(1);
      ptr_deref_2368_store_2_ack_0 <= ackL(0);
      reqR(15) <= ptr_deref_2404_store_1_req_1;
      reqR(14) <= ptr_deref_2404_store_2_req_1;
      reqR(13) <= ptr_deref_2431_store_2_req_1;
      reqR(12) <= ptr_deref_2431_store_0_req_1;
      reqR(11) <= ptr_deref_2404_store_0_req_1;
      reqR(10) <= ptr_deref_2404_store_3_req_1;
      reqR(9) <= ptr_deref_2431_store_1_req_1;
      reqR(8) <= ptr_deref_2431_store_3_req_1;
      reqR(7) <= ptr_deref_2347_store_0_req_1;
      reqR(6) <= ptr_deref_2347_store_1_req_1;
      reqR(5) <= ptr_deref_2347_store_2_req_1;
      reqR(4) <= ptr_deref_2347_store_3_req_1;
      reqR(3) <= ptr_deref_2368_store_0_req_1;
      reqR(2) <= ptr_deref_2368_store_3_req_1;
      reqR(1) <= ptr_deref_2368_store_1_req_1;
      reqR(0) <= ptr_deref_2368_store_2_req_1;
      ptr_deref_2404_store_1_ack_1 <= ackR(15);
      ptr_deref_2404_store_2_ack_1 <= ackR(14);
      ptr_deref_2431_store_2_ack_1 <= ackR(13);
      ptr_deref_2431_store_0_ack_1 <= ackR(12);
      ptr_deref_2404_store_0_ack_1 <= ackR(11);
      ptr_deref_2404_store_3_ack_1 <= ackR(10);
      ptr_deref_2431_store_1_ack_1 <= ackR(9);
      ptr_deref_2431_store_3_ack_1 <= ackR(8);
      ptr_deref_2347_store_0_ack_1 <= ackR(7);
      ptr_deref_2347_store_1_ack_1 <= ackR(6);
      ptr_deref_2347_store_2_ack_1 <= ackR(5);
      ptr_deref_2347_store_3_ack_1 <= ackR(4);
      ptr_deref_2368_store_0_ack_1 <= ackR(3);
      ptr_deref_2368_store_3_ack_1 <= ackR(2);
      ptr_deref_2368_store_1_ack_1 <= ackR(1);
      ptr_deref_2368_store_2_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2404_word_address_1 & ptr_deref_2404_word_address_2 & ptr_deref_2431_word_address_2 & ptr_deref_2431_word_address_0 & ptr_deref_2404_word_address_0 & ptr_deref_2404_word_address_3 & ptr_deref_2431_word_address_1 & ptr_deref_2431_word_address_3 & ptr_deref_2347_word_address_0 & ptr_deref_2347_word_address_1 & ptr_deref_2347_word_address_2 & ptr_deref_2347_word_address_3 & ptr_deref_2368_word_address_0 & ptr_deref_2368_word_address_3 & ptr_deref_2368_word_address_1 & ptr_deref_2368_word_address_2;
      data_in <= ptr_deref_2404_data_1 & ptr_deref_2404_data_2 & ptr_deref_2431_data_2 & ptr_deref_2431_data_0 & ptr_deref_2404_data_0 & ptr_deref_2404_data_3 & ptr_deref_2431_data_1 & ptr_deref_2431_data_3 & ptr_deref_2347_data_0 & ptr_deref_2347_data_1 & ptr_deref_2347_data_2 & ptr_deref_2347_data_3 & ptr_deref_2368_data_0 & ptr_deref_2368_data_3 & ptr_deref_2368_data_1 & ptr_deref_2368_data_2;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 16,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 16,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2311_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2311_inst_ack_0 then -- 
            assert false report " ReadPipe src_in0 to wire simple_obj_ref_2311_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2311_inst_req_0;
      simple_obj_ref_2311_inst_ack_0 <= ack(0);
      simple_obj_ref_2311_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => src_in0_pipe_read_req(0),
          oack => src_in0_pipe_read_ack(0),
          odata => src_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2434_inst_ack_0 then -- 
          assert false report " WritePipe chk_in0 from wire type_cast_2436_wire value="  &  convert_slv_to_hex_string(type_cast_2436_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2434_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2434_inst_req_0;
      simple_obj_ref_2434_inst_ack_0 <= ack(0);
      data_in <= type_cast_2436_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => chk_in0_pipe_write_req(0),
          oack => chk_in0_pipe_write_ack(0),
          odata => chk_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_2387_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_2387_call_req_0;
      call_stmt_2387_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_2387_call_req_1;
      call_stmt_2387_call_ack_1 <= ackR(0);
      data_in <= tmp12_2384;
      tmp13_2387 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 16,
        owidth => 16,
        twidth => 2,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 16, twidth => 2, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to0 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to0_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to0_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to0_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga0_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to0;
architecture Default of ahir_glue_to0 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to0_CP_11804_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_2510_base_resize_req_0 : boolean;
  signal ptr_deref_2514_root_address_inst_req_0 : boolean;
  signal ptr_deref_2514_addr_3_ack_1 : boolean;
  signal type_cast_2503_inst_ack_0 : boolean;
  signal ptr_deref_2514_load_3_ack_0 : boolean;
  signal array_obj_ref_2510_final_reg_req_0 : boolean;
  signal ptr_deref_2514_base_resize_ack_0 : boolean;
  signal ptr_deref_2514_load_1_ack_0 : boolean;
  signal ptr_deref_2514_load_3_req_0 : boolean;
  signal ptr_deref_2514_root_address_inst_ack_0 : boolean;
  signal type_cast_2503_inst_req_0 : boolean;
  signal array_obj_ref_2510_final_reg_ack_0 : boolean;
  signal array_obj_ref_2510_root_address_inst_ack_1 : boolean;
  signal ptr_deref_2514_addr_2_ack_1 : boolean;
  signal ptr_deref_2514_load_1_req_0 : boolean;
  signal array_obj_ref_2510_base_resize_ack_0 : boolean;
  signal array_obj_ref_2510_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2510_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2514_addr_2_req_1 : boolean;
  signal array_obj_ref_2510_root_address_inst_req_0 : boolean;
  signal ptr_deref_2514_load_0_ack_0 : boolean;
  signal ptr_deref_2514_addr_3_req_1 : boolean;
  signal ptr_deref_2514_addr_3_ack_0 : boolean;
  signal ptr_deref_2514_load_0_req_0 : boolean;
  signal ptr_deref_2514_load_2_ack_1 : boolean;
  signal ptr_deref_2514_addr_0_req_0 : boolean;
  signal ptr_deref_2514_addr_0_ack_0 : boolean;
  signal ptr_deref_2514_addr_0_req_1 : boolean;
  signal ptr_deref_2514_addr_0_ack_1 : boolean;
  signal ptr_deref_2514_addr_3_req_0 : boolean;
  signal ptr_deref_2514_addr_1_req_0 : boolean;
  signal ptr_deref_2514_addr_1_ack_0 : boolean;
  signal ptr_deref_2514_addr_1_req_1 : boolean;
  signal ptr_deref_2514_load_2_req_0 : boolean;
  signal ptr_deref_2514_addr_1_ack_1 : boolean;
  signal ptr_deref_2514_load_2_ack_0 : boolean;
  signal ptr_deref_2514_addr_2_req_0 : boolean;
  signal ptr_deref_2514_addr_2_ack_0 : boolean;
  signal ptr_deref_2514_load_0_req_1 : boolean;
  signal ptr_deref_2514_load_0_ack_1 : boolean;
  signal ptr_deref_2514_load_3_ack_1 : boolean;
  signal binary_2523_inst_req_0 : boolean;
  signal binary_2523_inst_ack_0 : boolean;
  signal ptr_deref_2514_load_1_req_1 : boolean;
  signal ptr_deref_2514_load_1_ack_1 : boolean;
  signal ptr_deref_2514_load_2_req_1 : boolean;
  signal ptr_deref_2514_load_3_req_1 : boolean;
  signal ptr_deref_2514_base_resize_req_0 : boolean;
  signal type_cast_2518_inst_req_0 : boolean;
  signal type_cast_2518_inst_ack_0 : boolean;
  signal ptr_deref_2514_gather_scatter_req_0 : boolean;
  signal ptr_deref_2514_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_2445_inst_req_0 : boolean;
  signal simple_obj_ref_2445_inst_ack_0 : boolean;
  signal type_cast_2446_inst_req_0 : boolean;
  signal type_cast_2446_inst_ack_0 : boolean;
  signal type_cast_2450_inst_req_0 : boolean;
  signal type_cast_2450_inst_ack_0 : boolean;
  signal binary_2456_inst_req_0 : boolean;
  signal binary_2456_inst_ack_0 : boolean;
  signal binary_2456_inst_req_1 : boolean;
  signal binary_2456_inst_ack_1 : boolean;
  signal type_cast_2460_inst_req_0 : boolean;
  signal type_cast_2460_inst_ack_0 : boolean;
  signal call_stmt_2465_call_req_0 : boolean;
  signal call_stmt_2465_call_ack_0 : boolean;
  signal call_stmt_2465_call_req_1 : boolean;
  signal call_stmt_2465_call_ack_1 : boolean;
  signal ptr_deref_2467_base_resize_req_0 : boolean;
  signal ptr_deref_2467_base_resize_ack_0 : boolean;
  signal ptr_deref_2467_root_address_inst_req_0 : boolean;
  signal ptr_deref_2467_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2467_addr_0_req_0 : boolean;
  signal ptr_deref_2467_addr_0_ack_0 : boolean;
  signal ptr_deref_2467_addr_0_req_1 : boolean;
  signal ptr_deref_2467_addr_0_ack_1 : boolean;
  signal ptr_deref_2467_addr_1_req_0 : boolean;
  signal ptr_deref_2467_addr_1_ack_0 : boolean;
  signal ptr_deref_2467_addr_1_req_1 : boolean;
  signal ptr_deref_2467_addr_1_ack_1 : boolean;
  signal ptr_deref_2467_gather_scatter_req_0 : boolean;
  signal ptr_deref_2467_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2467_store_0_req_0 : boolean;
  signal ptr_deref_2467_store_0_ack_0 : boolean;
  signal ptr_deref_2467_store_1_req_0 : boolean;
  signal ptr_deref_2467_store_1_ack_0 : boolean;
  signal ptr_deref_2467_store_0_req_1 : boolean;
  signal ptr_deref_2467_store_0_ack_1 : boolean;
  signal ptr_deref_2467_store_1_req_1 : boolean;
  signal ptr_deref_2467_store_1_ack_1 : boolean;
  signal binary_2474_inst_req_0 : boolean;
  signal binary_2474_inst_ack_0 : boolean;
  signal binary_2474_inst_req_1 : boolean;
  signal binary_2474_inst_ack_1 : boolean;
  signal type_cast_2478_inst_req_0 : boolean;
  signal type_cast_2478_inst_ack_0 : boolean;
  signal binary_2484_inst_req_0 : boolean;
  signal binary_2484_inst_ack_0 : boolean;
  signal binary_2484_inst_req_1 : boolean;
  signal binary_2484_inst_ack_1 : boolean;
  signal binary_2523_inst_req_1 : boolean;
  signal binary_2523_inst_ack_1 : boolean;
  signal type_cast_2488_inst_req_0 : boolean;
  signal type_cast_2488_inst_ack_0 : boolean;
  signal array_obj_ref_2495_base_resize_req_0 : boolean;
  signal array_obj_ref_2495_base_resize_ack_0 : boolean;
  signal array_obj_ref_2495_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2495_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2495_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2495_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2495_final_reg_req_0 : boolean;
  signal array_obj_ref_2495_final_reg_ack_0 : boolean;
  signal ptr_deref_2499_base_resize_req_0 : boolean;
  signal ptr_deref_2499_base_resize_ack_0 : boolean;
  signal ptr_deref_2499_root_address_inst_req_0 : boolean;
  signal ptr_deref_2499_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2499_addr_0_req_0 : boolean;
  signal ptr_deref_2499_addr_0_ack_0 : boolean;
  signal ptr_deref_2499_addr_0_req_1 : boolean;
  signal ptr_deref_2499_addr_0_ack_1 : boolean;
  signal ptr_deref_2499_addr_1_req_0 : boolean;
  signal ptr_deref_2499_addr_1_ack_0 : boolean;
  signal ptr_deref_2499_addr_1_req_1 : boolean;
  signal ptr_deref_2499_addr_1_ack_1 : boolean;
  signal ptr_deref_2499_addr_2_req_0 : boolean;
  signal ptr_deref_2499_addr_2_ack_0 : boolean;
  signal ptr_deref_2499_addr_2_req_1 : boolean;
  signal ptr_deref_2499_addr_2_ack_1 : boolean;
  signal ptr_deref_2499_addr_3_req_0 : boolean;
  signal ptr_deref_2499_addr_3_ack_0 : boolean;
  signal ptr_deref_2499_addr_3_req_1 : boolean;
  signal ptr_deref_2499_addr_3_ack_1 : boolean;
  signal ptr_deref_2499_load_0_req_0 : boolean;
  signal ptr_deref_2499_load_0_ack_0 : boolean;
  signal ptr_deref_2499_load_1_req_0 : boolean;
  signal ptr_deref_2499_load_1_ack_0 : boolean;
  signal ptr_deref_2499_load_2_req_0 : boolean;
  signal ptr_deref_2499_load_2_ack_0 : boolean;
  signal ptr_deref_2499_load_3_req_0 : boolean;
  signal ptr_deref_2499_load_3_ack_0 : boolean;
  signal ptr_deref_2499_load_0_req_1 : boolean;
  signal ptr_deref_2499_load_0_ack_1 : boolean;
  signal ptr_deref_2499_load_1_req_1 : boolean;
  signal ptr_deref_2499_load_1_ack_1 : boolean;
  signal ptr_deref_2499_load_2_req_1 : boolean;
  signal ptr_deref_2499_load_2_ack_1 : boolean;
  signal ptr_deref_2499_load_3_req_1 : boolean;
  signal ptr_deref_2499_load_3_ack_1 : boolean;
  signal ptr_deref_2499_gather_scatter_req_0 : boolean;
  signal ptr_deref_2499_gather_scatter_ack_0 : boolean;
  signal type_cast_2527_inst_req_0 : boolean;
  signal type_cast_2527_inst_ack_0 : boolean;
  signal binary_2533_inst_req_0 : boolean;
  signal binary_2533_inst_ack_0 : boolean;
  signal binary_2533_inst_req_1 : boolean;
  signal binary_2533_inst_ack_1 : boolean;
  signal type_cast_2537_inst_req_0 : boolean;
  signal type_cast_2537_inst_ack_0 : boolean;
  signal binary_2543_inst_req_0 : boolean;
  signal binary_2543_inst_ack_0 : boolean;
  signal binary_2543_inst_req_1 : boolean;
  signal binary_2543_inst_ack_1 : boolean;
  signal binary_2549_inst_req_0 : boolean;
  signal binary_2549_inst_ack_0 : boolean;
  signal binary_2549_inst_req_1 : boolean;
  signal binary_2549_inst_ack_1 : boolean;
  signal type_cast_2553_inst_req_0 : boolean;
  signal type_cast_2553_inst_ack_0 : boolean;
  signal binary_2557_inst_req_0 : boolean;
  signal binary_2557_inst_ack_0 : boolean;
  signal binary_2557_inst_req_1 : boolean;
  signal binary_2557_inst_ack_1 : boolean;
  signal type_cast_2561_inst_req_0 : boolean;
  signal type_cast_2561_inst_ack_0 : boolean;
  signal binary_2566_inst_req_0 : boolean;
  signal binary_2566_inst_ack_0 : boolean;
  signal binary_2566_inst_req_1 : boolean;
  signal binary_2566_inst_ack_1 : boolean;
  signal call_stmt_2570_call_req_0 : boolean;
  signal call_stmt_2570_call_ack_0 : boolean;
  signal call_stmt_2570_call_req_1 : boolean;
  signal call_stmt_2570_call_ack_1 : boolean;
  signal ptr_deref_2572_base_resize_req_0 : boolean;
  signal ptr_deref_2572_base_resize_ack_0 : boolean;
  signal ptr_deref_2572_root_address_inst_req_0 : boolean;
  signal ptr_deref_2572_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2572_addr_0_req_0 : boolean;
  signal ptr_deref_2572_addr_0_ack_0 : boolean;
  signal ptr_deref_2572_addr_0_req_1 : boolean;
  signal ptr_deref_2572_addr_0_ack_1 : boolean;
  signal ptr_deref_2572_addr_1_req_0 : boolean;
  signal ptr_deref_2572_addr_1_ack_0 : boolean;
  signal ptr_deref_2572_addr_1_req_1 : boolean;
  signal ptr_deref_2572_addr_1_ack_1 : boolean;
  signal ptr_deref_2572_gather_scatter_req_0 : boolean;
  signal ptr_deref_2572_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2572_store_0_req_0 : boolean;
  signal ptr_deref_2572_store_0_ack_0 : boolean;
  signal ptr_deref_2572_store_1_req_0 : boolean;
  signal ptr_deref_2572_store_1_ack_0 : boolean;
  signal ptr_deref_2572_store_0_req_1 : boolean;
  signal ptr_deref_2572_store_0_ack_1 : boolean;
  signal ptr_deref_2572_store_1_req_1 : boolean;
  signal ptr_deref_2572_store_1_ack_1 : boolean;
  signal call_stmt_2577_call_req_0 : boolean;
  signal call_stmt_2577_call_ack_0 : boolean;
  signal call_stmt_2577_call_req_1 : boolean;
  signal call_stmt_2577_call_ack_1 : boolean;
  signal ptr_deref_2579_base_resize_req_0 : boolean;
  signal ptr_deref_2579_base_resize_ack_0 : boolean;
  signal ptr_deref_2579_root_address_inst_req_0 : boolean;
  signal ptr_deref_2579_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2579_addr_0_req_0 : boolean;
  signal ptr_deref_2579_addr_0_ack_0 : boolean;
  signal ptr_deref_2579_addr_0_req_1 : boolean;
  signal ptr_deref_2579_addr_0_ack_1 : boolean;
  signal ptr_deref_2579_addr_1_req_0 : boolean;
  signal ptr_deref_2579_addr_1_ack_0 : boolean;
  signal ptr_deref_2579_addr_1_req_1 : boolean;
  signal ptr_deref_2579_addr_1_ack_1 : boolean;
  signal ptr_deref_2579_gather_scatter_req_0 : boolean;
  signal ptr_deref_2579_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2579_store_0_req_0 : boolean;
  signal ptr_deref_2579_store_0_ack_0 : boolean;
  signal ptr_deref_2579_store_1_req_0 : boolean;
  signal ptr_deref_2579_store_1_ack_0 : boolean;
  signal ptr_deref_2579_store_0_req_1 : boolean;
  signal ptr_deref_2579_store_0_ack_1 : boolean;
  signal ptr_deref_2579_store_1_req_1 : boolean;
  signal ptr_deref_2579_store_1_ack_1 : boolean;
  signal ptr_deref_2584_base_resize_req_0 : boolean;
  signal ptr_deref_2584_base_resize_ack_0 : boolean;
  signal ptr_deref_2584_root_address_inst_req_0 : boolean;
  signal ptr_deref_2584_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2584_addr_0_req_0 : boolean;
  signal ptr_deref_2584_addr_0_ack_0 : boolean;
  signal ptr_deref_2584_addr_0_req_1 : boolean;
  signal ptr_deref_2584_addr_0_ack_1 : boolean;
  signal ptr_deref_2584_addr_1_req_0 : boolean;
  signal ptr_deref_2584_addr_1_ack_0 : boolean;
  signal ptr_deref_2584_addr_1_req_1 : boolean;
  signal ptr_deref_2584_addr_1_ack_1 : boolean;
  signal ptr_deref_2584_addr_2_req_0 : boolean;
  signal ptr_deref_2584_addr_2_ack_0 : boolean;
  signal ptr_deref_2584_addr_2_req_1 : boolean;
  signal ptr_deref_2584_addr_2_ack_1 : boolean;
  signal ptr_deref_2584_addr_3_req_0 : boolean;
  signal ptr_deref_2584_addr_3_ack_0 : boolean;
  signal ptr_deref_2584_addr_3_req_1 : boolean;
  signal ptr_deref_2584_addr_3_ack_1 : boolean;
  signal ptr_deref_2584_load_0_req_0 : boolean;
  signal ptr_deref_2584_load_0_ack_0 : boolean;
  signal ptr_deref_2584_load_1_req_0 : boolean;
  signal ptr_deref_2584_load_1_ack_0 : boolean;
  signal ptr_deref_2584_load_2_req_0 : boolean;
  signal ptr_deref_2584_load_2_ack_0 : boolean;
  signal ptr_deref_2584_load_3_req_0 : boolean;
  signal ptr_deref_2584_load_3_ack_0 : boolean;
  signal ptr_deref_2584_load_0_req_1 : boolean;
  signal ptr_deref_2584_load_0_ack_1 : boolean;
  signal ptr_deref_2584_load_1_req_1 : boolean;
  signal ptr_deref_2584_load_1_ack_1 : boolean;
  signal ptr_deref_2584_load_2_req_1 : boolean;
  signal ptr_deref_2584_load_2_ack_1 : boolean;
  signal ptr_deref_2584_load_3_req_1 : boolean;
  signal ptr_deref_2584_load_3_ack_1 : boolean;
  signal ptr_deref_2584_gather_scatter_req_0 : boolean;
  signal ptr_deref_2584_gather_scatter_ack_0 : boolean;
  signal type_cast_2588_inst_req_0 : boolean;
  signal type_cast_2588_inst_ack_0 : boolean;
  signal simple_obj_ref_2590_inst_req_0 : boolean;
  signal simple_obj_ref_2590_inst_ack_0 : boolean;
  signal type_cast_2596_inst_req_0 : boolean;
  signal type_cast_2596_inst_ack_0 : boolean;
  signal simple_obj_ref_2594_inst_req_0 : boolean;
  signal simple_obj_ref_2594_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to0_CP_11804: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_11895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2465_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_12420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2570_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_12718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2590_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2446_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_11845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2445_inst_req_0); -- 
    ack_11846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2445_inst_ack_0, ack => cp_elements(8)); -- 
    ack_11851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2446_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2450_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_11864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2450_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11873_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2456_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_11874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2456_inst_ack_0, ack => cp_elements(18)); -- 
    cr_11875_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2456_inst_req_1); -- 
    ca_11876_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2456_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11885_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2460_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_11886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2460_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_11896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2465_call_ack_0, ack => cp_elements(24)); -- 
    ccr_11900_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2465_call_req_1); -- 
    cca_11901_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2465_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_11947_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2467_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_11920_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2467_base_resize_req_0); -- 
    base_resize_ack_11921_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_11925_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2467_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2467_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_11933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2467_addr_0_req_0); -- 
    ra_11934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_11935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2467_addr_0_req_1); -- 
    ca_11936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_11940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2467_addr_1_req_0); -- 
    ra_11941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_11942_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2467_addr_1_req_1); -- 
    ca_11943_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2467_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_11955_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2467_store_0_req_0); -- 
    ra_11956_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_11960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2467_store_1_req_0); -- 
    ra_11961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_11971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2467_store_0_req_1); -- 
    ca_11972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_11976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2467_store_1_req_1); -- 
    ca_11977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2467_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_11986_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2474_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_11987_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2474_inst_ack_0, ack => cp_elements(55)); -- 
    cr_11988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2474_inst_req_1); -- 
    ca_11989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2474_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_11998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2478_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_11999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2478_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2484_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_12009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2484_inst_ack_0, ack => cp_elements(63)); -- 
    cr_12010_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2484_inst_req_1); -- 
    ca_12011_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2484_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2488_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_12021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2488_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2495_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_12032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2495_base_resize_req_0); -- 
    base_resize_ack_12033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_12038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2495_root_address_inst_req_0); -- 
    plus_base_ra_12039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_12040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2495_root_address_inst_req_1); -- 
    plus_base_ca_12041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2495_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2495_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_12059_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2499_base_resize_req_0); -- 
    base_resize_ack_12060_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_12064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2499_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2499_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_12072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2499_addr_0_req_0); -- 
    ra_12073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_12074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2499_addr_0_req_1); -- 
    ca_12075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_12079_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2499_addr_1_req_0); -- 
    ra_12080_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_12081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2499_addr_1_req_1); -- 
    ca_12082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_12086_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2499_addr_2_req_0); -- 
    ra_12087_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_12088_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2499_addr_2_req_1); -- 
    ca_12089_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_12093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2499_addr_3_req_0); -- 
    ra_12094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_12095_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2499_addr_3_req_1); -- 
    ca_12096_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_12106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2499_load_0_req_0); -- 
    ra_12107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_12111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2499_load_1_req_0); -- 
    ra_12112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_12116_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2499_load_2_req_0); -- 
    ra_12117_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_12121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2499_load_3_req_0); -- 
    ra_12122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_12132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2499_load_0_req_1); -- 
    ca_12133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_12137_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2499_load_1_req_1); -- 
    ca_12138_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_12142_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2499_load_2_req_1); -- 
    ca_12143_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_12147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2499_load_3_req_1); -- 
    ca_12148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12149_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2499_gather_scatter_req_0); -- 
    merge_ack_12150_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2499_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2503_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_12160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2503_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2510_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_12171_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2510_base_resize_req_0); -- 
    base_resize_ack_12172_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2510_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_12177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2510_root_address_inst_req_0); -- 
    plus_base_ra_12178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2510_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_12179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2510_root_address_inst_req_1); -- 
    plus_base_ca_12180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2510_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2510_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_12198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2514_base_resize_req_0); -- 
    base_resize_ack_12199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_12203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2514_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2514_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_12211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2514_addr_0_req_0); -- 
    ra_12212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_12213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2514_addr_0_req_1); -- 
    ca_12214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_12218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2514_addr_1_req_0); -- 
    ra_12219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_12220_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2514_addr_1_req_1); -- 
    ca_12221_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_12225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2514_addr_2_req_0); -- 
    ra_12226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_12227_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2514_addr_2_req_1); -- 
    ca_12228_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_12232_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2514_addr_3_req_0); -- 
    ra_12233_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_12234_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2514_addr_3_req_1); -- 
    ca_12235_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_12245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2514_load_0_req_0); -- 
    ra_12246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_12250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2514_load_1_req_0); -- 
    ra_12251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_12255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2514_load_2_req_0); -- 
    ra_12256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_12260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2514_load_3_req_0); -- 
    ra_12261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_12271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2514_load_0_req_1); -- 
    ca_12272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_12276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2514_load_1_req_1); -- 
    ca_12277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_12281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2514_load_2_req_1); -- 
    ca_12282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_12286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2514_load_3_req_1); -- 
    ca_12287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12288_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2514_gather_scatter_req_0); -- 
    merge_ack_12289_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2514_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2518_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_12299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2518_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2523_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_12310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2523_inst_ack_0, ack => cp_elements(162)); -- 
    cr_12311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2523_inst_req_1); -- 
    cp_elements(163) <= binary_2523_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12321_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2527_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_12322_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2527_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2533_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_12332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2533_inst_ack_0, ack => cp_elements(171)); -- 
    cr_12333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2533_inst_req_1); -- 
    ca_12334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2533_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2537_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_12344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2537_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2543_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_12354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2543_inst_ack_0, ack => cp_elements(178)); -- 
    cr_12355_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2543_inst_req_1); -- 
    ca_12356_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2543_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2549_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_12366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2549_inst_ack_0, ack => cp_elements(183)); -- 
    cr_12367_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2549_inst_req_1); -- 
    ca_12368_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2549_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2557_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2553_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_12380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2553_inst_ack_0, ack => cp_elements(189)); -- 
    ra_12385_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2557_inst_ack_0, ack => cp_elements(190)); -- 
    cr_12386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2557_inst_req_1); -- 
    ca_12387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2557_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2561_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_12397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2561_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12407_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2566_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_12408_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2566_inst_ack_0, ack => cp_elements(197)); -- 
    cr_12409_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2566_inst_req_1); -- 
    ca_12410_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2566_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_12421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2570_call_ack_0, ack => cp_elements(200)); -- 
    ccr_12425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2570_call_req_1); -- 
    cca_12426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2570_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_12472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2572_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_12445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2572_base_resize_req_0); -- 
    base_resize_ack_12446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_12450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2572_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2572_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_12458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2572_addr_0_req_0); -- 
    ra_12459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_12460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2572_addr_0_req_1); -- 
    ca_12461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_12465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2572_addr_1_req_0); -- 
    ra_12466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_12467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2572_addr_1_req_1); -- 
    ca_12468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2572_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_12480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2572_store_0_req_0); -- 
    ra_12481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_12485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2572_store_1_req_0); -- 
    ra_12486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_12496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2572_store_0_req_1); -- 
    ca_12497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_12501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2572_store_1_req_1); -- 
    ca_12502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2572_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_12512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2577_call_req_0); -- 
    cra_12513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2577_call_ack_0, ack => cp_elements(227)); -- 
    ccr_12517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2577_call_req_1); -- 
    cca_12518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2577_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_12564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2579_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_12537_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2579_base_resize_req_0); -- 
    base_resize_ack_12538_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_12542_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2579_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2579_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_12550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2579_addr_0_req_0); -- 
    ra_12551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_12552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2579_addr_0_req_1); -- 
    ca_12553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_12557_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2579_addr_1_req_0); -- 
    ra_12558_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_12559_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2579_addr_1_req_1); -- 
    ca_12560_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2579_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_12572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2579_store_0_req_0); -- 
    ra_12573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_12577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2579_store_1_req_0); -- 
    ra_12578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_12588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2579_store_0_req_1); -- 
    ca_12589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_12593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2579_store_1_req_1); -- 
    ca_12594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2579_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_12607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2584_base_resize_req_0); -- 
    base_resize_ack_12608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_12612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2584_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2584_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_12620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2584_addr_0_req_0); -- 
    ra_12621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_12622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2584_addr_0_req_1); -- 
    ca_12623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_12627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2584_addr_1_req_0); -- 
    ra_12628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_12629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2584_addr_1_req_1); -- 
    ca_12630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_12634_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2584_addr_2_req_0); -- 
    ra_12635_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_12636_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2584_addr_2_req_1); -- 
    ca_12637_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_12641_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2584_addr_3_req_0); -- 
    ra_12642_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_12643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2584_addr_3_req_1); -- 
    ca_12644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_12654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2584_load_0_req_0); -- 
    ra_12655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_12659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2584_load_1_req_0); -- 
    ra_12660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_12664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2584_load_2_req_0); -- 
    ra_12665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_12669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2584_load_3_req_0); -- 
    ra_12670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_12680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2584_load_0_req_1); -- 
    ca_12681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_12685_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2584_load_1_req_1); -- 
    ca_12686_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_12690_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2584_load_2_req_1); -- 
    ca_12691_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_12695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2584_load_3_req_1); -- 
    ca_12696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_12697_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2584_gather_scatter_req_0); -- 
    merge_ack_12698_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2584_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2588_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_12708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2588_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_12719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2590_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2596_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_12732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2596_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_12737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2594_inst_req_0); -- 
    pipe_wack_12738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2594_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2495_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2495_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2495_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2510_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2510_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2510_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2558 : std_logic_vector(0 downto 0);
    signal ptr_deref_2467_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2467_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2467_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2467_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2499_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2499_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2499_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2499_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2499_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2514_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2514_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2514_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2514_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2514_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2572_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2572_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2572_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2579_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2579_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2579_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2584_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2584_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2584_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2584_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2584_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2445_wire : std_logic_vector(31 downto 0);
    signal tmp10_2500 : std_logic_vector(31 downto 0);
    signal tmp11_2504 : std_logic_vector(31 downto 0);
    signal tmp12_2511 : std_logic_vector(31 downto 0);
    signal tmp13_2515 : std_logic_vector(31 downto 0);
    signal tmp14_2519 : std_logic_vector(31 downto 0);
    signal tmp15_2524 : std_logic_vector(31 downto 0);
    signal tmp16_2528 : std_logic_vector(15 downto 0);
    signal tmp17_2534 : std_logic_vector(31 downto 0);
    signal tmp18_2544 : std_logic_vector(15 downto 0);
    signal tmp19_2550 : std_logic_vector(31 downto 0);
    signal tmp1_2451 : std_logic_vector(31 downto 0);
    signal tmp20_2562 : std_logic_vector(15 downto 0);
    signal tmp21_2567 : std_logic_vector(15 downto 0);
    signal tmp22_2570 : std_logic_vector(15 downto 0);
    signal tmp23_2577 : std_logic_vector(15 downto 0);
    signal tmp24_2585 : std_logic_vector(31 downto 0);
    signal tmp25_2589 : std_logic_vector(31 downto 0);
    signal tmp2_2457 : std_logic_vector(31 downto 0);
    signal tmp3_2461 : std_logic_vector(31 downto 0);
    signal tmp4_2465 : std_logic_vector(15 downto 0);
    signal tmp5_2475 : std_logic_vector(31 downto 0);
    signal tmp6_2479 : std_logic_vector(31 downto 0);
    signal tmp7_2485 : std_logic_vector(31 downto 0);
    signal tmp8_2489 : std_logic_vector(31 downto 0);
    signal tmp9_2496 : std_logic_vector(31 downto 0);
    signal tmp_2447 : std_logic_vector(31 downto 0);
    signal type_cast_2455_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2463_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2473_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2532_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2542_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2548_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2553_wire : std_logic_vector(31 downto 0);
    signal type_cast_2556_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2592_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2596_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2538 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2495_final_offset <= "0000000000010000";
    array_obj_ref_2510_final_offset <= "0000000000001100";
    ptr_deref_2467_word_offset_0 <= "0000000000000000";
    ptr_deref_2467_word_offset_1 <= "0000000000000001";
    ptr_deref_2499_word_offset_0 <= "0000000000000000";
    ptr_deref_2499_word_offset_1 <= "0000000000000001";
    ptr_deref_2499_word_offset_2 <= "0000000000000010";
    ptr_deref_2499_word_offset_3 <= "0000000000000011";
    ptr_deref_2514_word_offset_0 <= "0000000000000000";
    ptr_deref_2514_word_offset_1 <= "0000000000000001";
    ptr_deref_2514_word_offset_2 <= "0000000000000010";
    ptr_deref_2514_word_offset_3 <= "0000000000000011";
    ptr_deref_2572_word_offset_0 <= "0000000000000000";
    ptr_deref_2572_word_offset_1 <= "0000000000000001";
    ptr_deref_2579_word_offset_0 <= "0000000000000000";
    ptr_deref_2579_word_offset_1 <= "0000000000000001";
    ptr_deref_2584_word_offset_0 <= "0000000000000000";
    ptr_deref_2584_word_offset_1 <= "0000000000000001";
    ptr_deref_2584_word_offset_2 <= "0000000000000010";
    ptr_deref_2584_word_offset_3 <= "0000000000000011";
    type_cast_2455_wire_constant <= "11111111111111111111100000000000";
    type_cast_2463_wire_constant <= "0000000000000001";
    type_cast_2473_wire_constant <= "00000000000000000000000000000110";
    type_cast_2483_wire_constant <= "00000000000000000000000000000010";
    type_cast_2532_wire_constant <= "00000000000000000000000000000011";
    type_cast_2542_wire_constant <= "0001111111111111";
    type_cast_2548_wire_constant <= "00000000000000000000000000000111";
    type_cast_2556_wire_constant <= "00000000000000000000000000000000";
    type_cast_2592_wire_constant <= "00000000000000000000000000000001";
    array_obj_ref_2495_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2451, dout => array_obj_ref_2495_resized_base_address, req => array_obj_ref_2495_base_resize_req_0, ack => array_obj_ref_2495_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2495_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2495_root_address, dout => tmp9_2496, req => array_obj_ref_2495_final_reg_req_0, ack => array_obj_ref_2495_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2510_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2451, dout => array_obj_ref_2510_resized_base_address, req => array_obj_ref_2510_base_resize_req_0, ack => array_obj_ref_2510_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2510_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2510_root_address, dout => tmp12_2511, req => array_obj_ref_2510_final_reg_req_0, ack => array_obj_ref_2510_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2467_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2461, dout => ptr_deref_2467_resized_base_address, req => ptr_deref_2467_base_resize_req_0, ack => ptr_deref_2467_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2499_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2496, dout => ptr_deref_2499_resized_base_address, req => ptr_deref_2499_base_resize_req_0, ack => ptr_deref_2499_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2514_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2511, dout => ptr_deref_2514_resized_base_address, req => ptr_deref_2514_base_resize_req_0, ack => ptr_deref_2514_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2572_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2479, dout => ptr_deref_2572_resized_base_address, req => ptr_deref_2572_base_resize_req_0, ack => ptr_deref_2572_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2579_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2489, dout => ptr_deref_2579_resized_base_address, req => ptr_deref_2579_base_resize_req_0, ack => ptr_deref_2579_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2584_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2511, dout => ptr_deref_2584_resized_base_address, req => ptr_deref_2584_base_resize_req_0, ack => ptr_deref_2584_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2446_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2445_wire, dout => tmp_2447, req => type_cast_2446_inst_req_0, ack => type_cast_2446_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2450_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2447, dout => tmp1_2451, req => type_cast_2450_inst_req_0, ack => type_cast_2450_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2460_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2457, dout => tmp3_2461, req => type_cast_2460_inst_req_0, ack => type_cast_2460_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2478_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2475, dout => tmp6_2479, req => type_cast_2478_inst_req_0, ack => type_cast_2478_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2488_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2485, dout => tmp8_2489, req => type_cast_2488_inst_req_0, ack => type_cast_2488_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2503_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2500, dout => tmp11_2504, req => type_cast_2503_inst_req_0, ack => type_cast_2503_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2518_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2515, dout => tmp14_2519, req => type_cast_2518_inst_req_0, ack => type_cast_2518_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2527_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2524, dout => tmp16_2528, req => type_cast_2527_inst_req_0, ack => type_cast_2527_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2537_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2534, dout => xx_xtrx_xi_2538, req => type_cast_2537_inst_req_0, ack => type_cast_2537_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2553_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2550, dout => type_cast_2553_wire, req => type_cast_2553_inst_req_0, ack => type_cast_2553_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2561_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2558, dout => tmp20_2562, req => type_cast_2561_inst_req_0, ack => type_cast_2561_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2588_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2585, dout => tmp25_2589, req => type_cast_2588_inst_req_0, ack => type_cast_2588_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2596_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2589, dout => type_cast_2596_wire, req => type_cast_2596_inst_req_0, ack => type_cast_2596_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2467_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2467_gather_scatter_ack_0 <= ptr_deref_2467_gather_scatter_req_0;
      aggregated_sig <= tmp4_2465;
      ptr_deref_2467_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2467_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2467_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2467_root_address_inst_ack_0 <= ptr_deref_2467_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2467_resized_base_address;
      ptr_deref_2467_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2499_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2499_gather_scatter_ack_0 <= ptr_deref_2499_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2499_data_3 & ptr_deref_2499_data_2 & ptr_deref_2499_data_1 & ptr_deref_2499_data_0;
      tmp10_2500 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2499_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2499_root_address_inst_ack_0 <= ptr_deref_2499_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2499_resized_base_address;
      ptr_deref_2499_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2514_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2514_gather_scatter_ack_0 <= ptr_deref_2514_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2514_data_3 & ptr_deref_2514_data_2 & ptr_deref_2514_data_1 & ptr_deref_2514_data_0;
      tmp13_2515 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2514_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2514_root_address_inst_ack_0 <= ptr_deref_2514_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2514_resized_base_address;
      ptr_deref_2514_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2572_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2572_gather_scatter_ack_0 <= ptr_deref_2572_gather_scatter_req_0;
      aggregated_sig <= tmp22_2570;
      ptr_deref_2572_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2572_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2572_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2572_root_address_inst_ack_0 <= ptr_deref_2572_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2572_resized_base_address;
      ptr_deref_2572_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2579_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2579_gather_scatter_ack_0 <= ptr_deref_2579_gather_scatter_req_0;
      aggregated_sig <= tmp23_2577;
      ptr_deref_2579_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2579_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2579_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2579_root_address_inst_ack_0 <= ptr_deref_2579_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2579_resized_base_address;
      ptr_deref_2579_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2584_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2584_gather_scatter_ack_0 <= ptr_deref_2584_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2584_data_3 & ptr_deref_2584_data_2 & ptr_deref_2584_data_1 & ptr_deref_2584_data_0;
      tmp24_2585 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2584_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2584_root_address_inst_ack_0 <= ptr_deref_2584_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2584_resized_base_address;
      ptr_deref_2584_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2495_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2495_resized_base_address;
      array_obj_ref_2495_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2495_root_address_inst_req_0,
          ackL => array_obj_ref_2495_root_address_inst_ack_0,
          reqR => array_obj_ref_2495_root_address_inst_req_1,
          ackR => array_obj_ref_2495_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2510_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2510_resized_base_address;
      array_obj_ref_2510_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2510_root_address_inst_req_0,
          ackL => array_obj_ref_2510_root_address_inst_ack_0,
          reqR => array_obj_ref_2510_root_address_inst_req_1,
          ackR => array_obj_ref_2510_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2456_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2447;
      tmp2_2457 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2456_inst_req_0,
          ackL => binary_2456_inst_ack_0,
          reqR => binary_2456_inst_req_1,
          ackR => binary_2456_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2474_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2457;
      tmp5_2475 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2474_inst_req_0,
          ackL => binary_2474_inst_ack_0,
          reqR => binary_2474_inst_req_1,
          ackR => binary_2474_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2484_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2457;
      tmp7_2485 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2484_inst_req_0,
          ackL => binary_2484_inst_ack_0,
          reqR => binary_2484_inst_req_1,
          ackR => binary_2484_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2523_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2504 & tmp14_2519;
      tmp15_2524 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2523_inst_req_0,
          ackL => binary_2523_inst_ack_0,
          reqR => binary_2523_inst_req_1,
          ackR => binary_2523_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2533_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2524;
      tmp17_2534 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2533_inst_req_0,
          ackL => binary_2533_inst_ack_0,
          reqR => binary_2533_inst_req_1,
          ackR => binary_2533_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2543_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2538;
      tmp18_2544 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2543_inst_req_0,
          ackL => binary_2543_inst_ack_0,
          reqR => binary_2543_inst_req_1,
          ackR => binary_2543_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2549_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2524;
      tmp19_2550 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2549_inst_req_0,
          ackL => binary_2549_inst_ack_0,
          reqR => binary_2549_inst_req_1,
          ackR => binary_2549_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2557_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2553_wire;
      notx_xx_xi_2558 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2557_inst_req_0,
          ackL => binary_2557_inst_ack_0,
          reqR => binary_2557_inst_req_1,
          ackR => binary_2557_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2566_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2544 & tmp20_2562;
      tmp21_2567 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2566_inst_req_0,
          ackL => binary_2566_inst_ack_0,
          reqR => binary_2566_inst_req_1,
          ackR => binary_2566_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2467_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2467_root_address;
      ptr_deref_2467_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2467_addr_0_req_0,
          ackL => ptr_deref_2467_addr_0_ack_0,
          reqR => ptr_deref_2467_addr_0_req_1,
          ackR => ptr_deref_2467_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2467_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2467_root_address;
      ptr_deref_2467_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2467_addr_1_req_0,
          ackL => ptr_deref_2467_addr_1_ack_0,
          reqR => ptr_deref_2467_addr_1_req_1,
          ackR => ptr_deref_2467_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2499_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2499_root_address;
      ptr_deref_2499_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2499_addr_0_req_0,
          ackL => ptr_deref_2499_addr_0_ack_0,
          reqR => ptr_deref_2499_addr_0_req_1,
          ackR => ptr_deref_2499_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2499_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2499_root_address;
      ptr_deref_2499_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2499_addr_1_req_0,
          ackL => ptr_deref_2499_addr_1_ack_0,
          reqR => ptr_deref_2499_addr_1_req_1,
          ackR => ptr_deref_2499_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2499_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2499_root_address;
      ptr_deref_2499_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2499_addr_2_req_0,
          ackL => ptr_deref_2499_addr_2_ack_0,
          reqR => ptr_deref_2499_addr_2_req_1,
          ackR => ptr_deref_2499_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2499_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2499_root_address;
      ptr_deref_2499_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2499_addr_3_req_0,
          ackL => ptr_deref_2499_addr_3_ack_0,
          reqR => ptr_deref_2499_addr_3_req_1,
          ackR => ptr_deref_2499_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2514_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2514_root_address;
      ptr_deref_2514_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2514_addr_0_req_0,
          ackL => ptr_deref_2514_addr_0_ack_0,
          reqR => ptr_deref_2514_addr_0_req_1,
          ackR => ptr_deref_2514_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2514_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2514_root_address;
      ptr_deref_2514_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2514_addr_1_req_0,
          ackL => ptr_deref_2514_addr_1_ack_0,
          reqR => ptr_deref_2514_addr_1_req_1,
          ackR => ptr_deref_2514_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2514_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2514_root_address;
      ptr_deref_2514_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2514_addr_2_req_0,
          ackL => ptr_deref_2514_addr_2_ack_0,
          reqR => ptr_deref_2514_addr_2_req_1,
          ackR => ptr_deref_2514_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2514_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2514_root_address;
      ptr_deref_2514_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2514_addr_3_req_0,
          ackL => ptr_deref_2514_addr_3_ack_0,
          reqR => ptr_deref_2514_addr_3_req_1,
          ackR => ptr_deref_2514_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2572_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2572_root_address;
      ptr_deref_2572_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2572_addr_0_req_0,
          ackL => ptr_deref_2572_addr_0_ack_0,
          reqR => ptr_deref_2572_addr_0_req_1,
          ackR => ptr_deref_2572_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2572_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2572_root_address;
      ptr_deref_2572_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2572_addr_1_req_0,
          ackL => ptr_deref_2572_addr_1_ack_0,
          reqR => ptr_deref_2572_addr_1_req_1,
          ackR => ptr_deref_2572_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2579_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2579_root_address;
      ptr_deref_2579_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2579_addr_0_req_0,
          ackL => ptr_deref_2579_addr_0_ack_0,
          reqR => ptr_deref_2579_addr_0_req_1,
          ackR => ptr_deref_2579_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2579_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2579_root_address;
      ptr_deref_2579_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2579_addr_1_req_0,
          ackL => ptr_deref_2579_addr_1_ack_0,
          reqR => ptr_deref_2579_addr_1_req_1,
          ackR => ptr_deref_2579_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2584_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2584_root_address;
      ptr_deref_2584_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2584_addr_0_req_0,
          ackL => ptr_deref_2584_addr_0_ack_0,
          reqR => ptr_deref_2584_addr_0_req_1,
          ackR => ptr_deref_2584_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2584_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2584_root_address;
      ptr_deref_2584_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2584_addr_1_req_0,
          ackL => ptr_deref_2584_addr_1_ack_0,
          reqR => ptr_deref_2584_addr_1_req_1,
          ackR => ptr_deref_2584_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2584_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2584_root_address;
      ptr_deref_2584_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2584_addr_2_req_0,
          ackL => ptr_deref_2584_addr_2_ack_0,
          reqR => ptr_deref_2584_addr_2_req_1,
          ackR => ptr_deref_2584_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2584_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2584_root_address;
      ptr_deref_2584_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2584_addr_3_req_0,
          ackL => ptr_deref_2584_addr_3_ack_0,
          reqR => ptr_deref_2584_addr_3_req_1,
          ackR => ptr_deref_2584_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2499_load_0 ptr_deref_2584_load_1 ptr_deref_2499_load_3 ptr_deref_2499_load_2 ptr_deref_2584_load_2 ptr_deref_2584_load_3 ptr_deref_2499_load_1 ptr_deref_2514_load_0 ptr_deref_2514_load_1 ptr_deref_2514_load_2 ptr_deref_2514_load_3 ptr_deref_2584_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2499_load_0_req_0,
        ptr_deref_2499_load_0_ack_0,
        ptr_deref_2499_load_0_req_1,
        ptr_deref_2499_load_0_ack_1,
        "ptr_deref_2499_load_0",
        "memory_space_5" ,
        ptr_deref_2499_data_0,
        ptr_deref_2499_word_address_0,
        "ptr_deref_2499_data_0",
        "ptr_deref_2499_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2584_load_1_req_0,
        ptr_deref_2584_load_1_ack_0,
        ptr_deref_2584_load_1_req_1,
        ptr_deref_2584_load_1_ack_1,
        "ptr_deref_2584_load_1",
        "memory_space_5" ,
        ptr_deref_2584_data_1,
        ptr_deref_2584_word_address_1,
        "ptr_deref_2584_data_1",
        "ptr_deref_2584_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2499_load_3_req_0,
        ptr_deref_2499_load_3_ack_0,
        ptr_deref_2499_load_3_req_1,
        ptr_deref_2499_load_3_ack_1,
        "ptr_deref_2499_load_3",
        "memory_space_5" ,
        ptr_deref_2499_data_3,
        ptr_deref_2499_word_address_3,
        "ptr_deref_2499_data_3",
        "ptr_deref_2499_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2499_load_2_req_0,
        ptr_deref_2499_load_2_ack_0,
        ptr_deref_2499_load_2_req_1,
        ptr_deref_2499_load_2_ack_1,
        "ptr_deref_2499_load_2",
        "memory_space_5" ,
        ptr_deref_2499_data_2,
        ptr_deref_2499_word_address_2,
        "ptr_deref_2499_data_2",
        "ptr_deref_2499_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2584_load_2_req_0,
        ptr_deref_2584_load_2_ack_0,
        ptr_deref_2584_load_2_req_1,
        ptr_deref_2584_load_2_ack_1,
        "ptr_deref_2584_load_2",
        "memory_space_5" ,
        ptr_deref_2584_data_2,
        ptr_deref_2584_word_address_2,
        "ptr_deref_2584_data_2",
        "ptr_deref_2584_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2584_load_3_req_0,
        ptr_deref_2584_load_3_ack_0,
        ptr_deref_2584_load_3_req_1,
        ptr_deref_2584_load_3_ack_1,
        "ptr_deref_2584_load_3",
        "memory_space_5" ,
        ptr_deref_2584_data_3,
        ptr_deref_2584_word_address_3,
        "ptr_deref_2584_data_3",
        "ptr_deref_2584_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2499_load_1_req_0,
        ptr_deref_2499_load_1_ack_0,
        ptr_deref_2499_load_1_req_1,
        ptr_deref_2499_load_1_ack_1,
        "ptr_deref_2499_load_1",
        "memory_space_5" ,
        ptr_deref_2499_data_1,
        ptr_deref_2499_word_address_1,
        "ptr_deref_2499_data_1",
        "ptr_deref_2499_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2514_load_0_req_0,
        ptr_deref_2514_load_0_ack_0,
        ptr_deref_2514_load_0_req_1,
        ptr_deref_2514_load_0_ack_1,
        "ptr_deref_2514_load_0",
        "memory_space_5" ,
        ptr_deref_2514_data_0,
        ptr_deref_2514_word_address_0,
        "ptr_deref_2514_data_0",
        "ptr_deref_2514_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2514_load_1_req_0,
        ptr_deref_2514_load_1_ack_0,
        ptr_deref_2514_load_1_req_1,
        ptr_deref_2514_load_1_ack_1,
        "ptr_deref_2514_load_1",
        "memory_space_5" ,
        ptr_deref_2514_data_1,
        ptr_deref_2514_word_address_1,
        "ptr_deref_2514_data_1",
        "ptr_deref_2514_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2514_load_2_req_0,
        ptr_deref_2514_load_2_ack_0,
        ptr_deref_2514_load_2_req_1,
        ptr_deref_2514_load_2_ack_1,
        "ptr_deref_2514_load_2",
        "memory_space_5" ,
        ptr_deref_2514_data_2,
        ptr_deref_2514_word_address_2,
        "ptr_deref_2514_data_2",
        "ptr_deref_2514_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2514_load_3_req_0,
        ptr_deref_2514_load_3_ack_0,
        ptr_deref_2514_load_3_req_1,
        ptr_deref_2514_load_3_ack_1,
        "ptr_deref_2514_load_3",
        "memory_space_5" ,
        ptr_deref_2514_data_3,
        ptr_deref_2514_word_address_3,
        "ptr_deref_2514_data_3",
        "ptr_deref_2514_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2584_load_0_req_0,
        ptr_deref_2584_load_0_ack_0,
        ptr_deref_2584_load_0_req_1,
        ptr_deref_2584_load_0_ack_1,
        "ptr_deref_2584_load_0",
        "memory_space_5" ,
        ptr_deref_2584_data_0,
        ptr_deref_2584_word_address_0,
        "ptr_deref_2584_data_0",
        "ptr_deref_2584_word_address_0" -- 
      );
      reqL(11) <= ptr_deref_2499_load_0_req_0;
      reqL(10) <= ptr_deref_2584_load_1_req_0;
      reqL(9) <= ptr_deref_2499_load_3_req_0;
      reqL(8) <= ptr_deref_2499_load_2_req_0;
      reqL(7) <= ptr_deref_2584_load_2_req_0;
      reqL(6) <= ptr_deref_2584_load_3_req_0;
      reqL(5) <= ptr_deref_2499_load_1_req_0;
      reqL(4) <= ptr_deref_2514_load_0_req_0;
      reqL(3) <= ptr_deref_2514_load_1_req_0;
      reqL(2) <= ptr_deref_2514_load_2_req_0;
      reqL(1) <= ptr_deref_2514_load_3_req_0;
      reqL(0) <= ptr_deref_2584_load_0_req_0;
      ptr_deref_2499_load_0_ack_0 <= ackL(11);
      ptr_deref_2584_load_1_ack_0 <= ackL(10);
      ptr_deref_2499_load_3_ack_0 <= ackL(9);
      ptr_deref_2499_load_2_ack_0 <= ackL(8);
      ptr_deref_2584_load_2_ack_0 <= ackL(7);
      ptr_deref_2584_load_3_ack_0 <= ackL(6);
      ptr_deref_2499_load_1_ack_0 <= ackL(5);
      ptr_deref_2514_load_0_ack_0 <= ackL(4);
      ptr_deref_2514_load_1_ack_0 <= ackL(3);
      ptr_deref_2514_load_2_ack_0 <= ackL(2);
      ptr_deref_2514_load_3_ack_0 <= ackL(1);
      ptr_deref_2584_load_0_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2499_load_0_req_1;
      reqR(10) <= ptr_deref_2584_load_1_req_1;
      reqR(9) <= ptr_deref_2499_load_3_req_1;
      reqR(8) <= ptr_deref_2499_load_2_req_1;
      reqR(7) <= ptr_deref_2584_load_2_req_1;
      reqR(6) <= ptr_deref_2584_load_3_req_1;
      reqR(5) <= ptr_deref_2499_load_1_req_1;
      reqR(4) <= ptr_deref_2514_load_0_req_1;
      reqR(3) <= ptr_deref_2514_load_1_req_1;
      reqR(2) <= ptr_deref_2514_load_2_req_1;
      reqR(1) <= ptr_deref_2514_load_3_req_1;
      reqR(0) <= ptr_deref_2584_load_0_req_1;
      ptr_deref_2499_load_0_ack_1 <= ackR(11);
      ptr_deref_2584_load_1_ack_1 <= ackR(10);
      ptr_deref_2499_load_3_ack_1 <= ackR(9);
      ptr_deref_2499_load_2_ack_1 <= ackR(8);
      ptr_deref_2584_load_2_ack_1 <= ackR(7);
      ptr_deref_2584_load_3_ack_1 <= ackR(6);
      ptr_deref_2499_load_1_ack_1 <= ackR(5);
      ptr_deref_2514_load_0_ack_1 <= ackR(4);
      ptr_deref_2514_load_1_ack_1 <= ackR(3);
      ptr_deref_2514_load_2_ack_1 <= ackR(2);
      ptr_deref_2514_load_3_ack_1 <= ackR(1);
      ptr_deref_2584_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_2499_word_address_0 & ptr_deref_2584_word_address_1 & ptr_deref_2499_word_address_3 & ptr_deref_2499_word_address_2 & ptr_deref_2584_word_address_2 & ptr_deref_2584_word_address_3 & ptr_deref_2499_word_address_1 & ptr_deref_2514_word_address_0 & ptr_deref_2514_word_address_1 & ptr_deref_2514_word_address_2 & ptr_deref_2514_word_address_3 & ptr_deref_2584_word_address_0;
      ptr_deref_2499_data_0 <= data_out(95 downto 88);
      ptr_deref_2584_data_1 <= data_out(87 downto 80);
      ptr_deref_2499_data_3 <= data_out(79 downto 72);
      ptr_deref_2499_data_2 <= data_out(71 downto 64);
      ptr_deref_2584_data_2 <= data_out(63 downto 56);
      ptr_deref_2584_data_3 <= data_out(55 downto 48);
      ptr_deref_2499_data_1 <= data_out(47 downto 40);
      ptr_deref_2514_data_0 <= data_out(39 downto 32);
      ptr_deref_2514_data_1 <= data_out(31 downto 24);
      ptr_deref_2514_data_2 <= data_out(23 downto 16);
      ptr_deref_2514_data_3 <= data_out(15 downto 8);
      ptr_deref_2584_data_0 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2579_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2579_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2579_word_address_1) &  " data ptr_deref_2579_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2579_data_1) severity note; --
        end if;
        if ptr_deref_2467_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2467_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2467_word_address_0) &  " data ptr_deref_2467_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2467_data_0) severity note; --
        end if;
        if ptr_deref_2572_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2572_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2572_word_address_0) &  " data ptr_deref_2572_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2572_data_0) severity note; --
        end if;
        if ptr_deref_2467_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2467_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2467_word_address_1) &  " data ptr_deref_2467_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2467_data_1) severity note; --
        end if;
        if ptr_deref_2572_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2572_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2572_word_address_1) &  " data ptr_deref_2572_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2572_data_1) severity note; --
        end if;
        if ptr_deref_2579_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2579_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2579_word_address_0) &  " data ptr_deref_2579_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2579_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2579_store_1 ptr_deref_2467_store_0 ptr_deref_2572_store_0 ptr_deref_2467_store_1 ptr_deref_2572_store_1 ptr_deref_2579_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2579_store_1_req_0;
      reqL(4) <= ptr_deref_2467_store_0_req_0;
      reqL(3) <= ptr_deref_2572_store_0_req_0;
      reqL(2) <= ptr_deref_2467_store_1_req_0;
      reqL(1) <= ptr_deref_2572_store_1_req_0;
      reqL(0) <= ptr_deref_2579_store_0_req_0;
      ptr_deref_2579_store_1_ack_0 <= ackL(5);
      ptr_deref_2467_store_0_ack_0 <= ackL(4);
      ptr_deref_2572_store_0_ack_0 <= ackL(3);
      ptr_deref_2467_store_1_ack_0 <= ackL(2);
      ptr_deref_2572_store_1_ack_0 <= ackL(1);
      ptr_deref_2579_store_0_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2579_store_1_req_1;
      reqR(4) <= ptr_deref_2467_store_0_req_1;
      reqR(3) <= ptr_deref_2572_store_0_req_1;
      reqR(2) <= ptr_deref_2467_store_1_req_1;
      reqR(1) <= ptr_deref_2572_store_1_req_1;
      reqR(0) <= ptr_deref_2579_store_0_req_1;
      ptr_deref_2579_store_1_ack_1 <= ackR(5);
      ptr_deref_2467_store_0_ack_1 <= ackR(4);
      ptr_deref_2572_store_0_ack_1 <= ackR(3);
      ptr_deref_2467_store_1_ack_1 <= ackR(2);
      ptr_deref_2572_store_1_ack_1 <= ackR(1);
      ptr_deref_2579_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2579_word_address_1 & ptr_deref_2467_word_address_0 & ptr_deref_2572_word_address_0 & ptr_deref_2467_word_address_1 & ptr_deref_2572_word_address_1 & ptr_deref_2579_word_address_0;
      data_in <= ptr_deref_2579_data_1 & ptr_deref_2467_data_0 & ptr_deref_2572_data_0 & ptr_deref_2467_data_1 & ptr_deref_2572_data_1 & ptr_deref_2579_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2445_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2445_inst_ack_0 then -- 
            assert false report " ReadPipe to0_in0 to wire simple_obj_ref_2445_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2445_inst_req_0;
      simple_obj_ref_2445_inst_ack_0 <= ack(0);
      simple_obj_ref_2445_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to0_in0_pipe_read_req(0),
          oack => to0_in0_pipe_read_ack(0),
          odata => to0_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2590_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2592_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2592_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2590_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2590_inst_req_0;
      simple_obj_ref_2590_inst_ack_0 <= ack(0);
      data_in <= type_cast_2592_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2594_inst_ack_0 then -- 
          assert false report " WritePipe tofpga0_out0 from wire type_cast_2596_wire value="  &  convert_slv_to_hex_string(type_cast_2596_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2594_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2594_inst_req_0;
      simple_obj_ref_2594_inst_ack_0 <= ack(0);
      data_in <= type_cast_2596_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga0_out0_pipe_write_req(0),
          oack => tofpga0_out0_pipe_write_ack(0),
          odata => tofpga0_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2570_call call_stmt_2577_call call_stmt_2465_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2570_call_req_0;
      reqL(1) <= call_stmt_2577_call_req_0;
      reqL(0) <= call_stmt_2465_call_req_0;
      call_stmt_2570_call_ack_0 <= ackL(2);
      call_stmt_2577_call_ack_0 <= ackL(1);
      call_stmt_2465_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2570_call_req_1;
      reqR(1) <= call_stmt_2577_call_req_1;
      reqR(0) <= call_stmt_2465_call_req_1;
      call_stmt_2570_call_ack_1 <= ackR(2);
      call_stmt_2577_call_ack_1 <= ackR(1);
      call_stmt_2465_call_ack_1 <= ackR(0);
      data_in <= tmp16_2528 & tmp21_2567 & type_cast_2463_wire_constant;
      tmp22_2570 <= data_out(47 downto 32);
      tmp23_2577 <= data_out(31 downto 16);
      tmp4_2465 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to1 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to1_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to1_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to1_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga1_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to1;
architecture Default of ahir_glue_to1 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to1_CP_12747_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_2674_load_1_req_0 : boolean;
  signal ptr_deref_2674_load_2_req_1 : boolean;
  signal ptr_deref_2739_addr_0_req_0 : boolean;
  signal ptr_deref_2732_store_1_req_0 : boolean;
  signal binary_2726_inst_req_0 : boolean;
  signal type_cast_2678_inst_ack_0 : boolean;
  signal ptr_deref_2739_store_0_req_1 : boolean;
  signal binary_2703_inst_ack_0 : boolean;
  signal type_cast_2687_inst_req_0 : boolean;
  signal ptr_deref_2674_load_1_req_1 : boolean;
  signal ptr_deref_2739_addr_0_ack_1 : boolean;
  signal call_stmt_2737_call_ack_0 : boolean;
  signal array_obj_ref_2670_root_address_inst_req_1 : boolean;
  signal call_stmt_2737_call_ack_1 : boolean;
  signal type_cast_2721_inst_req_0 : boolean;
  signal ptr_deref_2739_addr_1_ack_1 : boolean;
  signal ptr_deref_2732_addr_1_req_0 : boolean;
  signal ptr_deref_2674_base_resize_req_0 : boolean;
  signal ptr_deref_2732_gather_scatter_req_0 : boolean;
  signal ptr_deref_2732_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2670_base_resize_ack_0 : boolean;
  signal ptr_deref_2739_store_0_ack_0 : boolean;
  signal binary_2709_inst_ack_0 : boolean;
  signal ptr_deref_2674_addr_3_ack_0 : boolean;
  signal ptr_deref_2744_base_resize_ack_0 : boolean;
  signal ptr_deref_2674_root_address_inst_ack_0 : boolean;
  signal type_cast_2721_inst_ack_0 : boolean;
  signal array_obj_ref_2670_base_resize_req_0 : boolean;
  signal type_cast_2687_inst_ack_0 : boolean;
  signal array_obj_ref_2670_root_address_inst_ack_0 : boolean;
  signal call_stmt_2737_call_req_1 : boolean;
  signal ptr_deref_2744_addr_0_ack_1 : boolean;
  signal ptr_deref_2739_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2739_addr_0_req_1 : boolean;
  signal type_cast_2697_inst_ack_0 : boolean;
  signal binary_2717_inst_req_0 : boolean;
  signal ptr_deref_2674_addr_3_req_0 : boolean;
  signal binary_2717_inst_ack_1 : boolean;
  signal ptr_deref_2674_addr_0_ack_1 : boolean;
  signal ptr_deref_2674_root_address_inst_req_0 : boolean;
  signal ptr_deref_2674_addr_1_ack_0 : boolean;
  signal ptr_deref_2674_addr_2_ack_0 : boolean;
  signal binary_2709_inst_req_0 : boolean;
  signal ptr_deref_2732_store_1_ack_0 : boolean;
  signal ptr_deref_2674_addr_1_ack_1 : boolean;
  signal ptr_deref_2744_addr_1_ack_0 : boolean;
  signal ptr_deref_2744_addr_2_req_0 : boolean;
  signal ptr_deref_2744_addr_1_req_0 : boolean;
  signal ptr_deref_2674_load_2_ack_0 : boolean;
  signal ptr_deref_2732_addr_0_req_1 : boolean;
  signal ptr_deref_2674_base_resize_ack_0 : boolean;
  signal binary_2703_inst_req_0 : boolean;
  signal array_obj_ref_2670_root_address_inst_ack_1 : boolean;
  signal type_cast_2697_inst_req_0 : boolean;
  signal binary_2726_inst_ack_0 : boolean;
  signal ptr_deref_2674_load_3_req_1 : boolean;
  signal ptr_deref_2674_load_0_req_0 : boolean;
  signal binary_2703_inst_req_1 : boolean;
  signal call_stmt_2730_call_ack_1 : boolean;
  signal array_obj_ref_2670_root_address_inst_req_0 : boolean;
  signal binary_2683_inst_ack_0 : boolean;
  signal ptr_deref_2744_addr_3_req_1 : boolean;
  signal ptr_deref_2744_addr_1_req_1 : boolean;
  signal ptr_deref_2744_addr_2_ack_0 : boolean;
  signal ptr_deref_2744_addr_2_req_1 : boolean;
  signal ptr_deref_2744_root_address_inst_req_0 : boolean;
  signal ptr_deref_2739_root_address_inst_req_0 : boolean;
  signal ptr_deref_2739_store_0_req_0 : boolean;
  signal ptr_deref_2732_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2744_addr_1_ack_1 : boolean;
  signal ptr_deref_2732_store_0_ack_0 : boolean;
  signal ptr_deref_2674_load_0_ack_0 : boolean;
  signal type_cast_2678_inst_req_0 : boolean;
  signal ptr_deref_2739_addr_1_req_1 : boolean;
  signal ptr_deref_2674_load_1_ack_1 : boolean;
  signal ptr_deref_2732_store_0_req_0 : boolean;
  signal binary_2709_inst_ack_1 : boolean;
  signal ptr_deref_2739_addr_0_ack_0 : boolean;
  signal binary_2683_inst_req_0 : boolean;
  signal binary_2703_inst_ack_1 : boolean;
  signal ptr_deref_2732_root_address_inst_req_0 : boolean;
  signal ptr_deref_2739_store_1_ack_1 : boolean;
  signal ptr_deref_2674_addr_0_req_1 : boolean;
  signal ptr_deref_2744_addr_0_req_0 : boolean;
  signal ptr_deref_2744_addr_3_ack_0 : boolean;
  signal binary_2683_inst_ack_1 : boolean;
  signal ptr_deref_2674_addr_1_req_1 : boolean;
  signal ptr_deref_2732_base_resize_ack_0 : boolean;
  signal ptr_deref_2739_store_1_req_1 : boolean;
  signal ptr_deref_2744_base_resize_req_0 : boolean;
  signal ptr_deref_2744_addr_0_req_1 : boolean;
  signal ptr_deref_2732_addr_0_ack_1 : boolean;
  signal binary_2709_inst_req_1 : boolean;
  signal ptr_deref_2744_root_address_inst_ack_0 : boolean;
  signal binary_2693_inst_ack_1 : boolean;
  signal binary_2683_inst_req_1 : boolean;
  signal ptr_deref_2744_addr_0_ack_0 : boolean;
  signal ptr_deref_2674_addr_1_req_0 : boolean;
  signal ptr_deref_2674_load_0_ack_1 : boolean;
  signal ptr_deref_2674_load_1_ack_0 : boolean;
  signal ptr_deref_2744_addr_2_ack_1 : boolean;
  signal ptr_deref_2744_addr_3_ack_1 : boolean;
  signal ptr_deref_2674_addr_2_ack_1 : boolean;
  signal binary_2726_inst_req_1 : boolean;
  signal ptr_deref_2739_base_resize_req_0 : boolean;
  signal type_cast_2713_inst_req_0 : boolean;
  signal binary_2726_inst_ack_1 : boolean;
  signal type_cast_2663_inst_req_0 : boolean;
  signal ptr_deref_2674_load_2_ack_1 : boolean;
  signal ptr_deref_2732_addr_1_ack_0 : boolean;
  signal ptr_deref_2732_store_0_req_1 : boolean;
  signal ptr_deref_2739_base_resize_ack_0 : boolean;
  signal ptr_deref_2732_addr_1_req_1 : boolean;
  signal ptr_deref_2732_store_0_ack_1 : boolean;
  signal ptr_deref_2744_addr_3_req_0 : boolean;
  signal ptr_deref_2674_addr_0_ack_0 : boolean;
  signal ptr_deref_2674_addr_0_req_0 : boolean;
  signal binary_2693_inst_req_1 : boolean;
  signal type_cast_2663_inst_ack_0 : boolean;
  signal ptr_deref_2732_store_1_req_1 : boolean;
  signal ptr_deref_2732_addr_0_req_0 : boolean;
  signal ptr_deref_2732_store_1_ack_1 : boolean;
  signal binary_2693_inst_req_0 : boolean;
  signal binary_2717_inst_ack_0 : boolean;
  signal ptr_deref_2739_addr_1_req_0 : boolean;
  signal ptr_deref_2674_addr_2_req_1 : boolean;
  signal ptr_deref_2674_load_2_req_0 : boolean;
  signal ptr_deref_2732_addr_1_ack_1 : boolean;
  signal ptr_deref_2739_store_0_ack_1 : boolean;
  signal ptr_deref_2744_load_0_req_0 : boolean;
  signal ptr_deref_2732_addr_0_ack_0 : boolean;
  signal ptr_deref_2732_base_resize_req_0 : boolean;
  signal ptr_deref_2674_addr_2_req_0 : boolean;
  signal binary_2717_inst_req_1 : boolean;
  signal ptr_deref_2739_addr_1_ack_0 : boolean;
  signal array_obj_ref_2670_final_reg_ack_0 : boolean;
  signal array_obj_ref_2670_final_reg_req_0 : boolean;
  signal call_stmt_2730_call_req_1 : boolean;
  signal type_cast_2713_inst_ack_0 : boolean;
  signal ptr_deref_2674_load_3_req_0 : boolean;
  signal ptr_deref_2674_addr_3_req_1 : boolean;
  signal ptr_deref_2674_load_3_ack_1 : boolean;
  signal ptr_deref_2674_addr_3_ack_1 : boolean;
  signal ptr_deref_2674_load_3_ack_0 : boolean;
  signal ptr_deref_2739_gather_scatter_req_0 : boolean;
  signal ptr_deref_2674_gather_scatter_req_0 : boolean;
  signal ptr_deref_2739_gather_scatter_ack_0 : boolean;
  signal call_stmt_2737_call_req_0 : boolean;
  signal call_stmt_2730_call_ack_0 : boolean;
  signal call_stmt_2730_call_req_0 : boolean;
  signal ptr_deref_2739_store_1_req_0 : boolean;
  signal ptr_deref_2674_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2674_load_0_req_1 : boolean;
  signal ptr_deref_2739_store_1_ack_0 : boolean;
  signal binary_2693_inst_ack_0 : boolean;
  signal simple_obj_ref_2605_inst_req_0 : boolean;
  signal simple_obj_ref_2605_inst_ack_0 : boolean;
  signal type_cast_2606_inst_req_0 : boolean;
  signal type_cast_2606_inst_ack_0 : boolean;
  signal type_cast_2610_inst_req_0 : boolean;
  signal type_cast_2610_inst_ack_0 : boolean;
  signal binary_2616_inst_req_0 : boolean;
  signal binary_2616_inst_ack_0 : boolean;
  signal binary_2616_inst_req_1 : boolean;
  signal binary_2616_inst_ack_1 : boolean;
  signal type_cast_2620_inst_req_0 : boolean;
  signal type_cast_2620_inst_ack_0 : boolean;
  signal call_stmt_2625_call_req_0 : boolean;
  signal call_stmt_2625_call_ack_0 : boolean;
  signal call_stmt_2625_call_req_1 : boolean;
  signal call_stmt_2625_call_ack_1 : boolean;
  signal ptr_deref_2627_base_resize_req_0 : boolean;
  signal ptr_deref_2627_base_resize_ack_0 : boolean;
  signal ptr_deref_2627_root_address_inst_req_0 : boolean;
  signal ptr_deref_2627_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2627_addr_0_req_0 : boolean;
  signal ptr_deref_2627_addr_0_ack_0 : boolean;
  signal ptr_deref_2627_addr_0_req_1 : boolean;
  signal ptr_deref_2627_addr_0_ack_1 : boolean;
  signal ptr_deref_2627_addr_1_req_0 : boolean;
  signal ptr_deref_2627_addr_1_ack_0 : boolean;
  signal ptr_deref_2627_addr_1_req_1 : boolean;
  signal ptr_deref_2627_addr_1_ack_1 : boolean;
  signal ptr_deref_2627_gather_scatter_req_0 : boolean;
  signal ptr_deref_2627_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2627_store_0_req_0 : boolean;
  signal ptr_deref_2627_store_0_ack_0 : boolean;
  signal ptr_deref_2627_store_1_req_0 : boolean;
  signal ptr_deref_2627_store_1_ack_0 : boolean;
  signal ptr_deref_2627_store_0_req_1 : boolean;
  signal ptr_deref_2627_store_0_ack_1 : boolean;
  signal ptr_deref_2627_store_1_req_1 : boolean;
  signal ptr_deref_2627_store_1_ack_1 : boolean;
  signal binary_2634_inst_req_0 : boolean;
  signal binary_2634_inst_ack_0 : boolean;
  signal binary_2634_inst_req_1 : boolean;
  signal binary_2634_inst_ack_1 : boolean;
  signal type_cast_2638_inst_req_0 : boolean;
  signal type_cast_2638_inst_ack_0 : boolean;
  signal binary_2644_inst_req_0 : boolean;
  signal binary_2644_inst_ack_0 : boolean;
  signal binary_2644_inst_req_1 : boolean;
  signal binary_2644_inst_ack_1 : boolean;
  signal ptr_deref_2744_load_0_ack_0 : boolean;
  signal type_cast_2648_inst_req_0 : boolean;
  signal type_cast_2648_inst_ack_0 : boolean;
  signal array_obj_ref_2655_base_resize_req_0 : boolean;
  signal array_obj_ref_2655_base_resize_ack_0 : boolean;
  signal array_obj_ref_2655_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2655_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2655_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2655_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2655_final_reg_req_0 : boolean;
  signal array_obj_ref_2655_final_reg_ack_0 : boolean;
  signal ptr_deref_2659_base_resize_req_0 : boolean;
  signal ptr_deref_2659_base_resize_ack_0 : boolean;
  signal ptr_deref_2659_root_address_inst_req_0 : boolean;
  signal ptr_deref_2659_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2659_addr_0_req_0 : boolean;
  signal ptr_deref_2659_addr_0_ack_0 : boolean;
  signal ptr_deref_2659_addr_0_req_1 : boolean;
  signal ptr_deref_2659_addr_0_ack_1 : boolean;
  signal ptr_deref_2659_addr_1_req_0 : boolean;
  signal ptr_deref_2659_addr_1_ack_0 : boolean;
  signal ptr_deref_2659_addr_1_req_1 : boolean;
  signal ptr_deref_2659_addr_1_ack_1 : boolean;
  signal ptr_deref_2659_addr_2_req_0 : boolean;
  signal ptr_deref_2659_addr_2_ack_0 : boolean;
  signal ptr_deref_2659_addr_2_req_1 : boolean;
  signal ptr_deref_2659_addr_2_ack_1 : boolean;
  signal ptr_deref_2659_addr_3_req_0 : boolean;
  signal ptr_deref_2659_addr_3_ack_0 : boolean;
  signal ptr_deref_2659_addr_3_req_1 : boolean;
  signal ptr_deref_2659_addr_3_ack_1 : boolean;
  signal ptr_deref_2659_load_0_req_0 : boolean;
  signal ptr_deref_2659_load_0_ack_0 : boolean;
  signal ptr_deref_2659_load_1_req_0 : boolean;
  signal ptr_deref_2659_load_1_ack_0 : boolean;
  signal ptr_deref_2659_load_2_req_0 : boolean;
  signal ptr_deref_2659_load_2_ack_0 : boolean;
  signal ptr_deref_2659_load_3_req_0 : boolean;
  signal ptr_deref_2659_load_3_ack_0 : boolean;
  signal ptr_deref_2659_load_0_req_1 : boolean;
  signal ptr_deref_2659_load_0_ack_1 : boolean;
  signal ptr_deref_2659_load_1_req_1 : boolean;
  signal ptr_deref_2659_load_1_ack_1 : boolean;
  signal ptr_deref_2659_load_2_req_1 : boolean;
  signal ptr_deref_2659_load_2_ack_1 : boolean;
  signal ptr_deref_2659_load_3_req_1 : boolean;
  signal ptr_deref_2659_load_3_ack_1 : boolean;
  signal ptr_deref_2659_gather_scatter_req_0 : boolean;
  signal ptr_deref_2659_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2744_load_1_req_0 : boolean;
  signal ptr_deref_2744_load_1_ack_0 : boolean;
  signal ptr_deref_2744_load_2_req_0 : boolean;
  signal ptr_deref_2744_load_2_ack_0 : boolean;
  signal ptr_deref_2744_load_3_req_0 : boolean;
  signal ptr_deref_2744_load_3_ack_0 : boolean;
  signal ptr_deref_2744_load_0_req_1 : boolean;
  signal ptr_deref_2744_load_0_ack_1 : boolean;
  signal ptr_deref_2744_load_1_req_1 : boolean;
  signal ptr_deref_2744_load_1_ack_1 : boolean;
  signal ptr_deref_2744_load_2_req_1 : boolean;
  signal ptr_deref_2744_load_2_ack_1 : boolean;
  signal ptr_deref_2744_load_3_req_1 : boolean;
  signal ptr_deref_2744_load_3_ack_1 : boolean;
  signal ptr_deref_2744_gather_scatter_req_0 : boolean;
  signal ptr_deref_2744_gather_scatter_ack_0 : boolean;
  signal type_cast_2748_inst_req_0 : boolean;
  signal type_cast_2748_inst_ack_0 : boolean;
  signal simple_obj_ref_2750_inst_req_0 : boolean;
  signal simple_obj_ref_2750_inst_ack_0 : boolean;
  signal type_cast_2756_inst_req_0 : boolean;
  signal type_cast_2756_inst_ack_0 : boolean;
  signal simple_obj_ref_2754_inst_req_0 : boolean;
  signal simple_obj_ref_2754_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to1_CP_12747: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_12838_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2625_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_13363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2730_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_13661_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2750_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2606_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_12788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2605_inst_req_0); -- 
    ack_12789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2605_inst_ack_0, ack => cp_elements(8)); -- 
    ack_12794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2606_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2610_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_12807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2610_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2616_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_12817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2616_inst_ack_0, ack => cp_elements(18)); -- 
    cr_12818_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2616_inst_req_1); -- 
    ca_12819_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2616_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2620_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_12829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2620_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_12839_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2625_call_ack_0, ack => cp_elements(24)); -- 
    ccr_12843_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2625_call_req_1); -- 
    cca_12844_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2625_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_12890_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2627_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_12863_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2627_base_resize_req_0); -- 
    base_resize_ack_12864_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_12868_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2627_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2627_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_12876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2627_addr_0_req_0); -- 
    ra_12877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_12878_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2627_addr_0_req_1); -- 
    ca_12879_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_12883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2627_addr_1_req_0); -- 
    ra_12884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_12885_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2627_addr_1_req_1); -- 
    ca_12886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2627_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_12898_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2627_store_0_req_0); -- 
    ra_12899_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_12903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2627_store_1_req_0); -- 
    ra_12904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_12914_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2627_store_0_req_1); -- 
    ca_12915_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_12919_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2627_store_1_req_1); -- 
    ca_12920_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2627_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2634_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_12930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2634_inst_ack_0, ack => cp_elements(55)); -- 
    cr_12931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2634_inst_req_1); -- 
    ca_12932_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2634_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2638_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_12942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2638_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_12951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2644_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_12952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2644_inst_ack_0, ack => cp_elements(63)); -- 
    cr_12953_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2644_inst_req_1); -- 
    ca_12954_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2644_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_12963_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2648_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_12964_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2648_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_12988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2655_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_12975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2655_base_resize_req_0); -- 
    base_resize_ack_12976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2655_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_12981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2655_root_address_inst_req_0); -- 
    plus_base_ra_12982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2655_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_12983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2655_root_address_inst_req_1); -- 
    plus_base_ca_12984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2655_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2655_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_13002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2659_base_resize_req_0); -- 
    base_resize_ack_13003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_13007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2659_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2659_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_13015_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2659_addr_0_req_0); -- 
    ra_13016_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_13017_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2659_addr_0_req_1); -- 
    ca_13018_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_13022_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2659_addr_1_req_0); -- 
    ra_13023_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_13024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2659_addr_1_req_1); -- 
    ca_13025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_13029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2659_addr_2_req_0); -- 
    ra_13030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_13031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2659_addr_2_req_1); -- 
    ca_13032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_13036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2659_addr_3_req_0); -- 
    ra_13037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_13038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2659_addr_3_req_1); -- 
    ca_13039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_13049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2659_load_0_req_0); -- 
    ra_13050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_13054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2659_load_1_req_0); -- 
    ra_13055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_13059_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2659_load_2_req_0); -- 
    ra_13060_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_13064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2659_load_3_req_0); -- 
    ra_13065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_13075_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2659_load_0_req_1); -- 
    ca_13076_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_13080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2659_load_1_req_1); -- 
    ca_13081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_13085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2659_load_2_req_1); -- 
    ca_13086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_13090_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2659_load_3_req_1); -- 
    ca_13091_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_13092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2659_gather_scatter_req_0); -- 
    merge_ack_13093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2659_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13102_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2663_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_13103_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2663_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_13127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2670_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_13114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2670_base_resize_req_0); -- 
    base_resize_ack_13115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2670_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_13120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2670_root_address_inst_req_0); -- 
    plus_base_ra_13121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2670_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_13122_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2670_root_address_inst_req_1); -- 
    plus_base_ca_13123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2670_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2670_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_13141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2674_base_resize_req_0); -- 
    base_resize_ack_13142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_13146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2674_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2674_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_13154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2674_addr_0_req_0); -- 
    ra_13155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_13156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2674_addr_0_req_1); -- 
    ca_13157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_13161_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2674_addr_1_req_0); -- 
    ra_13162_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_13163_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2674_addr_1_req_1); -- 
    ca_13164_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_13168_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2674_addr_2_req_0); -- 
    ra_13169_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_13170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2674_addr_2_req_1); -- 
    ca_13171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_13175_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2674_addr_3_req_0); -- 
    ra_13176_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_13177_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2674_addr_3_req_1); -- 
    ca_13178_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_13188_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2674_load_0_req_0); -- 
    ra_13189_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_13193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2674_load_1_req_0); -- 
    ra_13194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_13198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2674_load_2_req_0); -- 
    ra_13199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_13203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2674_load_3_req_0); -- 
    ra_13204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_13214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2674_load_0_req_1); -- 
    ca_13215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_13219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2674_load_1_req_1); -- 
    ca_13220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_13224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2674_load_2_req_1); -- 
    ca_13225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_13229_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2674_load_3_req_1); -- 
    ca_13230_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_13231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2674_gather_scatter_req_0); -- 
    merge_ack_13232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2674_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2678_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_13242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2678_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13252_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2683_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_13253_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2683_inst_ack_0, ack => cp_elements(162)); -- 
    cr_13254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2683_inst_req_1); -- 
    cp_elements(163) <= binary_2683_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13264_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2687_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_13265_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2687_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2693_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_13275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2693_inst_ack_0, ack => cp_elements(171)); -- 
    cr_13276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2693_inst_req_1); -- 
    ca_13277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2693_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2697_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_13287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2697_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2703_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_13297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2703_inst_ack_0, ack => cp_elements(178)); -- 
    cr_13298_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2703_inst_req_1); -- 
    ca_13299_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2703_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2709_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_13309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2709_inst_ack_0, ack => cp_elements(183)); -- 
    cr_13310_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2709_inst_req_1); -- 
    ca_13311_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2709_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2717_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13322_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2713_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_13323_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2713_inst_ack_0, ack => cp_elements(189)); -- 
    ra_13328_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2717_inst_ack_0, ack => cp_elements(190)); -- 
    cr_13329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2717_inst_req_1); -- 
    ca_13330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2717_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2721_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_13340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2721_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2726_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_13351_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2726_inst_ack_0, ack => cp_elements(197)); -- 
    cr_13352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2726_inst_req_1); -- 
    ca_13353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2726_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_13364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2730_call_ack_0, ack => cp_elements(200)); -- 
    ccr_13368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2730_call_req_1); -- 
    cca_13369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2730_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_13415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2732_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_13388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2732_base_resize_req_0); -- 
    base_resize_ack_13389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_13393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2732_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2732_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_13401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2732_addr_0_req_0); -- 
    ra_13402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_13403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2732_addr_0_req_1); -- 
    ca_13404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_13408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2732_addr_1_req_0); -- 
    ra_13409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_13410_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2732_addr_1_req_1); -- 
    ca_13411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2732_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_13423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2732_store_0_req_0); -- 
    ra_13424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_13428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2732_store_1_req_0); -- 
    ra_13429_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_13439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2732_store_0_req_1); -- 
    ca_13440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_13444_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2732_store_1_req_1); -- 
    ca_13445_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2732_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_13455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2737_call_req_0); -- 
    cra_13456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2737_call_ack_0, ack => cp_elements(227)); -- 
    ccr_13460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2737_call_req_1); -- 
    cca_13461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2737_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_13507_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2739_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_13480_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2739_base_resize_req_0); -- 
    base_resize_ack_13481_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_13485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2739_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2739_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_13493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2739_addr_0_req_0); -- 
    ra_13494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_13495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2739_addr_0_req_1); -- 
    ca_13496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_13500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2739_addr_1_req_0); -- 
    ra_13501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_13502_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2739_addr_1_req_1); -- 
    ca_13503_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2739_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_13515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2739_store_0_req_0); -- 
    ra_13516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_13520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2739_store_1_req_0); -- 
    ra_13521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_13531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2739_store_0_req_1); -- 
    ca_13532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_13536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2739_store_1_req_1); -- 
    ca_13537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2739_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_13550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2744_base_resize_req_0); -- 
    base_resize_ack_13551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_13555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2744_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2744_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_13563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2744_addr_0_req_0); -- 
    ra_13564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_13565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2744_addr_0_req_1); -- 
    ca_13566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_13570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2744_addr_1_req_0); -- 
    ra_13571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_13572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2744_addr_1_req_1); -- 
    ca_13573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_13577_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2744_addr_2_req_0); -- 
    ra_13578_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_13579_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2744_addr_2_req_1); -- 
    ca_13580_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_13584_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2744_addr_3_req_0); -- 
    ra_13585_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_13586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2744_addr_3_req_1); -- 
    ca_13587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_13597_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2744_load_0_req_0); -- 
    ra_13598_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_13602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2744_load_1_req_0); -- 
    ra_13603_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_13607_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2744_load_2_req_0); -- 
    ra_13608_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_13612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2744_load_3_req_0); -- 
    ra_13613_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_13623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2744_load_0_req_1); -- 
    ca_13624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_13628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2744_load_1_req_1); -- 
    ca_13629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_13633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2744_load_2_req_1); -- 
    ca_13634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_13638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2744_load_3_req_1); -- 
    ca_13639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_13640_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2744_gather_scatter_req_0); -- 
    merge_ack_13641_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2744_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2748_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_13651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2748_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_13662_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2750_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2756_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_13675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2756_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_13680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2754_inst_req_0); -- 
    pipe_wack_13681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2754_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2655_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2655_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2655_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2670_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2670_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2670_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2718 : std_logic_vector(0 downto 0);
    signal ptr_deref_2627_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2627_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2627_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2627_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2659_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2659_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2659_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2659_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2659_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2674_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2674_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2674_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2674_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2674_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2732_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2732_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2732_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2739_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2739_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2739_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2744_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2744_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2744_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2744_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2744_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2605_wire : std_logic_vector(31 downto 0);
    signal tmp10_2660 : std_logic_vector(31 downto 0);
    signal tmp11_2664 : std_logic_vector(31 downto 0);
    signal tmp12_2671 : std_logic_vector(31 downto 0);
    signal tmp13_2675 : std_logic_vector(31 downto 0);
    signal tmp14_2679 : std_logic_vector(31 downto 0);
    signal tmp15_2684 : std_logic_vector(31 downto 0);
    signal tmp16_2688 : std_logic_vector(15 downto 0);
    signal tmp17_2694 : std_logic_vector(31 downto 0);
    signal tmp18_2704 : std_logic_vector(15 downto 0);
    signal tmp19_2710 : std_logic_vector(31 downto 0);
    signal tmp1_2611 : std_logic_vector(31 downto 0);
    signal tmp20_2722 : std_logic_vector(15 downto 0);
    signal tmp21_2727 : std_logic_vector(15 downto 0);
    signal tmp22_2730 : std_logic_vector(15 downto 0);
    signal tmp23_2737 : std_logic_vector(15 downto 0);
    signal tmp24_2745 : std_logic_vector(31 downto 0);
    signal tmp25_2749 : std_logic_vector(31 downto 0);
    signal tmp2_2617 : std_logic_vector(31 downto 0);
    signal tmp3_2621 : std_logic_vector(31 downto 0);
    signal tmp4_2625 : std_logic_vector(15 downto 0);
    signal tmp5_2635 : std_logic_vector(31 downto 0);
    signal tmp6_2639 : std_logic_vector(31 downto 0);
    signal tmp7_2645 : std_logic_vector(31 downto 0);
    signal tmp8_2649 : std_logic_vector(31 downto 0);
    signal tmp9_2656 : std_logic_vector(31 downto 0);
    signal tmp_2607 : std_logic_vector(31 downto 0);
    signal type_cast_2615_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2623_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2633_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2643_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2692_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2702_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2708_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2713_wire : std_logic_vector(31 downto 0);
    signal type_cast_2716_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2752_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2756_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2698 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2655_final_offset <= "0000000000010000";
    array_obj_ref_2670_final_offset <= "0000000000001100";
    ptr_deref_2627_word_offset_0 <= "0000000000000000";
    ptr_deref_2627_word_offset_1 <= "0000000000000001";
    ptr_deref_2659_word_offset_0 <= "0000000000000000";
    ptr_deref_2659_word_offset_1 <= "0000000000000001";
    ptr_deref_2659_word_offset_2 <= "0000000000000010";
    ptr_deref_2659_word_offset_3 <= "0000000000000011";
    ptr_deref_2674_word_offset_0 <= "0000000000000000";
    ptr_deref_2674_word_offset_1 <= "0000000000000001";
    ptr_deref_2674_word_offset_2 <= "0000000000000010";
    ptr_deref_2674_word_offset_3 <= "0000000000000011";
    ptr_deref_2732_word_offset_0 <= "0000000000000000";
    ptr_deref_2732_word_offset_1 <= "0000000000000001";
    ptr_deref_2739_word_offset_0 <= "0000000000000000";
    ptr_deref_2739_word_offset_1 <= "0000000000000001";
    ptr_deref_2744_word_offset_0 <= "0000000000000000";
    ptr_deref_2744_word_offset_1 <= "0000000000000001";
    ptr_deref_2744_word_offset_2 <= "0000000000000010";
    ptr_deref_2744_word_offset_3 <= "0000000000000011";
    type_cast_2615_wire_constant <= "11111111111111111111100000000000";
    type_cast_2623_wire_constant <= "0000000000000010";
    type_cast_2633_wire_constant <= "00000000000000000000000000000110";
    type_cast_2643_wire_constant <= "00000000000000000000000000000010";
    type_cast_2692_wire_constant <= "00000000000000000000000000000011";
    type_cast_2702_wire_constant <= "0001111111111111";
    type_cast_2708_wire_constant <= "00000000000000000000000000000111";
    type_cast_2716_wire_constant <= "00000000000000000000000000000000";
    type_cast_2752_wire_constant <= "00000000000000000000000000000010";
    array_obj_ref_2655_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2611, dout => array_obj_ref_2655_resized_base_address, req => array_obj_ref_2655_base_resize_req_0, ack => array_obj_ref_2655_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2655_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2655_root_address, dout => tmp9_2656, req => array_obj_ref_2655_final_reg_req_0, ack => array_obj_ref_2655_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2670_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2611, dout => array_obj_ref_2670_resized_base_address, req => array_obj_ref_2670_base_resize_req_0, ack => array_obj_ref_2670_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2670_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2670_root_address, dout => tmp12_2671, req => array_obj_ref_2670_final_reg_req_0, ack => array_obj_ref_2670_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2627_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2621, dout => ptr_deref_2627_resized_base_address, req => ptr_deref_2627_base_resize_req_0, ack => ptr_deref_2627_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2659_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2656, dout => ptr_deref_2659_resized_base_address, req => ptr_deref_2659_base_resize_req_0, ack => ptr_deref_2659_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2674_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2671, dout => ptr_deref_2674_resized_base_address, req => ptr_deref_2674_base_resize_req_0, ack => ptr_deref_2674_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2732_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2639, dout => ptr_deref_2732_resized_base_address, req => ptr_deref_2732_base_resize_req_0, ack => ptr_deref_2732_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2739_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2649, dout => ptr_deref_2739_resized_base_address, req => ptr_deref_2739_base_resize_req_0, ack => ptr_deref_2739_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2744_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2671, dout => ptr_deref_2744_resized_base_address, req => ptr_deref_2744_base_resize_req_0, ack => ptr_deref_2744_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2606_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2605_wire, dout => tmp_2607, req => type_cast_2606_inst_req_0, ack => type_cast_2606_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2610_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2607, dout => tmp1_2611, req => type_cast_2610_inst_req_0, ack => type_cast_2610_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2620_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2617, dout => tmp3_2621, req => type_cast_2620_inst_req_0, ack => type_cast_2620_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2638_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2635, dout => tmp6_2639, req => type_cast_2638_inst_req_0, ack => type_cast_2638_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2648_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2645, dout => tmp8_2649, req => type_cast_2648_inst_req_0, ack => type_cast_2648_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2663_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2660, dout => tmp11_2664, req => type_cast_2663_inst_req_0, ack => type_cast_2663_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2678_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2675, dout => tmp14_2679, req => type_cast_2678_inst_req_0, ack => type_cast_2678_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2687_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2684, dout => tmp16_2688, req => type_cast_2687_inst_req_0, ack => type_cast_2687_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2697_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2694, dout => xx_xtrx_xi_2698, req => type_cast_2697_inst_req_0, ack => type_cast_2697_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2713_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2710, dout => type_cast_2713_wire, req => type_cast_2713_inst_req_0, ack => type_cast_2713_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2721_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2718, dout => tmp20_2722, req => type_cast_2721_inst_req_0, ack => type_cast_2721_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2748_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2745, dout => tmp25_2749, req => type_cast_2748_inst_req_0, ack => type_cast_2748_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2756_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2749, dout => type_cast_2756_wire, req => type_cast_2756_inst_req_0, ack => type_cast_2756_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2627_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2627_gather_scatter_ack_0 <= ptr_deref_2627_gather_scatter_req_0;
      aggregated_sig <= tmp4_2625;
      ptr_deref_2627_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2627_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2627_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2627_root_address_inst_ack_0 <= ptr_deref_2627_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2627_resized_base_address;
      ptr_deref_2627_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2659_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2659_gather_scatter_ack_0 <= ptr_deref_2659_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2659_data_3 & ptr_deref_2659_data_2 & ptr_deref_2659_data_1 & ptr_deref_2659_data_0;
      tmp10_2660 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2659_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2659_root_address_inst_ack_0 <= ptr_deref_2659_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2659_resized_base_address;
      ptr_deref_2659_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2674_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2674_gather_scatter_ack_0 <= ptr_deref_2674_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2674_data_3 & ptr_deref_2674_data_2 & ptr_deref_2674_data_1 & ptr_deref_2674_data_0;
      tmp13_2675 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2674_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2674_root_address_inst_ack_0 <= ptr_deref_2674_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2674_resized_base_address;
      ptr_deref_2674_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2732_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2732_gather_scatter_ack_0 <= ptr_deref_2732_gather_scatter_req_0;
      aggregated_sig <= tmp22_2730;
      ptr_deref_2732_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2732_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2732_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2732_root_address_inst_ack_0 <= ptr_deref_2732_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2732_resized_base_address;
      ptr_deref_2732_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2739_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2739_gather_scatter_ack_0 <= ptr_deref_2739_gather_scatter_req_0;
      aggregated_sig <= tmp23_2737;
      ptr_deref_2739_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2739_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2739_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2739_root_address_inst_ack_0 <= ptr_deref_2739_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2739_resized_base_address;
      ptr_deref_2739_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2744_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2744_gather_scatter_ack_0 <= ptr_deref_2744_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2744_data_3 & ptr_deref_2744_data_2 & ptr_deref_2744_data_1 & ptr_deref_2744_data_0;
      tmp24_2745 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2744_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2744_root_address_inst_ack_0 <= ptr_deref_2744_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2744_resized_base_address;
      ptr_deref_2744_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2655_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2655_resized_base_address;
      array_obj_ref_2655_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2655_root_address_inst_req_0,
          ackL => array_obj_ref_2655_root_address_inst_ack_0,
          reqR => array_obj_ref_2655_root_address_inst_req_1,
          ackR => array_obj_ref_2655_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2670_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2670_resized_base_address;
      array_obj_ref_2670_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2670_root_address_inst_req_0,
          ackL => array_obj_ref_2670_root_address_inst_ack_0,
          reqR => array_obj_ref_2670_root_address_inst_req_1,
          ackR => array_obj_ref_2670_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2616_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2607;
      tmp2_2617 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2616_inst_req_0,
          ackL => binary_2616_inst_ack_0,
          reqR => binary_2616_inst_req_1,
          ackR => binary_2616_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2634_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2617;
      tmp5_2635 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2634_inst_req_0,
          ackL => binary_2634_inst_ack_0,
          reqR => binary_2634_inst_req_1,
          ackR => binary_2634_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2644_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2617;
      tmp7_2645 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2644_inst_req_0,
          ackL => binary_2644_inst_ack_0,
          reqR => binary_2644_inst_req_1,
          ackR => binary_2644_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2683_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2664 & tmp14_2679;
      tmp15_2684 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2683_inst_req_0,
          ackL => binary_2683_inst_ack_0,
          reqR => binary_2683_inst_req_1,
          ackR => binary_2683_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2693_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2684;
      tmp17_2694 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2693_inst_req_0,
          ackL => binary_2693_inst_ack_0,
          reqR => binary_2693_inst_req_1,
          ackR => binary_2693_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2703_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2698;
      tmp18_2704 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2703_inst_req_0,
          ackL => binary_2703_inst_ack_0,
          reqR => binary_2703_inst_req_1,
          ackR => binary_2703_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2709_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2684;
      tmp19_2710 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2709_inst_req_0,
          ackL => binary_2709_inst_ack_0,
          reqR => binary_2709_inst_req_1,
          ackR => binary_2709_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2717_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2713_wire;
      notx_xx_xi_2718 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2717_inst_req_0,
          ackL => binary_2717_inst_ack_0,
          reqR => binary_2717_inst_req_1,
          ackR => binary_2717_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2726_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2704 & tmp20_2722;
      tmp21_2727 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2726_inst_req_0,
          ackL => binary_2726_inst_ack_0,
          reqR => binary_2726_inst_req_1,
          ackR => binary_2726_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2627_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2627_root_address;
      ptr_deref_2627_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2627_addr_0_req_0,
          ackL => ptr_deref_2627_addr_0_ack_0,
          reqR => ptr_deref_2627_addr_0_req_1,
          ackR => ptr_deref_2627_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2627_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2627_root_address;
      ptr_deref_2627_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2627_addr_1_req_0,
          ackL => ptr_deref_2627_addr_1_ack_0,
          reqR => ptr_deref_2627_addr_1_req_1,
          ackR => ptr_deref_2627_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2659_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2659_root_address;
      ptr_deref_2659_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2659_addr_0_req_0,
          ackL => ptr_deref_2659_addr_0_ack_0,
          reqR => ptr_deref_2659_addr_0_req_1,
          ackR => ptr_deref_2659_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2659_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2659_root_address;
      ptr_deref_2659_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2659_addr_1_req_0,
          ackL => ptr_deref_2659_addr_1_ack_0,
          reqR => ptr_deref_2659_addr_1_req_1,
          ackR => ptr_deref_2659_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2659_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2659_root_address;
      ptr_deref_2659_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2659_addr_2_req_0,
          ackL => ptr_deref_2659_addr_2_ack_0,
          reqR => ptr_deref_2659_addr_2_req_1,
          ackR => ptr_deref_2659_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2659_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2659_root_address;
      ptr_deref_2659_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2659_addr_3_req_0,
          ackL => ptr_deref_2659_addr_3_ack_0,
          reqR => ptr_deref_2659_addr_3_req_1,
          ackR => ptr_deref_2659_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2674_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2674_root_address;
      ptr_deref_2674_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2674_addr_0_req_0,
          ackL => ptr_deref_2674_addr_0_ack_0,
          reqR => ptr_deref_2674_addr_0_req_1,
          ackR => ptr_deref_2674_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2674_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2674_root_address;
      ptr_deref_2674_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2674_addr_1_req_0,
          ackL => ptr_deref_2674_addr_1_ack_0,
          reqR => ptr_deref_2674_addr_1_req_1,
          ackR => ptr_deref_2674_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2674_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2674_root_address;
      ptr_deref_2674_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2674_addr_2_req_0,
          ackL => ptr_deref_2674_addr_2_ack_0,
          reqR => ptr_deref_2674_addr_2_req_1,
          ackR => ptr_deref_2674_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2674_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2674_root_address;
      ptr_deref_2674_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2674_addr_3_req_0,
          ackL => ptr_deref_2674_addr_3_ack_0,
          reqR => ptr_deref_2674_addr_3_req_1,
          ackR => ptr_deref_2674_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2732_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2732_root_address;
      ptr_deref_2732_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2732_addr_0_req_0,
          ackL => ptr_deref_2732_addr_0_ack_0,
          reqR => ptr_deref_2732_addr_0_req_1,
          ackR => ptr_deref_2732_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2732_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2732_root_address;
      ptr_deref_2732_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2732_addr_1_req_0,
          ackL => ptr_deref_2732_addr_1_ack_0,
          reqR => ptr_deref_2732_addr_1_req_1,
          ackR => ptr_deref_2732_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2739_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2739_root_address;
      ptr_deref_2739_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2739_addr_0_req_0,
          ackL => ptr_deref_2739_addr_0_ack_0,
          reqR => ptr_deref_2739_addr_0_req_1,
          ackR => ptr_deref_2739_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2739_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2739_root_address;
      ptr_deref_2739_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2739_addr_1_req_0,
          ackL => ptr_deref_2739_addr_1_ack_0,
          reqR => ptr_deref_2739_addr_1_req_1,
          ackR => ptr_deref_2739_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2744_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2744_root_address;
      ptr_deref_2744_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2744_addr_0_req_0,
          ackL => ptr_deref_2744_addr_0_ack_0,
          reqR => ptr_deref_2744_addr_0_req_1,
          ackR => ptr_deref_2744_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2744_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2744_root_address;
      ptr_deref_2744_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2744_addr_1_req_0,
          ackL => ptr_deref_2744_addr_1_ack_0,
          reqR => ptr_deref_2744_addr_1_req_1,
          ackR => ptr_deref_2744_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2744_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2744_root_address;
      ptr_deref_2744_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2744_addr_2_req_0,
          ackL => ptr_deref_2744_addr_2_ack_0,
          reqR => ptr_deref_2744_addr_2_req_1,
          ackR => ptr_deref_2744_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2744_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2744_root_address;
      ptr_deref_2744_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2744_addr_3_req_0,
          ackL => ptr_deref_2744_addr_3_ack_0,
          reqR => ptr_deref_2744_addr_3_req_1,
          ackR => ptr_deref_2744_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2744_load_1 ptr_deref_2744_load_3 ptr_deref_2744_load_0 ptr_deref_2659_load_3 ptr_deref_2659_load_2 ptr_deref_2659_load_1 ptr_deref_2659_load_0 ptr_deref_2744_load_2 ptr_deref_2674_load_0 ptr_deref_2674_load_1 ptr_deref_2674_load_2 ptr_deref_2674_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2744_load_1_req_0,
        ptr_deref_2744_load_1_ack_0,
        ptr_deref_2744_load_1_req_1,
        ptr_deref_2744_load_1_ack_1,
        "ptr_deref_2744_load_1",
        "memory_space_5" ,
        ptr_deref_2744_data_1,
        ptr_deref_2744_word_address_1,
        "ptr_deref_2744_data_1",
        "ptr_deref_2744_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2744_load_3_req_0,
        ptr_deref_2744_load_3_ack_0,
        ptr_deref_2744_load_3_req_1,
        ptr_deref_2744_load_3_ack_1,
        "ptr_deref_2744_load_3",
        "memory_space_5" ,
        ptr_deref_2744_data_3,
        ptr_deref_2744_word_address_3,
        "ptr_deref_2744_data_3",
        "ptr_deref_2744_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2744_load_0_req_0,
        ptr_deref_2744_load_0_ack_0,
        ptr_deref_2744_load_0_req_1,
        ptr_deref_2744_load_0_ack_1,
        "ptr_deref_2744_load_0",
        "memory_space_5" ,
        ptr_deref_2744_data_0,
        ptr_deref_2744_word_address_0,
        "ptr_deref_2744_data_0",
        "ptr_deref_2744_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2659_load_3_req_0,
        ptr_deref_2659_load_3_ack_0,
        ptr_deref_2659_load_3_req_1,
        ptr_deref_2659_load_3_ack_1,
        "ptr_deref_2659_load_3",
        "memory_space_5" ,
        ptr_deref_2659_data_3,
        ptr_deref_2659_word_address_3,
        "ptr_deref_2659_data_3",
        "ptr_deref_2659_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2659_load_2_req_0,
        ptr_deref_2659_load_2_ack_0,
        ptr_deref_2659_load_2_req_1,
        ptr_deref_2659_load_2_ack_1,
        "ptr_deref_2659_load_2",
        "memory_space_5" ,
        ptr_deref_2659_data_2,
        ptr_deref_2659_word_address_2,
        "ptr_deref_2659_data_2",
        "ptr_deref_2659_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2659_load_1_req_0,
        ptr_deref_2659_load_1_ack_0,
        ptr_deref_2659_load_1_req_1,
        ptr_deref_2659_load_1_ack_1,
        "ptr_deref_2659_load_1",
        "memory_space_5" ,
        ptr_deref_2659_data_1,
        ptr_deref_2659_word_address_1,
        "ptr_deref_2659_data_1",
        "ptr_deref_2659_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2659_load_0_req_0,
        ptr_deref_2659_load_0_ack_0,
        ptr_deref_2659_load_0_req_1,
        ptr_deref_2659_load_0_ack_1,
        "ptr_deref_2659_load_0",
        "memory_space_5" ,
        ptr_deref_2659_data_0,
        ptr_deref_2659_word_address_0,
        "ptr_deref_2659_data_0",
        "ptr_deref_2659_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2744_load_2_req_0,
        ptr_deref_2744_load_2_ack_0,
        ptr_deref_2744_load_2_req_1,
        ptr_deref_2744_load_2_ack_1,
        "ptr_deref_2744_load_2",
        "memory_space_5" ,
        ptr_deref_2744_data_2,
        ptr_deref_2744_word_address_2,
        "ptr_deref_2744_data_2",
        "ptr_deref_2744_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2674_load_0_req_0,
        ptr_deref_2674_load_0_ack_0,
        ptr_deref_2674_load_0_req_1,
        ptr_deref_2674_load_0_ack_1,
        "ptr_deref_2674_load_0",
        "memory_space_5" ,
        ptr_deref_2674_data_0,
        ptr_deref_2674_word_address_0,
        "ptr_deref_2674_data_0",
        "ptr_deref_2674_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2674_load_1_req_0,
        ptr_deref_2674_load_1_ack_0,
        ptr_deref_2674_load_1_req_1,
        ptr_deref_2674_load_1_ack_1,
        "ptr_deref_2674_load_1",
        "memory_space_5" ,
        ptr_deref_2674_data_1,
        ptr_deref_2674_word_address_1,
        "ptr_deref_2674_data_1",
        "ptr_deref_2674_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2674_load_2_req_0,
        ptr_deref_2674_load_2_ack_0,
        ptr_deref_2674_load_2_req_1,
        ptr_deref_2674_load_2_ack_1,
        "ptr_deref_2674_load_2",
        "memory_space_5" ,
        ptr_deref_2674_data_2,
        ptr_deref_2674_word_address_2,
        "ptr_deref_2674_data_2",
        "ptr_deref_2674_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2674_load_3_req_0,
        ptr_deref_2674_load_3_ack_0,
        ptr_deref_2674_load_3_req_1,
        ptr_deref_2674_load_3_ack_1,
        "ptr_deref_2674_load_3",
        "memory_space_5" ,
        ptr_deref_2674_data_3,
        ptr_deref_2674_word_address_3,
        "ptr_deref_2674_data_3",
        "ptr_deref_2674_word_address_3" -- 
      );
      reqL(11) <= ptr_deref_2744_load_1_req_0;
      reqL(10) <= ptr_deref_2744_load_3_req_0;
      reqL(9) <= ptr_deref_2744_load_0_req_0;
      reqL(8) <= ptr_deref_2659_load_3_req_0;
      reqL(7) <= ptr_deref_2659_load_2_req_0;
      reqL(6) <= ptr_deref_2659_load_1_req_0;
      reqL(5) <= ptr_deref_2659_load_0_req_0;
      reqL(4) <= ptr_deref_2744_load_2_req_0;
      reqL(3) <= ptr_deref_2674_load_0_req_0;
      reqL(2) <= ptr_deref_2674_load_1_req_0;
      reqL(1) <= ptr_deref_2674_load_2_req_0;
      reqL(0) <= ptr_deref_2674_load_3_req_0;
      ptr_deref_2744_load_1_ack_0 <= ackL(11);
      ptr_deref_2744_load_3_ack_0 <= ackL(10);
      ptr_deref_2744_load_0_ack_0 <= ackL(9);
      ptr_deref_2659_load_3_ack_0 <= ackL(8);
      ptr_deref_2659_load_2_ack_0 <= ackL(7);
      ptr_deref_2659_load_1_ack_0 <= ackL(6);
      ptr_deref_2659_load_0_ack_0 <= ackL(5);
      ptr_deref_2744_load_2_ack_0 <= ackL(4);
      ptr_deref_2674_load_0_ack_0 <= ackL(3);
      ptr_deref_2674_load_1_ack_0 <= ackL(2);
      ptr_deref_2674_load_2_ack_0 <= ackL(1);
      ptr_deref_2674_load_3_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2744_load_1_req_1;
      reqR(10) <= ptr_deref_2744_load_3_req_1;
      reqR(9) <= ptr_deref_2744_load_0_req_1;
      reqR(8) <= ptr_deref_2659_load_3_req_1;
      reqR(7) <= ptr_deref_2659_load_2_req_1;
      reqR(6) <= ptr_deref_2659_load_1_req_1;
      reqR(5) <= ptr_deref_2659_load_0_req_1;
      reqR(4) <= ptr_deref_2744_load_2_req_1;
      reqR(3) <= ptr_deref_2674_load_0_req_1;
      reqR(2) <= ptr_deref_2674_load_1_req_1;
      reqR(1) <= ptr_deref_2674_load_2_req_1;
      reqR(0) <= ptr_deref_2674_load_3_req_1;
      ptr_deref_2744_load_1_ack_1 <= ackR(11);
      ptr_deref_2744_load_3_ack_1 <= ackR(10);
      ptr_deref_2744_load_0_ack_1 <= ackR(9);
      ptr_deref_2659_load_3_ack_1 <= ackR(8);
      ptr_deref_2659_load_2_ack_1 <= ackR(7);
      ptr_deref_2659_load_1_ack_1 <= ackR(6);
      ptr_deref_2659_load_0_ack_1 <= ackR(5);
      ptr_deref_2744_load_2_ack_1 <= ackR(4);
      ptr_deref_2674_load_0_ack_1 <= ackR(3);
      ptr_deref_2674_load_1_ack_1 <= ackR(2);
      ptr_deref_2674_load_2_ack_1 <= ackR(1);
      ptr_deref_2674_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_2744_word_address_1 & ptr_deref_2744_word_address_3 & ptr_deref_2744_word_address_0 & ptr_deref_2659_word_address_3 & ptr_deref_2659_word_address_2 & ptr_deref_2659_word_address_1 & ptr_deref_2659_word_address_0 & ptr_deref_2744_word_address_2 & ptr_deref_2674_word_address_0 & ptr_deref_2674_word_address_1 & ptr_deref_2674_word_address_2 & ptr_deref_2674_word_address_3;
      ptr_deref_2744_data_1 <= data_out(95 downto 88);
      ptr_deref_2744_data_3 <= data_out(87 downto 80);
      ptr_deref_2744_data_0 <= data_out(79 downto 72);
      ptr_deref_2659_data_3 <= data_out(71 downto 64);
      ptr_deref_2659_data_2 <= data_out(63 downto 56);
      ptr_deref_2659_data_1 <= data_out(55 downto 48);
      ptr_deref_2659_data_0 <= data_out(47 downto 40);
      ptr_deref_2744_data_2 <= data_out(39 downto 32);
      ptr_deref_2674_data_0 <= data_out(31 downto 24);
      ptr_deref_2674_data_1 <= data_out(23 downto 16);
      ptr_deref_2674_data_2 <= data_out(15 downto 8);
      ptr_deref_2674_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2732_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2732_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2732_word_address_0) &  " data ptr_deref_2732_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2732_data_0) severity note; --
        end if;
        if ptr_deref_2739_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2739_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2739_word_address_1) &  " data ptr_deref_2739_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2739_data_1) severity note; --
        end if;
        if ptr_deref_2627_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2627_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2627_word_address_0) &  " data ptr_deref_2627_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2627_data_0) severity note; --
        end if;
        if ptr_deref_2739_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2739_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2739_word_address_0) &  " data ptr_deref_2739_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2739_data_0) severity note; --
        end if;
        if ptr_deref_2732_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2732_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2732_word_address_1) &  " data ptr_deref_2732_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2732_data_1) severity note; --
        end if;
        if ptr_deref_2627_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2627_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2627_word_address_1) &  " data ptr_deref_2627_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2627_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2732_store_0 ptr_deref_2739_store_1 ptr_deref_2627_store_0 ptr_deref_2739_store_0 ptr_deref_2732_store_1 ptr_deref_2627_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2732_store_0_req_0;
      reqL(4) <= ptr_deref_2739_store_1_req_0;
      reqL(3) <= ptr_deref_2627_store_0_req_0;
      reqL(2) <= ptr_deref_2739_store_0_req_0;
      reqL(1) <= ptr_deref_2732_store_1_req_0;
      reqL(0) <= ptr_deref_2627_store_1_req_0;
      ptr_deref_2732_store_0_ack_0 <= ackL(5);
      ptr_deref_2739_store_1_ack_0 <= ackL(4);
      ptr_deref_2627_store_0_ack_0 <= ackL(3);
      ptr_deref_2739_store_0_ack_0 <= ackL(2);
      ptr_deref_2732_store_1_ack_0 <= ackL(1);
      ptr_deref_2627_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2732_store_0_req_1;
      reqR(4) <= ptr_deref_2739_store_1_req_1;
      reqR(3) <= ptr_deref_2627_store_0_req_1;
      reqR(2) <= ptr_deref_2739_store_0_req_1;
      reqR(1) <= ptr_deref_2732_store_1_req_1;
      reqR(0) <= ptr_deref_2627_store_1_req_1;
      ptr_deref_2732_store_0_ack_1 <= ackR(5);
      ptr_deref_2739_store_1_ack_1 <= ackR(4);
      ptr_deref_2627_store_0_ack_1 <= ackR(3);
      ptr_deref_2739_store_0_ack_1 <= ackR(2);
      ptr_deref_2732_store_1_ack_1 <= ackR(1);
      ptr_deref_2627_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2732_word_address_0 & ptr_deref_2739_word_address_1 & ptr_deref_2627_word_address_0 & ptr_deref_2739_word_address_0 & ptr_deref_2732_word_address_1 & ptr_deref_2627_word_address_1;
      data_in <= ptr_deref_2732_data_0 & ptr_deref_2739_data_1 & ptr_deref_2627_data_0 & ptr_deref_2739_data_0 & ptr_deref_2732_data_1 & ptr_deref_2627_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2605_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2605_inst_ack_0 then -- 
            assert false report " ReadPipe to1_in0 to wire simple_obj_ref_2605_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2605_inst_req_0;
      simple_obj_ref_2605_inst_ack_0 <= ack(0);
      simple_obj_ref_2605_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to1_in0_pipe_read_req(0),
          oack => to1_in0_pipe_read_ack(0),
          odata => to1_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2750_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2752_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2752_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2750_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2750_inst_req_0;
      simple_obj_ref_2750_inst_ack_0 <= ack(0);
      data_in <= type_cast_2752_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2754_inst_ack_0 then -- 
          assert false report " WritePipe tofpga1_out0 from wire type_cast_2756_wire value="  &  convert_slv_to_hex_string(type_cast_2756_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2754_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2754_inst_req_0;
      simple_obj_ref_2754_inst_ack_0 <= ack(0);
      data_in <= type_cast_2756_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga1_out0_pipe_write_req(0),
          oack => tofpga1_out0_pipe_write_ack(0),
          odata => tofpga1_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2737_call call_stmt_2730_call call_stmt_2625_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2737_call_req_0;
      reqL(1) <= call_stmt_2730_call_req_0;
      reqL(0) <= call_stmt_2625_call_req_0;
      call_stmt_2737_call_ack_0 <= ackL(2);
      call_stmt_2730_call_ack_0 <= ackL(1);
      call_stmt_2625_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2737_call_req_1;
      reqR(1) <= call_stmt_2730_call_req_1;
      reqR(0) <= call_stmt_2625_call_req_1;
      call_stmt_2737_call_ack_1 <= ackR(2);
      call_stmt_2730_call_ack_1 <= ackR(1);
      call_stmt_2625_call_ack_1 <= ackR(0);
      data_in <= tmp21_2727 & tmp16_2688 & type_cast_2623_wire_constant;
      tmp23_2737 <= data_out(47 downto 32);
      tmp22_2730 <= data_out(31 downto 16);
      tmp4_2625 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to2_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to2_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to2_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga2_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to2;
architecture Default of ahir_glue_to2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to2_CP_13690_start: Boolean;
  -- links between control-path and data-path
  signal binary_2843_inst_ack_0 : boolean;
  signal array_obj_ref_2830_root_address_inst_req_1 : boolean;
  signal ptr_deref_2834_addr_2_req_0 : boolean;
  signal ptr_deref_2834_addr_3_req_1 : boolean;
  signal binary_2853_inst_ack_0 : boolean;
  signal ptr_deref_2899_base_resize_ack_0 : boolean;
  signal ptr_deref_2899_addr_0_req_0 : boolean;
  signal ptr_deref_2892_store_0_req_1 : boolean;
  signal array_obj_ref_2830_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2892_base_resize_ack_0 : boolean;
  signal ptr_deref_2834_load_3_req_0 : boolean;
  signal ptr_deref_2834_load_1_ack_1 : boolean;
  signal array_obj_ref_2830_final_reg_ack_0 : boolean;
  signal ptr_deref_2904_base_resize_req_0 : boolean;
  signal binary_2853_inst_req_0 : boolean;
  signal ptr_deref_2904_load_0_req_0 : boolean;
  signal ptr_deref_2899_addr_0_ack_0 : boolean;
  signal ptr_deref_2892_store_0_ack_1 : boolean;
  signal binary_2843_inst_ack_1 : boolean;
  signal array_obj_ref_2830_base_resize_req_0 : boolean;
  signal ptr_deref_2834_addr_3_ack_0 : boolean;
  signal ptr_deref_2834_addr_0_req_1 : boolean;
  signal binary_2853_inst_req_1 : boolean;
  signal ptr_deref_2834_load_2_ack_1 : boolean;
  signal ptr_deref_2834_addr_1_ack_1 : boolean;
  signal binary_2877_inst_req_1 : boolean;
  signal ptr_deref_2834_addr_3_req_0 : boolean;
  signal binary_2853_inst_ack_1 : boolean;
  signal ptr_deref_2834_load_0_ack_0 : boolean;
  signal ptr_deref_2904_addr_3_ack_1 : boolean;
  signal ptr_deref_2899_store_1_ack_1 : boolean;
  signal ptr_deref_2904_addr_0_ack_1 : boolean;
  signal ptr_deref_2904_load_1_req_0 : boolean;
  signal ptr_deref_2904_load_0_ack_1 : boolean;
  signal ptr_deref_2904_load_1_ack_1 : boolean;
  signal ptr_deref_2892_base_resize_req_0 : boolean;
  signal call_stmt_2890_call_req_0 : boolean;
  signal ptr_deref_2834_addr_1_req_0 : boolean;
  signal ptr_deref_2904_addr_0_req_1 : boolean;
  signal type_cast_2838_inst_req_0 : boolean;
  signal binary_2886_inst_req_1 : boolean;
  signal call_stmt_2897_call_req_0 : boolean;
  signal ptr_deref_2899_root_address_inst_req_0 : boolean;
  signal ptr_deref_2899_addr_0_req_1 : boolean;
  signal binary_2886_inst_ack_0 : boolean;
  signal ptr_deref_2834_addr_1_ack_0 : boolean;
  signal type_cast_2847_inst_req_0 : boolean;
  signal array_obj_ref_2830_base_resize_ack_0 : boolean;
  signal ptr_deref_2834_addr_1_req_1 : boolean;
  signal ptr_deref_2834_load_1_req_1 : boolean;
  signal ptr_deref_2834_addr_0_ack_1 : boolean;
  signal ptr_deref_2834_load_2_req_1 : boolean;
  signal ptr_deref_2904_addr_2_req_0 : boolean;
  signal ptr_deref_2892_addr_0_ack_1 : boolean;
  signal ptr_deref_2899_store_1_req_1 : boolean;
  signal ptr_deref_2834_load_2_req_0 : boolean;
  signal ptr_deref_2904_addr_0_ack_0 : boolean;
  signal ptr_deref_2834_addr_2_ack_0 : boolean;
  signal array_obj_ref_2830_final_reg_req_0 : boolean;
  signal type_cast_2823_inst_req_0 : boolean;
  signal ptr_deref_2904_addr_3_ack_0 : boolean;
  signal type_cast_2838_inst_ack_0 : boolean;
  signal binary_2877_inst_ack_0 : boolean;
  signal type_cast_2847_inst_ack_0 : boolean;
  signal ptr_deref_2904_addr_1_ack_1 : boolean;
  signal type_cast_2823_inst_ack_0 : boolean;
  signal ptr_deref_2899_store_0_req_1 : boolean;
  signal ptr_deref_2904_addr_2_req_1 : boolean;
  signal ptr_deref_2904_base_resize_ack_0 : boolean;
  signal array_obj_ref_2830_root_address_inst_req_0 : boolean;
  signal binary_2863_inst_req_0 : boolean;
  signal binary_2869_inst_req_1 : boolean;
  signal type_cast_2857_inst_ack_0 : boolean;
  signal ptr_deref_2892_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_2830_root_address_inst_ack_1 : boolean;
  signal simple_obj_ref_2910_inst_req_0 : boolean;
  signal ptr_deref_2899_gather_scatter_req_0 : boolean;
  signal ptr_deref_2899_store_1_req_0 : boolean;
  signal binary_2863_inst_ack_1 : boolean;
  signal ptr_deref_2904_load_2_req_0 : boolean;
  signal ptr_deref_2904_addr_0_req_0 : boolean;
  signal binary_2863_inst_req_1 : boolean;
  signal binary_2843_inst_req_1 : boolean;
  signal ptr_deref_2834_load_0_req_0 : boolean;
  signal ptr_deref_2904_addr_3_req_1 : boolean;
  signal ptr_deref_2899_store_0_ack_1 : boolean;
  signal ptr_deref_2834_addr_0_ack_0 : boolean;
  signal binary_2886_inst_ack_1 : boolean;
  signal binary_2843_inst_req_0 : boolean;
  signal binary_2869_inst_ack_1 : boolean;
  signal type_cast_2857_inst_req_0 : boolean;
  signal ptr_deref_2904_load_2_ack_0 : boolean;
  signal ptr_deref_2834_gather_scatter_ack_0 : boolean;
  signal binary_2877_inst_req_0 : boolean;
  signal ptr_deref_2834_gather_scatter_req_0 : boolean;
  signal ptr_deref_2892_addr_0_req_1 : boolean;
  signal ptr_deref_2834_load_3_ack_1 : boolean;
  signal ptr_deref_2899_store_0_ack_0 : boolean;
  signal binary_2863_inst_ack_0 : boolean;
  signal ptr_deref_2892_gather_scatter_req_0 : boolean;
  signal ptr_deref_2892_addr_0_ack_0 : boolean;
  signal ptr_deref_2834_addr_0_req_0 : boolean;
  signal ptr_deref_2904_addr_1_req_1 : boolean;
  signal ptr_deref_2834_load_0_req_1 : boolean;
  signal ptr_deref_2904_addr_3_req_0 : boolean;
  signal ptr_deref_2834_load_3_req_1 : boolean;
  signal ptr_deref_2899_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2892_addr_0_req_0 : boolean;
  signal ptr_deref_2834_load_0_ack_1 : boolean;
  signal call_stmt_2890_call_ack_0 : boolean;
  signal ptr_deref_2899_root_address_inst_ack_0 : boolean;
  signal binary_2877_inst_ack_1 : boolean;
  signal binary_2869_inst_req_0 : boolean;
  signal ptr_deref_2892_root_address_inst_req_0 : boolean;
  signal call_stmt_2897_call_req_1 : boolean;
  signal ptr_deref_2904_addr_1_req_0 : boolean;
  signal type_cast_2873_inst_req_0 : boolean;
  signal call_stmt_2890_call_req_1 : boolean;
  signal ptr_deref_2892_addr_1_req_0 : boolean;
  signal type_cast_2908_inst_req_0 : boolean;
  signal ptr_deref_2834_addr_2_req_1 : boolean;
  signal ptr_deref_2892_root_address_inst_ack_0 : boolean;
  signal call_stmt_2890_call_ack_1 : boolean;
  signal ptr_deref_2892_addr_1_ack_0 : boolean;
  signal type_cast_2908_inst_ack_0 : boolean;
  signal ptr_deref_2904_load_1_req_1 : boolean;
  signal binary_2869_inst_ack_0 : boolean;
  signal ptr_deref_2904_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2904_load_3_ack_1 : boolean;
  signal ptr_deref_2904_load_3_ack_0 : boolean;
  signal call_stmt_2897_call_ack_0 : boolean;
  signal type_cast_2873_inst_ack_0 : boolean;
  signal ptr_deref_2892_addr_1_req_1 : boolean;
  signal ptr_deref_2892_store_0_req_0 : boolean;
  signal ptr_deref_2904_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2834_load_1_req_0 : boolean;
  signal ptr_deref_2834_addr_2_ack_1 : boolean;
  signal ptr_deref_2904_addr_1_ack_0 : boolean;
  signal ptr_deref_2892_addr_1_ack_1 : boolean;
  signal ptr_deref_2904_load_0_ack_0 : boolean;
  signal ptr_deref_2892_store_0_ack_0 : boolean;
  signal ptr_deref_2904_load_2_req_1 : boolean;
  signal ptr_deref_2899_base_resize_req_0 : boolean;
  signal ptr_deref_2904_load_2_ack_1 : boolean;
  signal ptr_deref_2904_load_0_req_1 : boolean;
  signal ptr_deref_2904_addr_2_ack_1 : boolean;
  signal ptr_deref_2899_store_1_ack_0 : boolean;
  signal ptr_deref_2834_base_resize_req_0 : boolean;
  signal ptr_deref_2834_addr_3_ack_1 : boolean;
  signal ptr_deref_2834_load_2_ack_0 : boolean;
  signal call_stmt_2897_call_ack_1 : boolean;
  signal ptr_deref_2834_base_resize_ack_0 : boolean;
  signal ptr_deref_2834_root_address_inst_req_0 : boolean;
  signal ptr_deref_2834_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2834_load_1_ack_0 : boolean;
  signal type_cast_2916_inst_ack_0 : boolean;
  signal ptr_deref_2904_gather_scatter_req_0 : boolean;
  signal ptr_deref_2892_store_1_ack_0 : boolean;
  signal ptr_deref_2904_root_address_inst_req_0 : boolean;
  signal ptr_deref_2904_load_3_req_0 : boolean;
  signal simple_obj_ref_2914_inst_ack_0 : boolean;
  signal ptr_deref_2904_load_3_req_1 : boolean;
  signal type_cast_2916_inst_req_0 : boolean;
  signal simple_obj_ref_2914_inst_req_0 : boolean;
  signal binary_2886_inst_req_0 : boolean;
  signal ptr_deref_2899_store_0_req_0 : boolean;
  signal simple_obj_ref_2910_inst_ack_0 : boolean;
  signal ptr_deref_2899_addr_1_ack_1 : boolean;
  signal ptr_deref_2899_addr_1_req_1 : boolean;
  signal ptr_deref_2899_addr_1_ack_0 : boolean;
  signal ptr_deref_2899_addr_1_req_0 : boolean;
  signal ptr_deref_2899_addr_0_ack_1 : boolean;
  signal simple_obj_ref_2765_inst_req_0 : boolean;
  signal simple_obj_ref_2765_inst_ack_0 : boolean;
  signal ptr_deref_2892_store_1_req_0 : boolean;
  signal type_cast_2766_inst_req_0 : boolean;
  signal type_cast_2881_inst_ack_0 : boolean;
  signal type_cast_2766_inst_ack_0 : boolean;
  signal ptr_deref_2834_load_3_ack_0 : boolean;
  signal ptr_deref_2904_load_1_ack_0 : boolean;
  signal type_cast_2881_inst_req_0 : boolean;
  signal ptr_deref_2892_store_1_ack_1 : boolean;
  signal type_cast_2770_inst_req_0 : boolean;
  signal type_cast_2770_inst_ack_0 : boolean;
  signal ptr_deref_2892_store_1_req_1 : boolean;
  signal binary_2776_inst_req_0 : boolean;
  signal binary_2776_inst_ack_0 : boolean;
  signal binary_2776_inst_req_1 : boolean;
  signal binary_2776_inst_ack_1 : boolean;
  signal type_cast_2780_inst_req_0 : boolean;
  signal type_cast_2780_inst_ack_0 : boolean;
  signal call_stmt_2785_call_req_0 : boolean;
  signal call_stmt_2785_call_ack_0 : boolean;
  signal call_stmt_2785_call_req_1 : boolean;
  signal call_stmt_2785_call_ack_1 : boolean;
  signal ptr_deref_2787_base_resize_req_0 : boolean;
  signal ptr_deref_2787_base_resize_ack_0 : boolean;
  signal ptr_deref_2787_root_address_inst_req_0 : boolean;
  signal ptr_deref_2787_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2787_addr_0_req_0 : boolean;
  signal ptr_deref_2787_addr_0_ack_0 : boolean;
  signal ptr_deref_2787_addr_0_req_1 : boolean;
  signal ptr_deref_2787_addr_0_ack_1 : boolean;
  signal ptr_deref_2787_addr_1_req_0 : boolean;
  signal ptr_deref_2787_addr_1_ack_0 : boolean;
  signal ptr_deref_2787_addr_1_req_1 : boolean;
  signal ptr_deref_2787_addr_1_ack_1 : boolean;
  signal ptr_deref_2787_gather_scatter_req_0 : boolean;
  signal ptr_deref_2787_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2787_store_0_req_0 : boolean;
  signal ptr_deref_2787_store_0_ack_0 : boolean;
  signal ptr_deref_2787_store_1_req_0 : boolean;
  signal ptr_deref_2787_store_1_ack_0 : boolean;
  signal ptr_deref_2787_store_0_req_1 : boolean;
  signal ptr_deref_2787_store_0_ack_1 : boolean;
  signal ptr_deref_2787_store_1_req_1 : boolean;
  signal ptr_deref_2787_store_1_ack_1 : boolean;
  signal binary_2794_inst_req_0 : boolean;
  signal binary_2794_inst_ack_0 : boolean;
  signal binary_2794_inst_req_1 : boolean;
  signal binary_2794_inst_ack_1 : boolean;
  signal type_cast_2798_inst_req_0 : boolean;
  signal type_cast_2798_inst_ack_0 : boolean;
  signal binary_2804_inst_req_0 : boolean;
  signal binary_2804_inst_ack_0 : boolean;
  signal binary_2804_inst_req_1 : boolean;
  signal binary_2804_inst_ack_1 : boolean;
  signal ptr_deref_2904_addr_2_ack_0 : boolean;
  signal type_cast_2808_inst_req_0 : boolean;
  signal type_cast_2808_inst_ack_0 : boolean;
  signal array_obj_ref_2815_base_resize_req_0 : boolean;
  signal array_obj_ref_2815_base_resize_ack_0 : boolean;
  signal array_obj_ref_2815_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2815_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2815_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2815_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2815_final_reg_req_0 : boolean;
  signal array_obj_ref_2815_final_reg_ack_0 : boolean;
  signal ptr_deref_2819_base_resize_req_0 : boolean;
  signal ptr_deref_2819_base_resize_ack_0 : boolean;
  signal ptr_deref_2819_root_address_inst_req_0 : boolean;
  signal ptr_deref_2819_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2819_addr_0_req_0 : boolean;
  signal ptr_deref_2819_addr_0_ack_0 : boolean;
  signal ptr_deref_2819_addr_0_req_1 : boolean;
  signal ptr_deref_2819_addr_0_ack_1 : boolean;
  signal ptr_deref_2819_addr_1_req_0 : boolean;
  signal ptr_deref_2819_addr_1_ack_0 : boolean;
  signal ptr_deref_2819_addr_1_req_1 : boolean;
  signal ptr_deref_2819_addr_1_ack_1 : boolean;
  signal ptr_deref_2819_addr_2_req_0 : boolean;
  signal ptr_deref_2819_addr_2_ack_0 : boolean;
  signal ptr_deref_2819_addr_2_req_1 : boolean;
  signal ptr_deref_2819_addr_2_ack_1 : boolean;
  signal ptr_deref_2819_addr_3_req_0 : boolean;
  signal ptr_deref_2819_addr_3_ack_0 : boolean;
  signal ptr_deref_2819_addr_3_req_1 : boolean;
  signal ptr_deref_2819_addr_3_ack_1 : boolean;
  signal ptr_deref_2819_load_0_req_0 : boolean;
  signal ptr_deref_2819_load_0_ack_0 : boolean;
  signal ptr_deref_2819_load_1_req_0 : boolean;
  signal ptr_deref_2819_load_1_ack_0 : boolean;
  signal ptr_deref_2819_load_2_req_0 : boolean;
  signal ptr_deref_2819_load_2_ack_0 : boolean;
  signal ptr_deref_2819_load_3_req_0 : boolean;
  signal ptr_deref_2819_load_3_ack_0 : boolean;
  signal ptr_deref_2819_load_0_req_1 : boolean;
  signal ptr_deref_2819_load_0_ack_1 : boolean;
  signal ptr_deref_2819_load_1_req_1 : boolean;
  signal ptr_deref_2819_load_1_ack_1 : boolean;
  signal ptr_deref_2819_load_2_req_1 : boolean;
  signal ptr_deref_2819_load_2_ack_1 : boolean;
  signal ptr_deref_2819_load_3_req_1 : boolean;
  signal ptr_deref_2819_load_3_ack_1 : boolean;
  signal ptr_deref_2819_gather_scatter_req_0 : boolean;
  signal ptr_deref_2819_gather_scatter_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to2_CP_13690: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_13781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2785_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_14306_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_2890_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_14604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_2910_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13736_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2766_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_13731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2765_inst_req_0); -- 
    ack_13732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2765_inst_ack_0, ack => cp_elements(8)); -- 
    ack_13737_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2766_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2770_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_13750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2770_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2776_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_13760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2776_inst_ack_0, ack => cp_elements(18)); -- 
    cr_13761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2776_inst_req_1); -- 
    ca_13762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2776_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2780_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_13772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2780_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_13782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2785_call_ack_0, ack => cp_elements(24)); -- 
    ccr_13786_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2785_call_req_1); -- 
    cca_13787_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2785_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_13833_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2787_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_13806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2787_base_resize_req_0); -- 
    base_resize_ack_13807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_13811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2787_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2787_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_13819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2787_addr_0_req_0); -- 
    ra_13820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_13821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2787_addr_0_req_1); -- 
    ca_13822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_13826_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2787_addr_1_req_0); -- 
    ra_13827_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_13828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2787_addr_1_req_1); -- 
    ca_13829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2787_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_13841_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2787_store_0_req_0); -- 
    ra_13842_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_13846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2787_store_1_req_0); -- 
    ra_13847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_13857_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2787_store_0_req_1); -- 
    ca_13858_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_13862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2787_store_1_req_1); -- 
    ca_13863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2787_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13872_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2794_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_13873_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2794_inst_ack_0, ack => cp_elements(55)); -- 
    cr_13874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2794_inst_req_1); -- 
    ca_13875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2794_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2798_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_13885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2798_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_13894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2804_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_13895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2804_inst_ack_0, ack => cp_elements(63)); -- 
    cr_13896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2804_inst_req_1); -- 
    ca_13897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2804_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_13906_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2808_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_13907_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2808_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_13931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2815_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_13918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2815_base_resize_req_0); -- 
    base_resize_ack_13919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2815_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_13924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2815_root_address_inst_req_0); -- 
    plus_base_ra_13925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2815_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_13926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2815_root_address_inst_req_1); -- 
    plus_base_ca_13927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2815_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2815_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_13945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2819_base_resize_req_0); -- 
    base_resize_ack_13946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_13950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2819_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2819_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_13958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2819_addr_0_req_0); -- 
    ra_13959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_13960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2819_addr_0_req_1); -- 
    ca_13961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_13965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2819_addr_1_req_0); -- 
    ra_13966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_13967_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2819_addr_1_req_1); -- 
    ca_13968_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_13972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2819_addr_2_req_0); -- 
    ra_13973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_13974_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2819_addr_2_req_1); -- 
    ca_13975_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_13979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2819_addr_3_req_0); -- 
    ra_13980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_13981_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2819_addr_3_req_1); -- 
    ca_13982_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_13992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2819_load_0_req_0); -- 
    ra_13993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_13997_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2819_load_1_req_0); -- 
    ra_13998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_14002_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2819_load_2_req_0); -- 
    ra_14003_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_14007_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2819_load_3_req_0); -- 
    ra_14008_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_14018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2819_load_0_req_1); -- 
    ca_14019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_14023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2819_load_1_req_1); -- 
    ca_14024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_14028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2819_load_2_req_1); -- 
    ca_14029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_14033_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2819_load_3_req_1); -- 
    ca_14034_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_14035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2819_gather_scatter_req_0); -- 
    merge_ack_14036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2819_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14045_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2823_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_14046_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2823_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_14070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2830_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_14057_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2830_base_resize_req_0); -- 
    base_resize_ack_14058_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2830_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_14063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2830_root_address_inst_req_0); -- 
    plus_base_ra_14064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2830_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_14065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2830_root_address_inst_req_1); -- 
    plus_base_ca_14066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2830_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2830_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_14084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2834_base_resize_req_0); -- 
    base_resize_ack_14085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_14089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2834_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2834_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_14097_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2834_addr_0_req_0); -- 
    ra_14098_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_14099_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2834_addr_0_req_1); -- 
    ca_14100_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_14104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2834_addr_1_req_0); -- 
    ra_14105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_14106_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2834_addr_1_req_1); -- 
    ca_14107_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_14111_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2834_addr_2_req_0); -- 
    ra_14112_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_14113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2834_addr_2_req_1); -- 
    ca_14114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_14118_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2834_addr_3_req_0); -- 
    ra_14119_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_14120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2834_addr_3_req_1); -- 
    ca_14121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_14131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2834_load_0_req_0); -- 
    ra_14132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_14136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2834_load_1_req_0); -- 
    ra_14137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_14141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2834_load_2_req_0); -- 
    ra_14142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_14146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2834_load_3_req_0); -- 
    ra_14147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_14157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2834_load_0_req_1); -- 
    ca_14158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_14162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2834_load_1_req_1); -- 
    ca_14163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_14167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2834_load_2_req_1); -- 
    ca_14168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_14172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2834_load_3_req_1); -- 
    ca_14173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_14174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2834_gather_scatter_req_0); -- 
    merge_ack_14175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2834_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2838_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_14185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2838_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_2843_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_14196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2843_inst_ack_0, ack => cp_elements(162)); -- 
    cr_14197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_2843_inst_req_1); -- 
    cp_elements(163) <= binary_2843_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14207_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_2847_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_14208_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2847_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14217_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_2853_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_14218_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2853_inst_ack_0, ack => cp_elements(171)); -- 
    cr_14219_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_2853_inst_req_1); -- 
    ca_14220_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2853_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14229_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_2857_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_14230_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2857_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14239_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_2863_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_14240_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2863_inst_ack_0, ack => cp_elements(178)); -- 
    cr_14241_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_2863_inst_req_1); -- 
    ca_14242_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2863_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_2869_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_14252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2869_inst_ack_0, ack => cp_elements(183)); -- 
    cr_14253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_2869_inst_req_1); -- 
    ca_14254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2869_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_2877_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_2873_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_14266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2873_inst_ack_0, ack => cp_elements(189)); -- 
    ra_14271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2877_inst_ack_0, ack => cp_elements(190)); -- 
    cr_14272_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_2877_inst_req_1); -- 
    ca_14273_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2877_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14282_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_2881_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_14283_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2881_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14293_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_2886_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_14294_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2886_inst_ack_0, ack => cp_elements(197)); -- 
    cr_14295_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_2886_inst_req_1); -- 
    ca_14296_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2886_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_14307_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2890_call_ack_0, ack => cp_elements(200)); -- 
    ccr_14311_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_2890_call_req_1); -- 
    cca_14312_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2890_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_14358_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_2892_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_14331_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_2892_base_resize_req_0); -- 
    base_resize_ack_14332_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_14336_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_2892_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_2892_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_14344_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_2892_addr_0_req_0); -- 
    ra_14345_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_14346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_2892_addr_0_req_1); -- 
    ca_14347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_14351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_2892_addr_1_req_0); -- 
    ra_14352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_14353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_2892_addr_1_req_1); -- 
    ca_14354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_2892_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_14366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_2892_store_0_req_0); -- 
    ra_14367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_14371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_2892_store_1_req_0); -- 
    ra_14372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_14382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_2892_store_0_req_1); -- 
    ca_14383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_14387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_2892_store_1_req_1); -- 
    ca_14388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2892_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_14398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_2897_call_req_0); -- 
    cra_14399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2897_call_ack_0, ack => cp_elements(227)); -- 
    ccr_14403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_2897_call_req_1); -- 
    cca_14404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2897_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_14450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_2899_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_14423_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_2899_base_resize_req_0); -- 
    base_resize_ack_14424_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_14428_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_2899_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_2899_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_14436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_2899_addr_0_req_0); -- 
    ra_14437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_14438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_2899_addr_0_req_1); -- 
    ca_14439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_14443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_2899_addr_1_req_0); -- 
    ra_14444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_14445_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_2899_addr_1_req_1); -- 
    ca_14446_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_2899_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_14458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_2899_store_0_req_0); -- 
    ra_14459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_14463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_2899_store_1_req_0); -- 
    ra_14464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_14474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_2899_store_0_req_1); -- 
    ca_14475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_14479_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_2899_store_1_req_1); -- 
    ca_14480_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2899_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_14493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_2904_base_resize_req_0); -- 
    base_resize_ack_14494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_14498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_2904_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_2904_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_14506_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_2904_addr_0_req_0); -- 
    ra_14507_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_14508_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_2904_addr_0_req_1); -- 
    ca_14509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_14513_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_2904_addr_1_req_0); -- 
    ra_14514_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_14515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_2904_addr_1_req_1); -- 
    ca_14516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_14520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_2904_addr_2_req_0); -- 
    ra_14521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_14522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_2904_addr_2_req_1); -- 
    ca_14523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_14527_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_2904_addr_3_req_0); -- 
    ra_14528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_14529_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_2904_addr_3_req_1); -- 
    ca_14530_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_14540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_2904_load_0_req_0); -- 
    ra_14541_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_14545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_2904_load_1_req_0); -- 
    ra_14546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_14550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_2904_load_2_req_0); -- 
    ra_14551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_14555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_2904_load_3_req_0); -- 
    ra_14556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_14566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_2904_load_0_req_1); -- 
    ca_14567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_14571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_2904_load_1_req_1); -- 
    ca_14572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_14576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_2904_load_2_req_1); -- 
    ca_14577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_14581_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_2904_load_3_req_1); -- 
    ca_14582_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_14583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_2904_gather_scatter_req_0); -- 
    merge_ack_14584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2904_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_2908_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_14594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2908_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_14605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2910_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_2916_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_14618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2916_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_14623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_2914_inst_req_0); -- 
    pipe_wack_14624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2914_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2815_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2815_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2815_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2830_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2830_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2830_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_2878 : std_logic_vector(0 downto 0);
    signal ptr_deref_2787_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2787_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2787_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2787_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2819_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2819_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2819_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2819_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2819_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2834_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2834_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2834_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2834_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2834_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2892_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2892_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2892_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2899_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2899_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2899_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2904_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2904_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2765_wire : std_logic_vector(31 downto 0);
    signal tmp10_2820 : std_logic_vector(31 downto 0);
    signal tmp11_2824 : std_logic_vector(31 downto 0);
    signal tmp12_2831 : std_logic_vector(31 downto 0);
    signal tmp13_2835 : std_logic_vector(31 downto 0);
    signal tmp14_2839 : std_logic_vector(31 downto 0);
    signal tmp15_2844 : std_logic_vector(31 downto 0);
    signal tmp16_2848 : std_logic_vector(15 downto 0);
    signal tmp17_2854 : std_logic_vector(31 downto 0);
    signal tmp18_2864 : std_logic_vector(15 downto 0);
    signal tmp19_2870 : std_logic_vector(31 downto 0);
    signal tmp1_2771 : std_logic_vector(31 downto 0);
    signal tmp20_2882 : std_logic_vector(15 downto 0);
    signal tmp21_2887 : std_logic_vector(15 downto 0);
    signal tmp22_2890 : std_logic_vector(15 downto 0);
    signal tmp23_2897 : std_logic_vector(15 downto 0);
    signal tmp24_2905 : std_logic_vector(31 downto 0);
    signal tmp25_2909 : std_logic_vector(31 downto 0);
    signal tmp2_2777 : std_logic_vector(31 downto 0);
    signal tmp3_2781 : std_logic_vector(31 downto 0);
    signal tmp4_2785 : std_logic_vector(15 downto 0);
    signal tmp5_2795 : std_logic_vector(31 downto 0);
    signal tmp6_2799 : std_logic_vector(31 downto 0);
    signal tmp7_2805 : std_logic_vector(31 downto 0);
    signal tmp8_2809 : std_logic_vector(31 downto 0);
    signal tmp9_2816 : std_logic_vector(31 downto 0);
    signal tmp_2767 : std_logic_vector(31 downto 0);
    signal type_cast_2775_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2783_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2793_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2803_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2852_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2862_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2868_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2873_wire : std_logic_vector(31 downto 0);
    signal type_cast_2876_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2912_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2916_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_2858 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2815_final_offset <= "0000000000010000";
    array_obj_ref_2830_final_offset <= "0000000000001100";
    ptr_deref_2787_word_offset_0 <= "0000000000000000";
    ptr_deref_2787_word_offset_1 <= "0000000000000001";
    ptr_deref_2819_word_offset_0 <= "0000000000000000";
    ptr_deref_2819_word_offset_1 <= "0000000000000001";
    ptr_deref_2819_word_offset_2 <= "0000000000000010";
    ptr_deref_2819_word_offset_3 <= "0000000000000011";
    ptr_deref_2834_word_offset_0 <= "0000000000000000";
    ptr_deref_2834_word_offset_1 <= "0000000000000001";
    ptr_deref_2834_word_offset_2 <= "0000000000000010";
    ptr_deref_2834_word_offset_3 <= "0000000000000011";
    ptr_deref_2892_word_offset_0 <= "0000000000000000";
    ptr_deref_2892_word_offset_1 <= "0000000000000001";
    ptr_deref_2899_word_offset_0 <= "0000000000000000";
    ptr_deref_2899_word_offset_1 <= "0000000000000001";
    ptr_deref_2904_word_offset_0 <= "0000000000000000";
    ptr_deref_2904_word_offset_1 <= "0000000000000001";
    ptr_deref_2904_word_offset_2 <= "0000000000000010";
    ptr_deref_2904_word_offset_3 <= "0000000000000011";
    type_cast_2775_wire_constant <= "11111111111111111111100000000000";
    type_cast_2783_wire_constant <= "0000000000000100";
    type_cast_2793_wire_constant <= "00000000000000000000000000000110";
    type_cast_2803_wire_constant <= "00000000000000000000000000000010";
    type_cast_2852_wire_constant <= "00000000000000000000000000000011";
    type_cast_2862_wire_constant <= "0001111111111111";
    type_cast_2868_wire_constant <= "00000000000000000000000000000111";
    type_cast_2876_wire_constant <= "00000000000000000000000000000000";
    type_cast_2912_wire_constant <= "00000000000000000000000000000011";
    array_obj_ref_2815_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2771, dout => array_obj_ref_2815_resized_base_address, req => array_obj_ref_2815_base_resize_req_0, ack => array_obj_ref_2815_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2815_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2815_root_address, dout => tmp9_2816, req => array_obj_ref_2815_final_reg_req_0, ack => array_obj_ref_2815_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2830_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2771, dout => array_obj_ref_2830_resized_base_address, req => array_obj_ref_2830_base_resize_req_0, ack => array_obj_ref_2830_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2830_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2830_root_address, dout => tmp12_2831, req => array_obj_ref_2830_final_reg_req_0, ack => array_obj_ref_2830_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2787_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2781, dout => ptr_deref_2787_resized_base_address, req => ptr_deref_2787_base_resize_req_0, ack => ptr_deref_2787_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2819_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2816, dout => ptr_deref_2819_resized_base_address, req => ptr_deref_2819_base_resize_req_0, ack => ptr_deref_2819_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2834_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2831, dout => ptr_deref_2834_resized_base_address, req => ptr_deref_2834_base_resize_req_0, ack => ptr_deref_2834_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2892_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2799, dout => ptr_deref_2892_resized_base_address, req => ptr_deref_2892_base_resize_req_0, ack => ptr_deref_2892_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2899_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2809, dout => ptr_deref_2899_resized_base_address, req => ptr_deref_2899_base_resize_req_0, ack => ptr_deref_2899_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2904_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2831, dout => ptr_deref_2904_resized_base_address, req => ptr_deref_2904_base_resize_req_0, ack => ptr_deref_2904_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2766_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2765_wire, dout => tmp_2767, req => type_cast_2766_inst_req_0, ack => type_cast_2766_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2770_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2767, dout => tmp1_2771, req => type_cast_2770_inst_req_0, ack => type_cast_2770_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2780_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2777, dout => tmp3_2781, req => type_cast_2780_inst_req_0, ack => type_cast_2780_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2798_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2795, dout => tmp6_2799, req => type_cast_2798_inst_req_0, ack => type_cast_2798_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2808_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2805, dout => tmp8_2809, req => type_cast_2808_inst_req_0, ack => type_cast_2808_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2823_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2820, dout => tmp11_2824, req => type_cast_2823_inst_req_0, ack => type_cast_2823_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2838_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2835, dout => tmp14_2839, req => type_cast_2838_inst_req_0, ack => type_cast_2838_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2847_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_2844, dout => tmp16_2848, req => type_cast_2847_inst_req_0, ack => type_cast_2847_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2857_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_2854, dout => xx_xtrx_xi_2858, req => type_cast_2857_inst_req_0, ack => type_cast_2857_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2873_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_2870, dout => type_cast_2873_wire, req => type_cast_2873_inst_req_0, ack => type_cast_2873_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2881_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_2878, dout => tmp20_2882, req => type_cast_2881_inst_req_0, ack => type_cast_2881_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2908_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_2905, dout => tmp25_2909, req => type_cast_2908_inst_req_0, ack => type_cast_2908_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2916_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_2909, dout => type_cast_2916_wire, req => type_cast_2916_inst_req_0, ack => type_cast_2916_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2787_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2787_gather_scatter_ack_0 <= ptr_deref_2787_gather_scatter_req_0;
      aggregated_sig <= tmp4_2785;
      ptr_deref_2787_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2787_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2787_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2787_root_address_inst_ack_0 <= ptr_deref_2787_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2787_resized_base_address;
      ptr_deref_2787_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2819_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2819_gather_scatter_ack_0 <= ptr_deref_2819_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2819_data_3 & ptr_deref_2819_data_2 & ptr_deref_2819_data_1 & ptr_deref_2819_data_0;
      tmp10_2820 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2819_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2819_root_address_inst_ack_0 <= ptr_deref_2819_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2819_resized_base_address;
      ptr_deref_2819_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2834_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2834_gather_scatter_ack_0 <= ptr_deref_2834_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2834_data_3 & ptr_deref_2834_data_2 & ptr_deref_2834_data_1 & ptr_deref_2834_data_0;
      tmp13_2835 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2834_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2834_root_address_inst_ack_0 <= ptr_deref_2834_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2834_resized_base_address;
      ptr_deref_2834_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2892_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2892_gather_scatter_ack_0 <= ptr_deref_2892_gather_scatter_req_0;
      aggregated_sig <= tmp22_2890;
      ptr_deref_2892_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2892_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2892_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2892_root_address_inst_ack_0 <= ptr_deref_2892_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2892_resized_base_address;
      ptr_deref_2892_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2899_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2899_gather_scatter_ack_0 <= ptr_deref_2899_gather_scatter_req_0;
      aggregated_sig <= tmp23_2897;
      ptr_deref_2899_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2899_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2899_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2899_root_address_inst_ack_0 <= ptr_deref_2899_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2899_resized_base_address;
      ptr_deref_2899_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2904_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2904_gather_scatter_ack_0 <= ptr_deref_2904_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2904_data_3 & ptr_deref_2904_data_2 & ptr_deref_2904_data_1 & ptr_deref_2904_data_0;
      tmp24_2905 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2904_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2904_root_address_inst_ack_0 <= ptr_deref_2904_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2904_resized_base_address;
      ptr_deref_2904_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2815_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2815_resized_base_address;
      array_obj_ref_2815_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2815_root_address_inst_req_0,
          ackL => array_obj_ref_2815_root_address_inst_ack_0,
          reqR => array_obj_ref_2815_root_address_inst_req_1,
          ackR => array_obj_ref_2815_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2830_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2830_resized_base_address;
      array_obj_ref_2830_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2830_root_address_inst_req_0,
          ackL => array_obj_ref_2830_root_address_inst_ack_0,
          reqR => array_obj_ref_2830_root_address_inst_req_1,
          ackR => array_obj_ref_2830_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2776_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2767;
      tmp2_2777 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2776_inst_req_0,
          ackL => binary_2776_inst_ack_0,
          reqR => binary_2776_inst_req_1,
          ackR => binary_2776_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2794_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2777;
      tmp5_2795 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2794_inst_req_0,
          ackL => binary_2794_inst_ack_0,
          reqR => binary_2794_inst_req_1,
          ackR => binary_2794_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2804_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2777;
      tmp7_2805 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2804_inst_req_0,
          ackL => binary_2804_inst_ack_0,
          reqR => binary_2804_inst_req_1,
          ackR => binary_2804_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_2843_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2824 & tmp14_2839;
      tmp15_2844 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2843_inst_req_0,
          ackL => binary_2843_inst_ack_0,
          reqR => binary_2843_inst_req_1,
          ackR => binary_2843_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_2853_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2844;
      tmp17_2854 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2853_inst_req_0,
          ackL => binary_2853_inst_ack_0,
          reqR => binary_2853_inst_req_1,
          ackR => binary_2853_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_2863_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_2858;
      tmp18_2864 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2863_inst_req_0,
          ackL => binary_2863_inst_ack_0,
          reqR => binary_2863_inst_req_1,
          ackR => binary_2863_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_2869_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_2844;
      tmp19_2870 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2869_inst_req_0,
          ackL => binary_2869_inst_ack_0,
          reqR => binary_2869_inst_req_1,
          ackR => binary_2869_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_2877_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_2873_wire;
      notx_xx_xi_2878 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2877_inst_req_0,
          ackL => binary_2877_inst_ack_0,
          reqR => binary_2877_inst_req_1,
          ackR => binary_2877_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_2886_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_2864 & tmp20_2882;
      tmp21_2887 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2886_inst_req_0,
          ackL => binary_2886_inst_ack_0,
          reqR => binary_2886_inst_req_1,
          ackR => binary_2886_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2787_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2787_root_address;
      ptr_deref_2787_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2787_addr_0_req_0,
          ackL => ptr_deref_2787_addr_0_ack_0,
          reqR => ptr_deref_2787_addr_0_req_1,
          ackR => ptr_deref_2787_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2787_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2787_root_address;
      ptr_deref_2787_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2787_addr_1_req_0,
          ackL => ptr_deref_2787_addr_1_ack_0,
          reqR => ptr_deref_2787_addr_1_req_1,
          ackR => ptr_deref_2787_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2819_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2819_root_address;
      ptr_deref_2819_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2819_addr_0_req_0,
          ackL => ptr_deref_2819_addr_0_ack_0,
          reqR => ptr_deref_2819_addr_0_req_1,
          ackR => ptr_deref_2819_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2819_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2819_root_address;
      ptr_deref_2819_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2819_addr_1_req_0,
          ackL => ptr_deref_2819_addr_1_ack_0,
          reqR => ptr_deref_2819_addr_1_req_1,
          ackR => ptr_deref_2819_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2819_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2819_root_address;
      ptr_deref_2819_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2819_addr_2_req_0,
          ackL => ptr_deref_2819_addr_2_ack_0,
          reqR => ptr_deref_2819_addr_2_req_1,
          ackR => ptr_deref_2819_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2819_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2819_root_address;
      ptr_deref_2819_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2819_addr_3_req_0,
          ackL => ptr_deref_2819_addr_3_ack_0,
          reqR => ptr_deref_2819_addr_3_req_1,
          ackR => ptr_deref_2819_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2834_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2834_root_address;
      ptr_deref_2834_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2834_addr_0_req_0,
          ackL => ptr_deref_2834_addr_0_ack_0,
          reqR => ptr_deref_2834_addr_0_req_1,
          ackR => ptr_deref_2834_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2834_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2834_root_address;
      ptr_deref_2834_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2834_addr_1_req_0,
          ackL => ptr_deref_2834_addr_1_ack_0,
          reqR => ptr_deref_2834_addr_1_req_1,
          ackR => ptr_deref_2834_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2834_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2834_root_address;
      ptr_deref_2834_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2834_addr_2_req_0,
          ackL => ptr_deref_2834_addr_2_ack_0,
          reqR => ptr_deref_2834_addr_2_req_1,
          ackR => ptr_deref_2834_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2834_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2834_root_address;
      ptr_deref_2834_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2834_addr_3_req_0,
          ackL => ptr_deref_2834_addr_3_ack_0,
          reqR => ptr_deref_2834_addr_3_req_1,
          ackR => ptr_deref_2834_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_2892_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2892_root_address;
      ptr_deref_2892_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2892_addr_0_req_0,
          ackL => ptr_deref_2892_addr_0_ack_0,
          reqR => ptr_deref_2892_addr_0_req_1,
          ackR => ptr_deref_2892_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_2892_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2892_root_address;
      ptr_deref_2892_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2892_addr_1_req_0,
          ackL => ptr_deref_2892_addr_1_ack_0,
          reqR => ptr_deref_2892_addr_1_req_1,
          ackR => ptr_deref_2892_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_2899_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2899_root_address;
      ptr_deref_2899_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2899_addr_0_req_0,
          ackL => ptr_deref_2899_addr_0_ack_0,
          reqR => ptr_deref_2899_addr_0_req_1,
          ackR => ptr_deref_2899_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_2899_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2899_root_address;
      ptr_deref_2899_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2899_addr_1_req_0,
          ackL => ptr_deref_2899_addr_1_ack_0,
          reqR => ptr_deref_2899_addr_1_req_1,
          ackR => ptr_deref_2899_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_2904_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_0_req_0,
          ackL => ptr_deref_2904_addr_0_ack_0,
          reqR => ptr_deref_2904_addr_0_req_1,
          ackR => ptr_deref_2904_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_2904_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_1_req_0,
          ackL => ptr_deref_2904_addr_1_ack_0,
          reqR => ptr_deref_2904_addr_1_req_1,
          ackR => ptr_deref_2904_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_2904_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_2_req_0,
          ackL => ptr_deref_2904_addr_2_ack_0,
          reqR => ptr_deref_2904_addr_2_req_1,
          ackR => ptr_deref_2904_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_2904_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2904_root_address;
      ptr_deref_2904_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2904_addr_3_req_0,
          ackL => ptr_deref_2904_addr_3_ack_0,
          reqR => ptr_deref_2904_addr_3_req_1,
          ackR => ptr_deref_2904_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2819_load_0 ptr_deref_2819_load_1 ptr_deref_2819_load_2 ptr_deref_2819_load_3 ptr_deref_2834_load_0 ptr_deref_2834_load_1 ptr_deref_2834_load_2 ptr_deref_2834_load_3 ptr_deref_2904_load_0 ptr_deref_2904_load_1 ptr_deref_2904_load_2 ptr_deref_2904_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2819_load_0_req_0,
        ptr_deref_2819_load_0_ack_0,
        ptr_deref_2819_load_0_req_1,
        ptr_deref_2819_load_0_ack_1,
        "ptr_deref_2819_load_0",
        "memory_space_5" ,
        ptr_deref_2819_data_0,
        ptr_deref_2819_word_address_0,
        "ptr_deref_2819_data_0",
        "ptr_deref_2819_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2819_load_1_req_0,
        ptr_deref_2819_load_1_ack_0,
        ptr_deref_2819_load_1_req_1,
        ptr_deref_2819_load_1_ack_1,
        "ptr_deref_2819_load_1",
        "memory_space_5" ,
        ptr_deref_2819_data_1,
        ptr_deref_2819_word_address_1,
        "ptr_deref_2819_data_1",
        "ptr_deref_2819_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2819_load_2_req_0,
        ptr_deref_2819_load_2_ack_0,
        ptr_deref_2819_load_2_req_1,
        ptr_deref_2819_load_2_ack_1,
        "ptr_deref_2819_load_2",
        "memory_space_5" ,
        ptr_deref_2819_data_2,
        ptr_deref_2819_word_address_2,
        "ptr_deref_2819_data_2",
        "ptr_deref_2819_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2819_load_3_req_0,
        ptr_deref_2819_load_3_ack_0,
        ptr_deref_2819_load_3_req_1,
        ptr_deref_2819_load_3_ack_1,
        "ptr_deref_2819_load_3",
        "memory_space_5" ,
        ptr_deref_2819_data_3,
        ptr_deref_2819_word_address_3,
        "ptr_deref_2819_data_3",
        "ptr_deref_2819_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2834_load_0_req_0,
        ptr_deref_2834_load_0_ack_0,
        ptr_deref_2834_load_0_req_1,
        ptr_deref_2834_load_0_ack_1,
        "ptr_deref_2834_load_0",
        "memory_space_5" ,
        ptr_deref_2834_data_0,
        ptr_deref_2834_word_address_0,
        "ptr_deref_2834_data_0",
        "ptr_deref_2834_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2834_load_1_req_0,
        ptr_deref_2834_load_1_ack_0,
        ptr_deref_2834_load_1_req_1,
        ptr_deref_2834_load_1_ack_1,
        "ptr_deref_2834_load_1",
        "memory_space_5" ,
        ptr_deref_2834_data_1,
        ptr_deref_2834_word_address_1,
        "ptr_deref_2834_data_1",
        "ptr_deref_2834_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2834_load_2_req_0,
        ptr_deref_2834_load_2_ack_0,
        ptr_deref_2834_load_2_req_1,
        ptr_deref_2834_load_2_ack_1,
        "ptr_deref_2834_load_2",
        "memory_space_5" ,
        ptr_deref_2834_data_2,
        ptr_deref_2834_word_address_2,
        "ptr_deref_2834_data_2",
        "ptr_deref_2834_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2834_load_3_req_0,
        ptr_deref_2834_load_3_ack_0,
        ptr_deref_2834_load_3_req_1,
        ptr_deref_2834_load_3_ack_1,
        "ptr_deref_2834_load_3",
        "memory_space_5" ,
        ptr_deref_2834_data_3,
        ptr_deref_2834_word_address_3,
        "ptr_deref_2834_data_3",
        "ptr_deref_2834_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2904_load_0_req_0,
        ptr_deref_2904_load_0_ack_0,
        ptr_deref_2904_load_0_req_1,
        ptr_deref_2904_load_0_ack_1,
        "ptr_deref_2904_load_0",
        "memory_space_5" ,
        ptr_deref_2904_data_0,
        ptr_deref_2904_word_address_0,
        "ptr_deref_2904_data_0",
        "ptr_deref_2904_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2904_load_1_req_0,
        ptr_deref_2904_load_1_ack_0,
        ptr_deref_2904_load_1_req_1,
        ptr_deref_2904_load_1_ack_1,
        "ptr_deref_2904_load_1",
        "memory_space_5" ,
        ptr_deref_2904_data_1,
        ptr_deref_2904_word_address_1,
        "ptr_deref_2904_data_1",
        "ptr_deref_2904_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2904_load_2_req_0,
        ptr_deref_2904_load_2_ack_0,
        ptr_deref_2904_load_2_req_1,
        ptr_deref_2904_load_2_ack_1,
        "ptr_deref_2904_load_2",
        "memory_space_5" ,
        ptr_deref_2904_data_2,
        ptr_deref_2904_word_address_2,
        "ptr_deref_2904_data_2",
        "ptr_deref_2904_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2904_load_3_req_0,
        ptr_deref_2904_load_3_ack_0,
        ptr_deref_2904_load_3_req_1,
        ptr_deref_2904_load_3_ack_1,
        "ptr_deref_2904_load_3",
        "memory_space_5" ,
        ptr_deref_2904_data_3,
        ptr_deref_2904_word_address_3,
        "ptr_deref_2904_data_3",
        "ptr_deref_2904_word_address_3" -- 
      );
      reqL(11) <= ptr_deref_2819_load_0_req_0;
      reqL(10) <= ptr_deref_2819_load_1_req_0;
      reqL(9) <= ptr_deref_2819_load_2_req_0;
      reqL(8) <= ptr_deref_2819_load_3_req_0;
      reqL(7) <= ptr_deref_2834_load_0_req_0;
      reqL(6) <= ptr_deref_2834_load_1_req_0;
      reqL(5) <= ptr_deref_2834_load_2_req_0;
      reqL(4) <= ptr_deref_2834_load_3_req_0;
      reqL(3) <= ptr_deref_2904_load_0_req_0;
      reqL(2) <= ptr_deref_2904_load_1_req_0;
      reqL(1) <= ptr_deref_2904_load_2_req_0;
      reqL(0) <= ptr_deref_2904_load_3_req_0;
      ptr_deref_2819_load_0_ack_0 <= ackL(11);
      ptr_deref_2819_load_1_ack_0 <= ackL(10);
      ptr_deref_2819_load_2_ack_0 <= ackL(9);
      ptr_deref_2819_load_3_ack_0 <= ackL(8);
      ptr_deref_2834_load_0_ack_0 <= ackL(7);
      ptr_deref_2834_load_1_ack_0 <= ackL(6);
      ptr_deref_2834_load_2_ack_0 <= ackL(5);
      ptr_deref_2834_load_3_ack_0 <= ackL(4);
      ptr_deref_2904_load_0_ack_0 <= ackL(3);
      ptr_deref_2904_load_1_ack_0 <= ackL(2);
      ptr_deref_2904_load_2_ack_0 <= ackL(1);
      ptr_deref_2904_load_3_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2819_load_0_req_1;
      reqR(10) <= ptr_deref_2819_load_1_req_1;
      reqR(9) <= ptr_deref_2819_load_2_req_1;
      reqR(8) <= ptr_deref_2819_load_3_req_1;
      reqR(7) <= ptr_deref_2834_load_0_req_1;
      reqR(6) <= ptr_deref_2834_load_1_req_1;
      reqR(5) <= ptr_deref_2834_load_2_req_1;
      reqR(4) <= ptr_deref_2834_load_3_req_1;
      reqR(3) <= ptr_deref_2904_load_0_req_1;
      reqR(2) <= ptr_deref_2904_load_1_req_1;
      reqR(1) <= ptr_deref_2904_load_2_req_1;
      reqR(0) <= ptr_deref_2904_load_3_req_1;
      ptr_deref_2819_load_0_ack_1 <= ackR(11);
      ptr_deref_2819_load_1_ack_1 <= ackR(10);
      ptr_deref_2819_load_2_ack_1 <= ackR(9);
      ptr_deref_2819_load_3_ack_1 <= ackR(8);
      ptr_deref_2834_load_0_ack_1 <= ackR(7);
      ptr_deref_2834_load_1_ack_1 <= ackR(6);
      ptr_deref_2834_load_2_ack_1 <= ackR(5);
      ptr_deref_2834_load_3_ack_1 <= ackR(4);
      ptr_deref_2904_load_0_ack_1 <= ackR(3);
      ptr_deref_2904_load_1_ack_1 <= ackR(2);
      ptr_deref_2904_load_2_ack_1 <= ackR(1);
      ptr_deref_2904_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_2819_word_address_0 & ptr_deref_2819_word_address_1 & ptr_deref_2819_word_address_2 & ptr_deref_2819_word_address_3 & ptr_deref_2834_word_address_0 & ptr_deref_2834_word_address_1 & ptr_deref_2834_word_address_2 & ptr_deref_2834_word_address_3 & ptr_deref_2904_word_address_0 & ptr_deref_2904_word_address_1 & ptr_deref_2904_word_address_2 & ptr_deref_2904_word_address_3;
      ptr_deref_2819_data_0 <= data_out(95 downto 88);
      ptr_deref_2819_data_1 <= data_out(87 downto 80);
      ptr_deref_2819_data_2 <= data_out(79 downto 72);
      ptr_deref_2819_data_3 <= data_out(71 downto 64);
      ptr_deref_2834_data_0 <= data_out(63 downto 56);
      ptr_deref_2834_data_1 <= data_out(55 downto 48);
      ptr_deref_2834_data_2 <= data_out(47 downto 40);
      ptr_deref_2834_data_3 <= data_out(39 downto 32);
      ptr_deref_2904_data_0 <= data_out(31 downto 24);
      ptr_deref_2904_data_1 <= data_out(23 downto 16);
      ptr_deref_2904_data_2 <= data_out(15 downto 8);
      ptr_deref_2904_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2787_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2787_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2787_word_address_0) &  " data ptr_deref_2787_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2787_data_0) severity note; --
        end if;
        if ptr_deref_2787_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2787_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2787_word_address_1) &  " data ptr_deref_2787_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2787_data_1) severity note; --
        end if;
        if ptr_deref_2892_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2892_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2892_word_address_0) &  " data ptr_deref_2892_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2892_data_0) severity note; --
        end if;
        if ptr_deref_2892_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2892_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2892_word_address_1) &  " data ptr_deref_2892_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2892_data_1) severity note; --
        end if;
        if ptr_deref_2899_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2899_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2899_word_address_0) &  " data ptr_deref_2899_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2899_data_0) severity note; --
        end if;
        if ptr_deref_2899_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2899_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2899_word_address_1) &  " data ptr_deref_2899_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2899_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2787_store_0 ptr_deref_2787_store_1 ptr_deref_2892_store_0 ptr_deref_2892_store_1 ptr_deref_2899_store_0 ptr_deref_2899_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2787_store_0_req_0;
      reqL(4) <= ptr_deref_2787_store_1_req_0;
      reqL(3) <= ptr_deref_2892_store_0_req_0;
      reqL(2) <= ptr_deref_2892_store_1_req_0;
      reqL(1) <= ptr_deref_2899_store_0_req_0;
      reqL(0) <= ptr_deref_2899_store_1_req_0;
      ptr_deref_2787_store_0_ack_0 <= ackL(5);
      ptr_deref_2787_store_1_ack_0 <= ackL(4);
      ptr_deref_2892_store_0_ack_0 <= ackL(3);
      ptr_deref_2892_store_1_ack_0 <= ackL(2);
      ptr_deref_2899_store_0_ack_0 <= ackL(1);
      ptr_deref_2899_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2787_store_0_req_1;
      reqR(4) <= ptr_deref_2787_store_1_req_1;
      reqR(3) <= ptr_deref_2892_store_0_req_1;
      reqR(2) <= ptr_deref_2892_store_1_req_1;
      reqR(1) <= ptr_deref_2899_store_0_req_1;
      reqR(0) <= ptr_deref_2899_store_1_req_1;
      ptr_deref_2787_store_0_ack_1 <= ackR(5);
      ptr_deref_2787_store_1_ack_1 <= ackR(4);
      ptr_deref_2892_store_0_ack_1 <= ackR(3);
      ptr_deref_2892_store_1_ack_1 <= ackR(2);
      ptr_deref_2899_store_0_ack_1 <= ackR(1);
      ptr_deref_2899_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2787_word_address_0 & ptr_deref_2787_word_address_1 & ptr_deref_2892_word_address_0 & ptr_deref_2892_word_address_1 & ptr_deref_2899_word_address_0 & ptr_deref_2899_word_address_1;
      data_in <= ptr_deref_2787_data_0 & ptr_deref_2787_data_1 & ptr_deref_2892_data_0 & ptr_deref_2892_data_1 & ptr_deref_2899_data_0 & ptr_deref_2899_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2765_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2765_inst_ack_0 then -- 
            assert false report " ReadPipe to2_in0 to wire simple_obj_ref_2765_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2765_inst_req_0;
      simple_obj_ref_2765_inst_ack_0 <= ack(0);
      simple_obj_ref_2765_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to2_in0_pipe_read_req(0),
          oack => to2_in0_pipe_read_ack(0),
          odata => to2_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2910_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_2912_wire_constant value="  &  convert_slv_to_hex_string(type_cast_2912_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_2910_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2910_inst_req_0;
      simple_obj_ref_2910_inst_ack_0 <= ack(0);
      data_in <= type_cast_2912_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_2914_inst_ack_0 then -- 
          assert false report " WritePipe tofpga2_out0 from wire type_cast_2916_wire value="  &  convert_slv_to_hex_string(type_cast_2916_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_2914_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_2914_inst_req_0;
      simple_obj_ref_2914_inst_ack_0 <= ack(0);
      data_in <= type_cast_2916_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga2_out0_pipe_write_req(0),
          oack => tofpga2_out0_pipe_write_ack(0),
          odata => tofpga2_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2785_call call_stmt_2890_call call_stmt_2897_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2785_call_req_0;
      reqL(1) <= call_stmt_2890_call_req_0;
      reqL(0) <= call_stmt_2897_call_req_0;
      call_stmt_2785_call_ack_0 <= ackL(2);
      call_stmt_2890_call_ack_0 <= ackL(1);
      call_stmt_2897_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2785_call_req_1;
      reqR(1) <= call_stmt_2890_call_req_1;
      reqR(0) <= call_stmt_2897_call_req_1;
      call_stmt_2785_call_ack_1 <= ackR(2);
      call_stmt_2890_call_ack_1 <= ackR(1);
      call_stmt_2897_call_ack_1 <= ackR(0);
      data_in <= type_cast_2783_wire_constant & tmp16_2848 & tmp21_2887;
      tmp4_2785 <= data_out(47 downto 32);
      tmp22_2890 <= data_out(31 downto 16);
      tmp23_2897 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_glue_to3 is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    to3_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
    to3_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    to3_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga3_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
    ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
    ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
    ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
    ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity ahir_glue_to3;
architecture Default of ahir_glue_to3 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal ahir_glue_to3_CP_14633_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3064_addr_0_req_1 : boolean;
  signal binary_3037_inst_req_0 : boolean;
  signal ptr_deref_3052_store_1_req_1 : boolean;
  signal type_cast_3041_inst_ack_0 : boolean;
  signal binary_3023_inst_ack_1 : boolean;
  signal binary_3037_inst_ack_1 : boolean;
  signal ptr_deref_3059_addr_1_ack_1 : boolean;
  signal binary_3023_inst_req_1 : boolean;
  signal binary_3037_inst_req_1 : boolean;
  signal ptr_deref_3059_store_0_req_1 : boolean;
  signal ptr_deref_3064_addr_1_ack_1 : boolean;
  signal binary_3029_inst_ack_0 : boolean;
  signal ptr_deref_3059_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3064_addr_1_req_1 : boolean;
  signal ptr_deref_3059_addr_1_req_1 : boolean;
  signal ptr_deref_3064_addr_0_ack_0 : boolean;
  signal binary_3037_inst_ack_0 : boolean;
  signal ptr_deref_3064_load_0_req_0 : boolean;
  signal ptr_deref_3064_load_2_req_1 : boolean;
  signal ptr_deref_3059_addr_0_req_0 : boolean;
  signal ptr_deref_3052_store_1_ack_0 : boolean;
  signal ptr_deref_3059_addr_1_ack_0 : boolean;
  signal ptr_deref_3064_load_1_ack_0 : boolean;
  signal ptr_deref_3064_load_3_ack_1 : boolean;
  signal ptr_deref_3064_load_2_req_0 : boolean;
  signal ptr_deref_3059_store_0_ack_1 : boolean;
  signal ptr_deref_3064_addr_0_ack_1 : boolean;
  signal ptr_deref_3059_store_1_req_1 : boolean;
  signal simple_obj_ref_3070_inst_req_0 : boolean;
  signal ptr_deref_3064_addr_3_ack_0 : boolean;
  signal ptr_deref_3064_gather_scatter_req_0 : boolean;
  signal ptr_deref_3064_addr_1_req_0 : boolean;
  signal ptr_deref_3059_store_1_ack_1 : boolean;
  signal ptr_deref_3064_addr_0_req_0 : boolean;
  signal call_stmt_3057_call_req_0 : boolean;
  signal binary_3029_inst_req_0 : boolean;
  signal ptr_deref_3064_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3064_load_1_req_0 : boolean;
  signal type_cast_3068_inst_ack_0 : boolean;
  signal type_cast_3068_inst_req_0 : boolean;
  signal ptr_deref_3052_base_resize_req_0 : boolean;
  signal simple_obj_ref_3070_inst_ack_0 : boolean;
  signal ptr_deref_3052_store_1_req_0 : boolean;
  signal ptr_deref_3059_gather_scatter_req_0 : boolean;
  signal ptr_deref_3052_store_0_ack_1 : boolean;
  signal ptr_deref_3064_load_2_ack_1 : boolean;
  signal binary_3046_inst_req_0 : boolean;
  signal ptr_deref_3052_gather_scatter_ack_0 : boolean;
  signal binary_3029_inst_req_1 : boolean;
  signal binary_3029_inst_ack_1 : boolean;
  signal call_stmt_3057_call_ack_1 : boolean;
  signal call_stmt_3057_call_ack_0 : boolean;
  signal ptr_deref_3052_store_0_req_0 : boolean;
  signal binary_3046_inst_req_1 : boolean;
  signal call_stmt_3057_call_req_1 : boolean;
  signal binary_3023_inst_req_0 : boolean;
  signal type_cast_3033_inst_ack_0 : boolean;
  signal ptr_deref_3064_addr_2_req_0 : boolean;
  signal ptr_deref_3052_base_resize_ack_0 : boolean;
  signal call_stmt_3050_call_req_0 : boolean;
  signal type_cast_3041_inst_req_0 : boolean;
  signal ptr_deref_3059_addr_0_req_1 : boolean;
  signal ptr_deref_3052_root_address_inst_req_0 : boolean;
  signal binary_3023_inst_ack_0 : boolean;
  signal binary_3046_inst_ack_0 : boolean;
  signal simple_obj_ref_3074_inst_req_0 : boolean;
  signal ptr_deref_3064_addr_1_ack_0 : boolean;
  signal ptr_deref_3059_addr_0_ack_1 : boolean;
  signal ptr_deref_3052_store_1_ack_1 : boolean;
  signal ptr_deref_3064_load_0_ack_1 : boolean;
  signal ptr_deref_3059_addr_0_ack_0 : boolean;
  signal ptr_deref_3059_addr_1_req_0 : boolean;
  signal ptr_deref_3052_root_address_inst_ack_0 : boolean;
  signal type_cast_3033_inst_req_0 : boolean;
  signal ptr_deref_3064_load_2_ack_0 : boolean;
  signal ptr_deref_3064_addr_2_ack_0 : boolean;
  signal call_stmt_3050_call_ack_0 : boolean;
  signal ptr_deref_3064_addr_2_req_1 : boolean;
  signal call_stmt_3050_call_req_1 : boolean;
  signal call_stmt_3050_call_ack_1 : boolean;
  signal ptr_deref_3064_base_resize_req_0 : boolean;
  signal ptr_deref_3064_base_resize_ack_0 : boolean;
  signal ptr_deref_3052_store_0_req_1 : boolean;
  signal ptr_deref_3059_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3064_root_address_inst_req_0 : boolean;
  signal ptr_deref_3064_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3064_addr_2_ack_1 : boolean;
  signal binary_3046_inst_ack_1 : boolean;
  signal ptr_deref_3064_load_0_ack_0 : boolean;
  signal ptr_deref_3059_store_0_req_0 : boolean;
  signal ptr_deref_3059_store_0_ack_0 : boolean;
  signal ptr_deref_3059_base_resize_req_0 : boolean;
  signal ptr_deref_3064_load_1_req_1 : boolean;
  signal ptr_deref_3059_base_resize_ack_0 : boolean;
  signal ptr_deref_3064_addr_3_req_0 : boolean;
  signal simple_obj_ref_3074_inst_ack_0 : boolean;
  signal ptr_deref_3064_load_3_req_0 : boolean;
  signal ptr_deref_3064_load_3_ack_0 : boolean;
  signal ptr_deref_3052_addr_0_req_0 : boolean;
  signal ptr_deref_3052_addr_0_ack_0 : boolean;
  signal ptr_deref_3064_load_0_req_1 : boolean;
  signal ptr_deref_3064_addr_3_req_1 : boolean;
  signal ptr_deref_3052_addr_0_req_1 : boolean;
  signal ptr_deref_3064_addr_3_ack_1 : boolean;
  signal type_cast_3076_inst_ack_0 : boolean;
  signal type_cast_3076_inst_req_0 : boolean;
  signal ptr_deref_3064_load_1_ack_1 : boolean;
  signal ptr_deref_3052_addr_0_ack_1 : boolean;
  signal ptr_deref_3059_store_1_req_0 : boolean;
  signal ptr_deref_3052_store_0_ack_0 : boolean;
  signal ptr_deref_3052_addr_1_req_0 : boolean;
  signal ptr_deref_3052_addr_1_ack_0 : boolean;
  signal ptr_deref_3052_addr_1_req_1 : boolean;
  signal ptr_deref_3059_store_1_ack_0 : boolean;
  signal ptr_deref_3052_addr_1_ack_1 : boolean;
  signal ptr_deref_3059_root_address_inst_req_0 : boolean;
  signal ptr_deref_3064_load_3_req_1 : boolean;
  signal ptr_deref_3052_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_2925_inst_req_0 : boolean;
  signal simple_obj_ref_2925_inst_ack_0 : boolean;
  signal type_cast_2926_inst_req_0 : boolean;
  signal type_cast_2926_inst_ack_0 : boolean;
  signal type_cast_2930_inst_req_0 : boolean;
  signal type_cast_2930_inst_ack_0 : boolean;
  signal binary_2936_inst_req_0 : boolean;
  signal binary_2936_inst_ack_0 : boolean;
  signal binary_2936_inst_req_1 : boolean;
  signal binary_2936_inst_ack_1 : boolean;
  signal type_cast_2940_inst_req_0 : boolean;
  signal type_cast_2940_inst_ack_0 : boolean;
  signal call_stmt_2945_call_req_0 : boolean;
  signal call_stmt_2945_call_ack_0 : boolean;
  signal call_stmt_2945_call_req_1 : boolean;
  signal call_stmt_2945_call_ack_1 : boolean;
  signal ptr_deref_2947_base_resize_req_0 : boolean;
  signal ptr_deref_2947_base_resize_ack_0 : boolean;
  signal ptr_deref_2947_root_address_inst_req_0 : boolean;
  signal ptr_deref_2947_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2947_addr_0_req_0 : boolean;
  signal ptr_deref_2947_addr_0_ack_0 : boolean;
  signal ptr_deref_2947_addr_0_req_1 : boolean;
  signal ptr_deref_2947_addr_0_ack_1 : boolean;
  signal ptr_deref_2947_addr_1_req_0 : boolean;
  signal ptr_deref_2947_addr_1_ack_0 : boolean;
  signal ptr_deref_2947_addr_1_req_1 : boolean;
  signal ptr_deref_2947_addr_1_ack_1 : boolean;
  signal ptr_deref_2947_gather_scatter_req_0 : boolean;
  signal ptr_deref_2947_gather_scatter_ack_0 : boolean;
  signal ptr_deref_2947_store_0_req_0 : boolean;
  signal ptr_deref_2947_store_0_ack_0 : boolean;
  signal ptr_deref_2947_store_1_req_0 : boolean;
  signal ptr_deref_2947_store_1_ack_0 : boolean;
  signal ptr_deref_2947_store_0_req_1 : boolean;
  signal ptr_deref_2947_store_0_ack_1 : boolean;
  signal ptr_deref_2947_store_1_req_1 : boolean;
  signal ptr_deref_2947_store_1_ack_1 : boolean;
  signal binary_2954_inst_req_0 : boolean;
  signal binary_2954_inst_ack_0 : boolean;
  signal binary_2954_inst_req_1 : boolean;
  signal binary_2954_inst_ack_1 : boolean;
  signal type_cast_2958_inst_req_0 : boolean;
  signal type_cast_2958_inst_ack_0 : boolean;
  signal binary_2964_inst_req_0 : boolean;
  signal binary_2964_inst_ack_0 : boolean;
  signal binary_2964_inst_req_1 : boolean;
  signal binary_2964_inst_ack_1 : boolean;
  signal type_cast_2968_inst_req_0 : boolean;
  signal type_cast_2968_inst_ack_0 : boolean;
  signal array_obj_ref_2975_base_resize_req_0 : boolean;
  signal array_obj_ref_2975_base_resize_ack_0 : boolean;
  signal array_obj_ref_2975_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2975_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2975_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2975_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2975_final_reg_req_0 : boolean;
  signal array_obj_ref_2975_final_reg_ack_0 : boolean;
  signal ptr_deref_2979_base_resize_req_0 : boolean;
  signal ptr_deref_2979_base_resize_ack_0 : boolean;
  signal ptr_deref_2979_root_address_inst_req_0 : boolean;
  signal ptr_deref_2979_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2979_addr_0_req_0 : boolean;
  signal ptr_deref_2979_addr_0_ack_0 : boolean;
  signal ptr_deref_2979_addr_0_req_1 : boolean;
  signal ptr_deref_2979_addr_0_ack_1 : boolean;
  signal ptr_deref_2979_addr_1_req_0 : boolean;
  signal ptr_deref_2979_addr_1_ack_0 : boolean;
  signal ptr_deref_2979_addr_1_req_1 : boolean;
  signal ptr_deref_2979_addr_1_ack_1 : boolean;
  signal ptr_deref_2979_addr_2_req_0 : boolean;
  signal ptr_deref_2979_addr_2_ack_0 : boolean;
  signal ptr_deref_2979_addr_2_req_1 : boolean;
  signal ptr_deref_2979_addr_2_ack_1 : boolean;
  signal ptr_deref_2979_addr_3_req_0 : boolean;
  signal ptr_deref_2979_addr_3_ack_0 : boolean;
  signal ptr_deref_2979_addr_3_req_1 : boolean;
  signal ptr_deref_2979_addr_3_ack_1 : boolean;
  signal ptr_deref_2979_load_0_req_0 : boolean;
  signal ptr_deref_2979_load_0_ack_0 : boolean;
  signal ptr_deref_2979_load_1_req_0 : boolean;
  signal ptr_deref_2979_load_1_ack_0 : boolean;
  signal ptr_deref_2979_load_2_req_0 : boolean;
  signal ptr_deref_2979_load_2_ack_0 : boolean;
  signal ptr_deref_2979_load_3_req_0 : boolean;
  signal ptr_deref_2979_load_3_ack_0 : boolean;
  signal ptr_deref_2979_load_0_req_1 : boolean;
  signal ptr_deref_2979_load_0_ack_1 : boolean;
  signal ptr_deref_2979_load_1_req_1 : boolean;
  signal ptr_deref_2979_load_1_ack_1 : boolean;
  signal ptr_deref_2979_load_2_req_1 : boolean;
  signal ptr_deref_2979_load_2_ack_1 : boolean;
  signal ptr_deref_2979_load_3_req_1 : boolean;
  signal ptr_deref_2979_load_3_ack_1 : boolean;
  signal ptr_deref_2979_gather_scatter_req_0 : boolean;
  signal ptr_deref_2979_gather_scatter_ack_0 : boolean;
  signal type_cast_2983_inst_req_0 : boolean;
  signal type_cast_2983_inst_ack_0 : boolean;
  signal array_obj_ref_2990_base_resize_req_0 : boolean;
  signal array_obj_ref_2990_base_resize_ack_0 : boolean;
  signal array_obj_ref_2990_root_address_inst_req_0 : boolean;
  signal array_obj_ref_2990_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_2990_root_address_inst_req_1 : boolean;
  signal array_obj_ref_2990_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_2990_final_reg_req_0 : boolean;
  signal array_obj_ref_2990_final_reg_ack_0 : boolean;
  signal ptr_deref_2994_base_resize_req_0 : boolean;
  signal ptr_deref_2994_base_resize_ack_0 : boolean;
  signal ptr_deref_2994_root_address_inst_req_0 : boolean;
  signal ptr_deref_2994_root_address_inst_ack_0 : boolean;
  signal ptr_deref_2994_addr_0_req_0 : boolean;
  signal ptr_deref_2994_addr_0_ack_0 : boolean;
  signal ptr_deref_2994_addr_0_req_1 : boolean;
  signal ptr_deref_2994_addr_0_ack_1 : boolean;
  signal ptr_deref_2994_addr_1_req_0 : boolean;
  signal ptr_deref_2994_addr_1_ack_0 : boolean;
  signal ptr_deref_2994_addr_1_req_1 : boolean;
  signal ptr_deref_2994_addr_1_ack_1 : boolean;
  signal ptr_deref_2994_addr_2_req_0 : boolean;
  signal ptr_deref_2994_addr_2_ack_0 : boolean;
  signal ptr_deref_2994_addr_2_req_1 : boolean;
  signal ptr_deref_2994_addr_2_ack_1 : boolean;
  signal ptr_deref_2994_addr_3_req_0 : boolean;
  signal ptr_deref_2994_addr_3_ack_0 : boolean;
  signal ptr_deref_2994_addr_3_req_1 : boolean;
  signal ptr_deref_2994_addr_3_ack_1 : boolean;
  signal ptr_deref_2994_load_0_req_0 : boolean;
  signal ptr_deref_2994_load_0_ack_0 : boolean;
  signal ptr_deref_2994_load_1_req_0 : boolean;
  signal ptr_deref_2994_load_1_ack_0 : boolean;
  signal ptr_deref_2994_load_2_req_0 : boolean;
  signal ptr_deref_2994_load_2_ack_0 : boolean;
  signal ptr_deref_2994_load_3_req_0 : boolean;
  signal ptr_deref_2994_load_3_ack_0 : boolean;
  signal ptr_deref_2994_load_0_req_1 : boolean;
  signal ptr_deref_2994_load_0_ack_1 : boolean;
  signal ptr_deref_2994_load_1_req_1 : boolean;
  signal ptr_deref_2994_load_1_ack_1 : boolean;
  signal ptr_deref_2994_load_2_req_1 : boolean;
  signal ptr_deref_2994_load_2_ack_1 : boolean;
  signal ptr_deref_2994_load_3_req_1 : boolean;
  signal ptr_deref_2994_load_3_ack_1 : boolean;
  signal ptr_deref_2994_gather_scatter_req_0 : boolean;
  signal ptr_deref_2994_gather_scatter_ack_0 : boolean;
  signal type_cast_2998_inst_req_0 : boolean;
  signal type_cast_2998_inst_ack_0 : boolean;
  signal binary_3003_inst_req_0 : boolean;
  signal binary_3003_inst_ack_0 : boolean;
  signal binary_3003_inst_req_1 : boolean;
  signal binary_3003_inst_ack_1 : boolean;
  signal type_cast_3007_inst_req_0 : boolean;
  signal type_cast_3007_inst_ack_0 : boolean;
  signal binary_3013_inst_req_0 : boolean;
  signal binary_3013_inst_ack_0 : boolean;
  signal binary_3013_inst_req_1 : boolean;
  signal binary_3013_inst_ack_1 : boolean;
  signal type_cast_3017_inst_req_0 : boolean;
  signal type_cast_3017_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  ahir_glue_to3_CP_14633: Block -- control-path 
    signal cp_elements: BooleanArray(302 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(302);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(302), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(23);
    crr_14724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_2945_call_req_0); -- 
    cp_elements(2) <= cp_elements(199);
    crr_15249_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_3050_call_req_0); -- 
    cp_elements(3) <= cp_elements(295);
    pipe_wreq_15547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_3070_inst_req_0); -- 
    cp_elements(4) <= cp_elements(0);
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => type_cast_2926_inst_req_0); -- 
    cp_elements(6) <= cp_elements(4);
    cp_elements(7) <= cp_elements(4);
    req_14674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => simple_obj_ref_2925_inst_req_0); -- 
    ack_14675_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_2925_inst_ack_0, ack => cp_elements(8)); -- 
    ack_14680_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2926_inst_ack_0, ack => cp_elements(9)); -- 
    cp_elements(10) <= cp_elements(9);
    cpelement_group_11 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(13));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(11),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14692_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => type_cast_2930_inst_req_0); -- 
    cp_elements(12) <= cp_elements(10);
    cp_elements(13) <= cp_elements(10);
    ack_14693_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2930_inst_ack_0, ack => cp_elements(14)); -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => binary_2936_inst_req_0); -- 
    cp_elements(16) <= cp_elements(10);
    cp_elements(17) <= cp_elements(10);
    ra_14703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2936_inst_ack_0, ack => cp_elements(18)); -- 
    cr_14704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_2936_inst_req_1); -- 
    ca_14705_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2936_inst_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(21));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14714_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_2940_inst_req_0); -- 
    cp_elements(21) <= cp_elements(10);
    ack_14715_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2940_inst_ack_0, ack => cp_elements(22)); -- 
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_14725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2945_call_ack_0, ack => cp_elements(24)); -- 
    ccr_14729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => call_stmt_2945_call_req_1); -- 
    cca_14730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2945_call_ack_1, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(25);
    cp_elements(27) <= cp_elements(26);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(29) & cp_elements(39));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_14776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_2947_gather_scatter_req_0); -- 
    cp_elements(29) <= cp_elements(26);
    cp_elements(30) <= cp_elements(29);
    base_resize_req_14749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => ptr_deref_2947_base_resize_req_0); -- 
    base_resize_ack_14750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_base_resize_ack_0, ack => cp_elements(31)); -- 
    sum_rename_req_14754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_2947_root_address_inst_req_0); -- 
    cp_elements(32) <= ptr_deref_2947_root_address_inst_ack_0;
    cp_elements(33) <= cp_elements(32);
    rr_14762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => ptr_deref_2947_addr_0_req_0); -- 
    ra_14763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_addr_0_ack_0, ack => cp_elements(34)); -- 
    cr_14764_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => ptr_deref_2947_addr_0_req_1); -- 
    ca_14765_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_addr_0_ack_1, ack => cp_elements(35)); -- 
    cp_elements(36) <= cp_elements(32);
    rr_14769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_2947_addr_1_req_0); -- 
    ra_14770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_addr_1_ack_0, ack => cp_elements(37)); -- 
    cr_14771_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_2947_addr_1_req_1); -- 
    ca_14772_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_addr_1_ack_1, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(35) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= ptr_deref_2947_gather_scatter_ack_0;
    cp_elements(41) <= cp_elements(40);
    rr_14784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_2947_store_0_req_0); -- 
    ra_14785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_store_0_ack_0, ack => cp_elements(42)); -- 
    cp_elements(43) <= cp_elements(40);
    rr_14789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_2947_store_1_req_0); -- 
    ra_14790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_store_1_ack_0, ack => cp_elements(44)); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(42) & cp_elements(44));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(46) <= cp_elements(45);
    cp_elements(47) <= cp_elements(46);
    cr_14800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => ptr_deref_2947_store_0_req_1); -- 
    ca_14801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_store_0_ack_1, ack => cp_elements(48)); -- 
    cp_elements(49) <= cp_elements(46);
    cr_14805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => ptr_deref_2947_store_1_req_1); -- 
    ca_14806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2947_store_1_ack_1, ack => cp_elements(50)); -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(48) & cp_elements(50));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14815_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_2954_inst_req_0); -- 
    cp_elements(53) <= cp_elements(26);
    cp_elements(54) <= cp_elements(26);
    ra_14816_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2954_inst_ack_0, ack => cp_elements(55)); -- 
    cr_14817_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => binary_2954_inst_req_1); -- 
    ca_14818_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2954_inst_ack_1, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(56) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14827_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => type_cast_2958_inst_req_0); -- 
    cp_elements(58) <= cp_elements(26);
    ack_14828_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2958_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(62));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_14837_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => binary_2964_inst_req_0); -- 
    cp_elements(61) <= cp_elements(26);
    cp_elements(62) <= cp_elements(26);
    ra_14838_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2964_inst_ack_0, ack => cp_elements(63)); -- 
    cr_14839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => binary_2964_inst_req_1); -- 
    ca_14840_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_2964_inst_ack_1, ack => cp_elements(64)); -- 
    cpelement_group_65 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(64) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(65),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14849_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_2968_inst_req_0); -- 
    cp_elements(66) <= cp_elements(26);
    ack_14850_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2968_inst_ack_0, ack => cp_elements(67)); -- 
    cp_elements(68) <= cp_elements(26);
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(68) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_14874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => array_obj_ref_2975_final_reg_req_0); -- 
    cp_elements(70) <= cp_elements(26);
    base_resize_req_14861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => array_obj_ref_2975_base_resize_req_0); -- 
    base_resize_ack_14862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2975_base_resize_ack_0, ack => cp_elements(71)); -- 
    plus_base_rr_14867_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_2975_root_address_inst_req_0); -- 
    plus_base_ra_14868_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2975_root_address_inst_ack_0, ack => cp_elements(72)); -- 
    plus_base_cr_14869_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_2975_root_address_inst_req_1); -- 
    plus_base_ca_14870_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2975_root_address_inst_ack_1, ack => cp_elements(73)); -- 
    cp_elements(74) <= array_obj_ref_2975_final_reg_ack_0;
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(74) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(76) <= cp_elements(74);
    base_resize_req_14888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_2979_base_resize_req_0); -- 
    base_resize_ack_14889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_14893_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_2979_root_address_inst_req_0); -- 
    cp_elements(78) <= ptr_deref_2979_root_address_inst_ack_0;
    cp_elements(79) <= cp_elements(78);
    rr_14901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_2979_addr_0_req_0); -- 
    ra_14902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_0_ack_0, ack => cp_elements(80)); -- 
    cr_14903_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_2979_addr_0_req_1); -- 
    ca_14904_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_0_ack_1, ack => cp_elements(81)); -- 
    cp_elements(82) <= cp_elements(78);
    rr_14908_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_2979_addr_1_req_0); -- 
    ra_14909_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_1_ack_0, ack => cp_elements(83)); -- 
    cr_14910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_2979_addr_1_req_1); -- 
    ca_14911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_1_ack_1, ack => cp_elements(84)); -- 
    cp_elements(85) <= cp_elements(78);
    rr_14915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_2979_addr_2_req_0); -- 
    ra_14916_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_2_ack_0, ack => cp_elements(86)); -- 
    cr_14917_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_2979_addr_2_req_1); -- 
    ca_14918_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_2_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= cp_elements(78);
    rr_14922_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => ptr_deref_2979_addr_3_req_0); -- 
    ra_14923_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_3_ack_0, ack => cp_elements(89)); -- 
    cr_14924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => ptr_deref_2979_addr_3_req_1); -- 
    ca_14925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_addr_3_ack_1, ack => cp_elements(90)); -- 
    cpelement_group_91 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(84) & cp_elements(87) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(91),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(92) <= cp_elements(75);
    rr_14935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_2979_load_0_req_0); -- 
    ra_14936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_0_ack_0, ack => cp_elements(93)); -- 
    cp_elements(94) <= cp_elements(75);
    rr_14940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_2979_load_1_req_0); -- 
    ra_14941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_1_ack_0, ack => cp_elements(95)); -- 
    cp_elements(96) <= cp_elements(75);
    rr_14945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_2979_load_2_req_0); -- 
    ra_14946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_2_ack_0, ack => cp_elements(97)); -- 
    cp_elements(98) <= cp_elements(75);
    rr_14950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_2979_load_3_req_0); -- 
    ra_14951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_3_ack_0, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(93) & cp_elements(95) & cp_elements(97) & cp_elements(99));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(101) <= cp_elements(100);
    cr_14961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => ptr_deref_2979_load_0_req_1); -- 
    ca_14962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_0_ack_1, ack => cp_elements(102)); -- 
    cp_elements(103) <= cp_elements(100);
    cr_14966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => ptr_deref_2979_load_1_req_1); -- 
    ca_14967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_1_ack_1, ack => cp_elements(104)); -- 
    cp_elements(105) <= cp_elements(100);
    cr_14971_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => ptr_deref_2979_load_2_req_1); -- 
    ca_14972_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_2_ack_1, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(100);
    cr_14976_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_2979_load_3_req_1); -- 
    ca_14977_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_load_3_ack_1, ack => cp_elements(108)); -- 
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(104) & cp_elements(106) & cp_elements(108));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_14978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_2979_gather_scatter_req_0); -- 
    merge_ack_14979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2979_gather_scatter_ack_0, ack => cp_elements(110)); -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_14988_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => type_cast_2983_inst_req_0); -- 
    cp_elements(112) <= cp_elements(26);
    ack_14989_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2983_inst_ack_0, ack => cp_elements(113)); -- 
    cp_elements(114) <= cp_elements(26);
    cpelement_group_115 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(114) & cp_elements(119));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(115),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => array_obj_ref_2990_final_reg_req_0); -- 
    cp_elements(116) <= cp_elements(26);
    base_resize_req_15000_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => array_obj_ref_2990_base_resize_req_0); -- 
    base_resize_ack_15001_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2990_base_resize_ack_0, ack => cp_elements(117)); -- 
    plus_base_rr_15006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_2990_root_address_inst_req_0); -- 
    plus_base_ra_15007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2990_root_address_inst_ack_0, ack => cp_elements(118)); -- 
    plus_base_cr_15008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_2990_root_address_inst_req_1); -- 
    plus_base_ca_15009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2990_root_address_inst_ack_1, ack => cp_elements(119)); -- 
    cp_elements(120) <= array_obj_ref_2990_final_reg_ack_0;
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(120) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(120);
    base_resize_req_15027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_2994_base_resize_req_0); -- 
    base_resize_ack_15028_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_base_resize_ack_0, ack => cp_elements(123)); -- 
    sum_rename_req_15032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => ptr_deref_2994_root_address_inst_req_0); -- 
    cp_elements(124) <= ptr_deref_2994_root_address_inst_ack_0;
    cp_elements(125) <= cp_elements(124);
    rr_15040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(125), ack => ptr_deref_2994_addr_0_req_0); -- 
    ra_15041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_0_ack_0, ack => cp_elements(126)); -- 
    cr_15042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => ptr_deref_2994_addr_0_req_1); -- 
    ca_15043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_0_ack_1, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(124);
    rr_15047_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => ptr_deref_2994_addr_1_req_0); -- 
    ra_15048_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_1_ack_0, ack => cp_elements(129)); -- 
    cr_15049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_2994_addr_1_req_1); -- 
    ca_15050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_1_ack_1, ack => cp_elements(130)); -- 
    cp_elements(131) <= cp_elements(124);
    rr_15054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_2994_addr_2_req_0); -- 
    ra_15055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_2_ack_0, ack => cp_elements(132)); -- 
    cr_15056_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => ptr_deref_2994_addr_2_req_1); -- 
    ca_15057_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_2_ack_1, ack => cp_elements(133)); -- 
    cp_elements(134) <= cp_elements(124);
    rr_15061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => ptr_deref_2994_addr_3_req_0); -- 
    ra_15062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_3_ack_0, ack => cp_elements(135)); -- 
    cr_15063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(135), ack => ptr_deref_2994_addr_3_req_1); -- 
    ca_15064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_addr_3_ack_1, ack => cp_elements(136)); -- 
    cpelement_group_137 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(130) & cp_elements(133) & cp_elements(136));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(137),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(138) <= cp_elements(121);
    rr_15074_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => ptr_deref_2994_load_0_req_0); -- 
    ra_15075_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_0_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(121);
    rr_15079_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => ptr_deref_2994_load_1_req_0); -- 
    ra_15080_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_1_ack_0, ack => cp_elements(141)); -- 
    cp_elements(142) <= cp_elements(121);
    rr_15084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_2994_load_2_req_0); -- 
    ra_15085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_2_ack_0, ack => cp_elements(143)); -- 
    cp_elements(144) <= cp_elements(121);
    rr_15089_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => ptr_deref_2994_load_3_req_0); -- 
    ra_15090_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_3_ack_0, ack => cp_elements(145)); -- 
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(139) & cp_elements(141) & cp_elements(143) & cp_elements(145));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(147) <= cp_elements(146);
    cr_15100_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(147), ack => ptr_deref_2994_load_0_req_1); -- 
    ca_15101_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_0_ack_1, ack => cp_elements(148)); -- 
    cp_elements(149) <= cp_elements(146);
    cr_15105_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_2994_load_1_req_1); -- 
    ca_15106_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_1_ack_1, ack => cp_elements(150)); -- 
    cp_elements(151) <= cp_elements(146);
    cr_15110_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(151), ack => ptr_deref_2994_load_2_req_1); -- 
    ca_15111_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_2_ack_1, ack => cp_elements(152)); -- 
    cp_elements(153) <= cp_elements(146);
    cr_15115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => ptr_deref_2994_load_3_req_1); -- 
    ca_15116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_load_3_ack_1, ack => cp_elements(154)); -- 
    cpelement_group_155 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(148) & cp_elements(150) & cp_elements(152) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_15117_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => ptr_deref_2994_gather_scatter_req_0); -- 
    merge_ack_15118_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_2994_gather_scatter_ack_0, ack => cp_elements(156)); -- 
    cpelement_group_157 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(156) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(157),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => type_cast_2998_inst_req_0); -- 
    cp_elements(158) <= cp_elements(26);
    ack_15128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_2998_inst_ack_0, ack => cp_elements(159)); -- 
    cpelement_group_160 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(159) & cp_elements(161));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(160),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_3003_inst_req_0); -- 
    cp_elements(161) <= cp_elements(26);
    ra_15139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3003_inst_ack_0, ack => cp_elements(162)); -- 
    cr_15140_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => binary_3003_inst_req_1); -- 
    cp_elements(163) <= binary_3003_inst_ack_1;
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15150_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(164), ack => type_cast_3007_inst_req_0); -- 
    cp_elements(165) <= cp_elements(26);
    cp_elements(166) <= cp_elements(163);
    ack_15151_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3007_inst_ack_0, ack => cp_elements(167)); -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(170));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15160_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_3013_inst_req_0); -- 
    cp_elements(169) <= cp_elements(26);
    cp_elements(170) <= cp_elements(163);
    ra_15161_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3013_inst_ack_0, ack => cp_elements(171)); -- 
    cr_15162_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_3013_inst_req_1); -- 
    ca_15163_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3013_inst_ack_1, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_3017_inst_req_0); -- 
    cp_elements(174) <= cp_elements(26);
    ack_15173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3017_inst_ack_0, ack => cp_elements(175)); -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(175) & cp_elements(177));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15182_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(176), ack => binary_3023_inst_req_0); -- 
    cp_elements(177) <= cp_elements(26);
    ra_15183_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3023_inst_ack_0, ack => cp_elements(178)); -- 
    cr_15184_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(178), ack => binary_3023_inst_req_1); -- 
    ca_15185_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3023_inst_ack_1, ack => cp_elements(179)); -- 
    cpelement_group_180 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(181) & cp_elements(182));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(180),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15194_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_3029_inst_req_0); -- 
    cp_elements(181) <= cp_elements(26);
    cp_elements(182) <= cp_elements(163);
    ra_15195_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3029_inst_ack_0, ack => cp_elements(183)); -- 
    cr_15196_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_3029_inst_req_1); -- 
    ca_15197_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3029_inst_ack_1, ack => cp_elements(184)); -- 
    cpelement_group_185 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(185),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_3037_inst_req_0); -- 
    cp_elements(186) <= cp_elements(26);
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(184) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_3033_inst_req_0); -- 
    cp_elements(188) <= cp_elements(26);
    ack_15209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3033_inst_ack_0, ack => cp_elements(189)); -- 
    ra_15214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3037_inst_ack_0, ack => cp_elements(190)); -- 
    cr_15215_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => binary_3037_inst_req_1); -- 
    ca_15216_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3037_inst_ack_1, ack => cp_elements(191)); -- 
    cpelement_group_192 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(191) & cp_elements(193));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(192),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(192), ack => type_cast_3041_inst_req_0); -- 
    cp_elements(193) <= cp_elements(26);
    ack_15226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3041_inst_ack_0, ack => cp_elements(194)); -- 
    cpelement_group_195 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(179) & cp_elements(194) & cp_elements(196));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(195),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => binary_3046_inst_req_0); -- 
    cp_elements(196) <= cp_elements(26);
    ra_15237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3046_inst_ack_0, ack => cp_elements(197)); -- 
    cr_15238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => binary_3046_inst_req_1); -- 
    ca_15239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3046_inst_ack_1, ack => cp_elements(198)); -- 
    cpelement_group_199 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67) & cp_elements(167) & cp_elements(198));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(199),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cra_15250_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3050_call_ack_0, ack => cp_elements(200)); -- 
    ccr_15254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => call_stmt_3050_call_req_1); -- 
    cca_15255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3050_call_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(201);
    cp_elements(203) <= cp_elements(202);
    cpelement_group_204 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(203) & cp_elements(205) & cp_elements(215));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(204),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_15301_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => ptr_deref_3052_gather_scatter_req_0); -- 
    cp_elements(205) <= cp_elements(202);
    cp_elements(206) <= cp_elements(205);
    base_resize_req_15274_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_3052_base_resize_req_0); -- 
    base_resize_ack_15275_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_base_resize_ack_0, ack => cp_elements(207)); -- 
    sum_rename_req_15279_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => ptr_deref_3052_root_address_inst_req_0); -- 
    cp_elements(208) <= ptr_deref_3052_root_address_inst_ack_0;
    cp_elements(209) <= cp_elements(208);
    rr_15287_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_3052_addr_0_req_0); -- 
    ra_15288_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_addr_0_ack_0, ack => cp_elements(210)); -- 
    cr_15289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(210), ack => ptr_deref_3052_addr_0_req_1); -- 
    ca_15290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_addr_0_ack_1, ack => cp_elements(211)); -- 
    cp_elements(212) <= cp_elements(208);
    rr_15294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_3052_addr_1_req_0); -- 
    ra_15295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_addr_1_ack_0, ack => cp_elements(213)); -- 
    cr_15296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(213), ack => ptr_deref_3052_addr_1_req_1); -- 
    ca_15297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_addr_1_ack_1, ack => cp_elements(214)); -- 
    cpelement_group_215 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(211) & cp_elements(214));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(215),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(216) <= ptr_deref_3052_gather_scatter_ack_0;
    cp_elements(217) <= cp_elements(216);
    rr_15309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_3052_store_0_req_0); -- 
    ra_15310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_store_0_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(216);
    rr_15314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_3052_store_1_req_0); -- 
    ra_15315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_store_1_ack_0, ack => cp_elements(220)); -- 
    cpelement_group_221 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(218) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(221),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(222) <= cp_elements(221);
    cr_15325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(222), ack => ptr_deref_3052_store_0_req_1); -- 
    ca_15326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_store_0_ack_1, ack => cp_elements(223)); -- 
    cp_elements(224) <= cp_elements(221);
    cr_15330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(224), ack => ptr_deref_3052_store_1_req_1); -- 
    ca_15331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3052_store_1_ack_1, ack => cp_elements(225)); -- 
    cpelement_group_226 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(223) & cp_elements(225));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(226),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    crr_15341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(226), ack => call_stmt_3057_call_req_0); -- 
    cra_15342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3057_call_ack_0, ack => cp_elements(227)); -- 
    ccr_15346_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => call_stmt_3057_call_req_1); -- 
    cca_15347_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3057_call_ack_1, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(228);
    cp_elements(230) <= cp_elements(229);
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(230) & cp_elements(232) & cp_elements(242));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_15393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(231), ack => ptr_deref_3059_gather_scatter_req_0); -- 
    cp_elements(232) <= cp_elements(229);
    cp_elements(233) <= cp_elements(232);
    base_resize_req_15366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => ptr_deref_3059_base_resize_req_0); -- 
    base_resize_ack_15367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_base_resize_ack_0, ack => cp_elements(234)); -- 
    sum_rename_req_15371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_3059_root_address_inst_req_0); -- 
    cp_elements(235) <= ptr_deref_3059_root_address_inst_ack_0;
    cp_elements(236) <= cp_elements(235);
    rr_15379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_3059_addr_0_req_0); -- 
    ra_15380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_addr_0_ack_0, ack => cp_elements(237)); -- 
    cr_15381_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(237), ack => ptr_deref_3059_addr_0_req_1); -- 
    ca_15382_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_addr_0_ack_1, ack => cp_elements(238)); -- 
    cp_elements(239) <= cp_elements(235);
    rr_15386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(239), ack => ptr_deref_3059_addr_1_req_0); -- 
    ra_15387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_addr_1_ack_0, ack => cp_elements(240)); -- 
    cr_15388_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_3059_addr_1_req_1); -- 
    ca_15389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_addr_1_ack_1, ack => cp_elements(241)); -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(238) & cp_elements(241));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(243) <= ptr_deref_3059_gather_scatter_ack_0;
    cp_elements(244) <= cp_elements(243);
    rr_15401_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_3059_store_0_req_0); -- 
    ra_15402_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_store_0_ack_0, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(243);
    rr_15406_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_3059_store_1_req_0); -- 
    ra_15407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_store_1_ack_0, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(249) <= cp_elements(248);
    cp_elements(250) <= cp_elements(249);
    cr_15417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => ptr_deref_3059_store_0_req_1); -- 
    ca_15418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_store_0_ack_1, ack => cp_elements(251)); -- 
    cp_elements(252) <= cp_elements(249);
    cr_15422_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => ptr_deref_3059_store_1_req_1); -- 
    ca_15423_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3059_store_1_ack_1, ack => cp_elements(253)); -- 
    cpelement_group_254 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(251) & cp_elements(253));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(254),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cpelement_group_255 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(248) & cp_elements(256) & cp_elements(272));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(255),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(256) <= cp_elements(229);
    cp_elements(257) <= cp_elements(256);
    base_resize_req_15436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(257), ack => ptr_deref_3064_base_resize_req_0); -- 
    base_resize_ack_15437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_base_resize_ack_0, ack => cp_elements(258)); -- 
    sum_rename_req_15441_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(258), ack => ptr_deref_3064_root_address_inst_req_0); -- 
    cp_elements(259) <= ptr_deref_3064_root_address_inst_ack_0;
    cp_elements(260) <= cp_elements(259);
    rr_15449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => ptr_deref_3064_addr_0_req_0); -- 
    ra_15450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_0_ack_0, ack => cp_elements(261)); -- 
    cr_15451_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(261), ack => ptr_deref_3064_addr_0_req_1); -- 
    ca_15452_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_0_ack_1, ack => cp_elements(262)); -- 
    cp_elements(263) <= cp_elements(259);
    rr_15456_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => ptr_deref_3064_addr_1_req_0); -- 
    ra_15457_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_1_ack_0, ack => cp_elements(264)); -- 
    cr_15458_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(264), ack => ptr_deref_3064_addr_1_req_1); -- 
    ca_15459_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_1_ack_1, ack => cp_elements(265)); -- 
    cp_elements(266) <= cp_elements(259);
    rr_15463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_3064_addr_2_req_0); -- 
    ra_15464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_2_ack_0, ack => cp_elements(267)); -- 
    cr_15465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(267), ack => ptr_deref_3064_addr_2_req_1); -- 
    ca_15466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_2_ack_1, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(259);
    rr_15470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_3064_addr_3_req_0); -- 
    ra_15471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_3_ack_0, ack => cp_elements(270)); -- 
    cr_15472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => ptr_deref_3064_addr_3_req_1); -- 
    ca_15473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_addr_3_ack_1, ack => cp_elements(271)); -- 
    cpelement_group_272 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(262) & cp_elements(265) & cp_elements(268) & cp_elements(271));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(272),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(273) <= cp_elements(255);
    rr_15483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => ptr_deref_3064_load_0_req_0); -- 
    ra_15484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_0_ack_0, ack => cp_elements(274)); -- 
    cp_elements(275) <= cp_elements(255);
    rr_15488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_3064_load_1_req_0); -- 
    ra_15489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_1_ack_0, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(255);
    rr_15493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_3064_load_2_req_0); -- 
    ra_15494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_2_ack_0, ack => cp_elements(278)); -- 
    cp_elements(279) <= cp_elements(255);
    rr_15498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(279), ack => ptr_deref_3064_load_3_req_0); -- 
    ra_15499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_3_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(276) & cp_elements(278) & cp_elements(280));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(282) <= cp_elements(281);
    cr_15509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(282), ack => ptr_deref_3064_load_0_req_1); -- 
    ca_15510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_0_ack_1, ack => cp_elements(283)); -- 
    cp_elements(284) <= cp_elements(281);
    cr_15514_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_3064_load_1_req_1); -- 
    ca_15515_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_1_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(281);
    cr_15519_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_3064_load_2_req_1); -- 
    ca_15520_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_2_ack_1, ack => cp_elements(287)); -- 
    cp_elements(288) <= cp_elements(281);
    cr_15524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => ptr_deref_3064_load_3_req_1); -- 
    ca_15525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_load_3_ack_1, ack => cp_elements(289)); -- 
    cpelement_group_290 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(283) & cp_elements(285) & cp_elements(287) & cp_elements(289));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(290),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_15526_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_3064_gather_scatter_req_0); -- 
    merge_ack_15527_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3064_gather_scatter_ack_0, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(291) & cp_elements(293));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => type_cast_3068_inst_req_0); -- 
    cp_elements(293) <= cp_elements(229);
    ack_15537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3068_inst_ack_0, ack => cp_elements(294)); -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(254) & cp_elements(294));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_15548_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3070_inst_ack_0, ack => cp_elements(296)); -- 
    cp_elements(297) <= cp_elements(296);
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(299) & cp_elements(300));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15560_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => type_cast_3076_inst_req_0); -- 
    cp_elements(299) <= cp_elements(297);
    cp_elements(300) <= cp_elements(297);
    ack_15561_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3076_inst_ack_0, ack => cp_elements(301)); -- 
    pipe_wreq_15566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => simple_obj_ref_3074_inst_req_0); -- 
    pipe_wack_15567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3074_inst_ack_0, ack => cp_elements(302)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_2975_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2975_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2975_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2990_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_2990_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_2990_root_address : std_logic_vector(15 downto 0);
    signal notx_xx_xi_3038 : std_logic_vector(0 downto 0);
    signal ptr_deref_2947_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2947_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2947_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2947_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2979_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2979_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2979_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2979_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2979_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_2994_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_2994_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_2994_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_2994_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_2994_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3052_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3052_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3052_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3059_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3059_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_wire : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3059_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3064_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3064_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_3064_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_3064_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3064_word_offset_3 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_2925_wire : std_logic_vector(31 downto 0);
    signal tmp10_2980 : std_logic_vector(31 downto 0);
    signal tmp11_2984 : std_logic_vector(31 downto 0);
    signal tmp12_2991 : std_logic_vector(31 downto 0);
    signal tmp13_2995 : std_logic_vector(31 downto 0);
    signal tmp14_2999 : std_logic_vector(31 downto 0);
    signal tmp15_3004 : std_logic_vector(31 downto 0);
    signal tmp16_3008 : std_logic_vector(15 downto 0);
    signal tmp17_3014 : std_logic_vector(31 downto 0);
    signal tmp18_3024 : std_logic_vector(15 downto 0);
    signal tmp19_3030 : std_logic_vector(31 downto 0);
    signal tmp1_2931 : std_logic_vector(31 downto 0);
    signal tmp20_3042 : std_logic_vector(15 downto 0);
    signal tmp21_3047 : std_logic_vector(15 downto 0);
    signal tmp22_3050 : std_logic_vector(15 downto 0);
    signal tmp23_3057 : std_logic_vector(15 downto 0);
    signal tmp24_3065 : std_logic_vector(31 downto 0);
    signal tmp25_3069 : std_logic_vector(31 downto 0);
    signal tmp2_2937 : std_logic_vector(31 downto 0);
    signal tmp3_2941 : std_logic_vector(31 downto 0);
    signal tmp4_2945 : std_logic_vector(15 downto 0);
    signal tmp5_2955 : std_logic_vector(31 downto 0);
    signal tmp6_2959 : std_logic_vector(31 downto 0);
    signal tmp7_2965 : std_logic_vector(31 downto 0);
    signal tmp8_2969 : std_logic_vector(31 downto 0);
    signal tmp9_2976 : std_logic_vector(31 downto 0);
    signal tmp_2927 : std_logic_vector(31 downto 0);
    signal type_cast_2935_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2943_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_2953_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2963_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3012_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3022_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3028_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3033_wire : std_logic_vector(31 downto 0);
    signal type_cast_3036_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3072_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3076_wire : std_logic_vector(31 downto 0);
    signal xx_xtrx_xi_3018 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_2975_final_offset <= "0000000000010000";
    array_obj_ref_2990_final_offset <= "0000000000001100";
    ptr_deref_2947_word_offset_0 <= "0000000000000000";
    ptr_deref_2947_word_offset_1 <= "0000000000000001";
    ptr_deref_2979_word_offset_0 <= "0000000000000000";
    ptr_deref_2979_word_offset_1 <= "0000000000000001";
    ptr_deref_2979_word_offset_2 <= "0000000000000010";
    ptr_deref_2979_word_offset_3 <= "0000000000000011";
    ptr_deref_2994_word_offset_0 <= "0000000000000000";
    ptr_deref_2994_word_offset_1 <= "0000000000000001";
    ptr_deref_2994_word_offset_2 <= "0000000000000010";
    ptr_deref_2994_word_offset_3 <= "0000000000000011";
    ptr_deref_3052_word_offset_0 <= "0000000000000000";
    ptr_deref_3052_word_offset_1 <= "0000000000000001";
    ptr_deref_3059_word_offset_0 <= "0000000000000000";
    ptr_deref_3059_word_offset_1 <= "0000000000000001";
    ptr_deref_3064_word_offset_0 <= "0000000000000000";
    ptr_deref_3064_word_offset_1 <= "0000000000000001";
    ptr_deref_3064_word_offset_2 <= "0000000000000010";
    ptr_deref_3064_word_offset_3 <= "0000000000000011";
    type_cast_2935_wire_constant <= "11111111111111111111100000000000";
    type_cast_2943_wire_constant <= "0000000000001000";
    type_cast_2953_wire_constant <= "00000000000000000000000000000110";
    type_cast_2963_wire_constant <= "00000000000000000000000000000010";
    type_cast_3012_wire_constant <= "00000000000000000000000000000011";
    type_cast_3022_wire_constant <= "0001111111111111";
    type_cast_3028_wire_constant <= "00000000000000000000000000000111";
    type_cast_3036_wire_constant <= "00000000000000000000000000000000";
    type_cast_3072_wire_constant <= "00000000000000000000000000000100";
    array_obj_ref_2975_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2931, dout => array_obj_ref_2975_resized_base_address, req => array_obj_ref_2975_base_resize_req_0, ack => array_obj_ref_2975_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2975_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2975_root_address, dout => tmp9_2976, req => array_obj_ref_2975_final_reg_req_0, ack => array_obj_ref_2975_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2990_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp1_2931, dout => array_obj_ref_2990_resized_base_address, req => array_obj_ref_2990_base_resize_req_0, ack => array_obj_ref_2990_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_2990_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_2990_root_address, dout => tmp12_2991, req => array_obj_ref_2990_final_reg_req_0, ack => array_obj_ref_2990_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2947_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp3_2941, dout => ptr_deref_2947_resized_base_address, req => ptr_deref_2947_base_resize_req_0, ack => ptr_deref_2947_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2979_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp9_2976, dout => ptr_deref_2979_resized_base_address, req => ptr_deref_2979_base_resize_req_0, ack => ptr_deref_2979_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2994_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2991, dout => ptr_deref_2994_resized_base_address, req => ptr_deref_2994_base_resize_req_0, ack => ptr_deref_2994_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3052_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp6_2959, dout => ptr_deref_3052_resized_base_address, req => ptr_deref_3052_base_resize_req_0, ack => ptr_deref_3052_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3059_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp8_2969, dout => ptr_deref_3059_resized_base_address, req => ptr_deref_3059_base_resize_req_0, ack => ptr_deref_3059_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3064_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => tmp12_2991, dout => ptr_deref_3064_resized_base_address, req => ptr_deref_3064_base_resize_req_0, ack => ptr_deref_3064_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_2926_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => simple_obj_ref_2925_wire, dout => tmp_2927, req => type_cast_2926_inst_req_0, ack => type_cast_2926_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2930_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp_2927, dout => tmp1_2931, req => type_cast_2930_inst_req_0, ack => type_cast_2930_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2940_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp2_2937, dout => tmp3_2941, req => type_cast_2940_inst_req_0, ack => type_cast_2940_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2958_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp5_2955, dout => tmp6_2959, req => type_cast_2958_inst_req_0, ack => type_cast_2958_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2968_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp7_2965, dout => tmp8_2969, req => type_cast_2968_inst_req_0, ack => type_cast_2968_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2983_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp10_2980, dout => tmp11_2984, req => type_cast_2983_inst_req_0, ack => type_cast_2983_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_2998_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp13_2995, dout => tmp14_2999, req => type_cast_2998_inst_req_0, ack => type_cast_2998_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3007_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp15_3004, dout => tmp16_3008, req => type_cast_3007_inst_req_0, ack => type_cast_3007_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3017_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => tmp17_3014, dout => xx_xtrx_xi_3018, req => type_cast_3017_inst_req_0, ack => type_cast_3017_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3033_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp19_3030, dout => type_cast_3033_wire, req => type_cast_3033_inst_req_0, ack => type_cast_3033_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3041_inst: RegisterBase --
      generic map(in_data_width => 1,out_data_width => 16, flow_through => false ) 
      port map( din => notx_xx_xi_3038, dout => tmp20_3042, req => type_cast_3041_inst_req_0, ack => type_cast_3041_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3068_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => tmp24_3065, dout => tmp25_3069, req => type_cast_3068_inst_req_0, ack => type_cast_3068_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3076_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => tmp25_3069, dout => type_cast_3076_wire, req => type_cast_3076_inst_req_0, ack => type_cast_3076_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_2947_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2947_gather_scatter_ack_0 <= ptr_deref_2947_gather_scatter_req_0;
      aggregated_sig <= tmp4_2945;
      ptr_deref_2947_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_2947_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_2947_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2947_root_address_inst_ack_0 <= ptr_deref_2947_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2947_resized_base_address;
      ptr_deref_2947_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2979_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2979_gather_scatter_ack_0 <= ptr_deref_2979_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2979_data_3 & ptr_deref_2979_data_2 & ptr_deref_2979_data_1 & ptr_deref_2979_data_0;
      tmp10_2980 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2979_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2979_root_address_inst_ack_0 <= ptr_deref_2979_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2979_resized_base_address;
      ptr_deref_2979_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_2994_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_2994_gather_scatter_ack_0 <= ptr_deref_2994_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_2994_data_3 & ptr_deref_2994_data_2 & ptr_deref_2994_data_1 & ptr_deref_2994_data_0;
      tmp13_2995 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_2994_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_2994_root_address_inst_ack_0 <= ptr_deref_2994_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_2994_resized_base_address;
      ptr_deref_2994_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3052_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3052_gather_scatter_ack_0 <= ptr_deref_3052_gather_scatter_req_0;
      aggregated_sig <= tmp22_3050;
      ptr_deref_3052_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_3052_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_3052_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3052_root_address_inst_ack_0 <= ptr_deref_3052_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3052_resized_base_address;
      ptr_deref_3052_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3059_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3059_gather_scatter_ack_0 <= ptr_deref_3059_gather_scatter_req_0;
      aggregated_sig <= tmp23_3057;
      ptr_deref_3059_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_3059_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_3059_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3059_root_address_inst_ack_0 <= ptr_deref_3059_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3059_resized_base_address;
      ptr_deref_3059_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3064_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3064_gather_scatter_ack_0 <= ptr_deref_3064_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3064_data_3 & ptr_deref_3064_data_2 & ptr_deref_3064_data_1 & ptr_deref_3064_data_0;
      tmp24_3065 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3064_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3064_root_address_inst_ack_0 <= ptr_deref_3064_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3064_resized_base_address;
      ptr_deref_3064_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_2975_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2975_resized_base_address;
      array_obj_ref_2975_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000010000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2975_root_address_inst_req_0,
          ackL => array_obj_ref_2975_root_address_inst_ack_0,
          reqR => array_obj_ref_2975_root_address_inst_req_1,
          ackR => array_obj_ref_2975_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_2990_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_2990_resized_base_address;
      array_obj_ref_2990_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_2990_root_address_inst_req_0,
          ackL => array_obj_ref_2990_root_address_inst_ack_0,
          reqR => array_obj_ref_2990_root_address_inst_req_1,
          ackR => array_obj_ref_2990_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_2936_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp_2927;
      tmp2_2937 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2936_inst_req_0,
          ackL => binary_2936_inst_ack_0,
          reqR => binary_2936_inst_req_1,
          ackR => binary_2936_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_2954_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2937;
      tmp5_2955 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2954_inst_req_0,
          ackL => binary_2954_inst_ack_0,
          reqR => binary_2954_inst_req_1,
          ackR => binary_2954_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_2964_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_2937;
      tmp7_2965 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_2964_inst_req_0,
          ackL => binary_2964_inst_ack_0,
          reqR => binary_2964_inst_req_1,
          ackR => binary_2964_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_3003_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp11_2984 & tmp14_2999;
      tmp15_3004 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3003_inst_req_0,
          ackL => binary_3003_inst_ack_0,
          reqR => binary_3003_inst_req_1,
          ackR => binary_3003_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_3013_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_3004;
      tmp17_3014 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3013_inst_req_0,
          ackL => binary_3013_inst_ack_0,
          reqR => binary_3013_inst_req_1,
          ackR => binary_3013_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_3023_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= xx_xtrx_xi_3018;
      tmp18_3024 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0001111111111111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3023_inst_req_0,
          ackL => binary_3023_inst_ack_0,
          reqR => binary_3023_inst_req_1,
          ackR => binary_3023_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_3029_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp15_3004;
      tmp19_3030 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3029_inst_req_0,
          ackL => binary_3029_inst_ack_0,
          reqR => binary_3029_inst_req_1,
          ackR => binary_3029_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_3037_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3033_wire;
      notx_xx_xi_3038 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3037_inst_req_0,
          ackL => binary_3037_inst_ack_0,
          reqR => binary_3037_inst_req_1,
          ackR => binary_3037_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_3046_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp18_3024 & tmp20_3042;
      tmp21_3047 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3046_inst_req_0,
          ackL => binary_3046_inst_ack_0,
          reqR => binary_3046_inst_req_1,
          ackR => binary_3046_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_2947_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2947_root_address;
      ptr_deref_2947_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2947_addr_0_req_0,
          ackL => ptr_deref_2947_addr_0_ack_0,
          reqR => ptr_deref_2947_addr_0_req_1,
          ackR => ptr_deref_2947_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_2947_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2947_root_address;
      ptr_deref_2947_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2947_addr_1_req_0,
          ackL => ptr_deref_2947_addr_1_ack_0,
          reqR => ptr_deref_2947_addr_1_req_1,
          ackR => ptr_deref_2947_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_2979_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2979_root_address;
      ptr_deref_2979_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2979_addr_0_req_0,
          ackL => ptr_deref_2979_addr_0_ack_0,
          reqR => ptr_deref_2979_addr_0_req_1,
          ackR => ptr_deref_2979_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_2979_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2979_root_address;
      ptr_deref_2979_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2979_addr_1_req_0,
          ackL => ptr_deref_2979_addr_1_ack_0,
          reqR => ptr_deref_2979_addr_1_req_1,
          ackR => ptr_deref_2979_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_2979_addr_2 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2979_root_address;
      ptr_deref_2979_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2979_addr_2_req_0,
          ackL => ptr_deref_2979_addr_2_ack_0,
          reqR => ptr_deref_2979_addr_2_req_1,
          ackR => ptr_deref_2979_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_2979_addr_3 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2979_root_address;
      ptr_deref_2979_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2979_addr_3_req_0,
          ackL => ptr_deref_2979_addr_3_ack_0,
          reqR => ptr_deref_2979_addr_3_req_1,
          ackR => ptr_deref_2979_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_2994_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2994_root_address;
      ptr_deref_2994_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2994_addr_0_req_0,
          ackL => ptr_deref_2994_addr_0_ack_0,
          reqR => ptr_deref_2994_addr_0_req_1,
          ackR => ptr_deref_2994_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_2994_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2994_root_address;
      ptr_deref_2994_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2994_addr_1_req_0,
          ackL => ptr_deref_2994_addr_1_ack_0,
          reqR => ptr_deref_2994_addr_1_req_1,
          ackR => ptr_deref_2994_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : ptr_deref_2994_addr_2 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2994_root_address;
      ptr_deref_2994_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2994_addr_2_req_0,
          ackL => ptr_deref_2994_addr_2_ack_0,
          reqR => ptr_deref_2994_addr_2_req_1,
          ackR => ptr_deref_2994_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : ptr_deref_2994_addr_3 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_2994_root_address;
      ptr_deref_2994_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_2994_addr_3_req_0,
          ackL => ptr_deref_2994_addr_3_ack_0,
          reqR => ptr_deref_2994_addr_3_req_1,
          ackR => ptr_deref_2994_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_3052_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3052_root_address;
      ptr_deref_3052_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3052_addr_0_req_0,
          ackL => ptr_deref_3052_addr_0_ack_0,
          reqR => ptr_deref_3052_addr_0_req_1,
          ackR => ptr_deref_3052_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_3052_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3052_root_address;
      ptr_deref_3052_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3052_addr_1_req_0,
          ackL => ptr_deref_3052_addr_1_ack_0,
          reqR => ptr_deref_3052_addr_1_req_1,
          ackR => ptr_deref_3052_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_3059_addr_0 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3059_root_address;
      ptr_deref_3059_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3059_addr_0_req_0,
          ackL => ptr_deref_3059_addr_0_ack_0,
          reqR => ptr_deref_3059_addr_0_req_1,
          ackR => ptr_deref_3059_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_3059_addr_1 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3059_root_address;
      ptr_deref_3059_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3059_addr_1_req_0,
          ackL => ptr_deref_3059_addr_1_ack_0,
          reqR => ptr_deref_3059_addr_1_req_1,
          ackR => ptr_deref_3059_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_3064_addr_0 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3064_root_address;
      ptr_deref_3064_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3064_addr_0_req_0,
          ackL => ptr_deref_3064_addr_0_ack_0,
          reqR => ptr_deref_3064_addr_0_req_1,
          ackR => ptr_deref_3064_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_3064_addr_1 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3064_root_address;
      ptr_deref_3064_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3064_addr_1_req_0,
          ackL => ptr_deref_3064_addr_1_ack_0,
          reqR => ptr_deref_3064_addr_1_req_1,
          ackR => ptr_deref_3064_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_3064_addr_2 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3064_root_address;
      ptr_deref_3064_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3064_addr_2_req_0,
          ackL => ptr_deref_3064_addr_2_ack_0,
          reqR => ptr_deref_3064_addr_2_req_1,
          ackR => ptr_deref_3064_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_3064_addr_3 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3064_root_address;
      ptr_deref_3064_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3064_addr_3_req_0,
          ackL => ptr_deref_3064_addr_3_ack_0,
          reqR => ptr_deref_3064_addr_3_req_1,
          ackR => ptr_deref_3064_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared load operator group (0) : ptr_deref_2979_load_0 ptr_deref_2979_load_1 ptr_deref_2979_load_2 ptr_deref_2979_load_3 ptr_deref_2994_load_0 ptr_deref_2994_load_1 ptr_deref_2994_load_2 ptr_deref_2994_load_3 ptr_deref_3064_load_0 ptr_deref_3064_load_1 ptr_deref_3064_load_2 ptr_deref_3064_load_3 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(191 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 11 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_2979_load_0_req_0,
        ptr_deref_2979_load_0_ack_0,
        ptr_deref_2979_load_0_req_1,
        ptr_deref_2979_load_0_ack_1,
        "ptr_deref_2979_load_0",
        "memory_space_5" ,
        ptr_deref_2979_data_0,
        ptr_deref_2979_word_address_0,
        "ptr_deref_2979_data_0",
        "ptr_deref_2979_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2979_load_1_req_0,
        ptr_deref_2979_load_1_ack_0,
        ptr_deref_2979_load_1_req_1,
        ptr_deref_2979_load_1_ack_1,
        "ptr_deref_2979_load_1",
        "memory_space_5" ,
        ptr_deref_2979_data_1,
        ptr_deref_2979_word_address_1,
        "ptr_deref_2979_data_1",
        "ptr_deref_2979_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2979_load_2_req_0,
        ptr_deref_2979_load_2_ack_0,
        ptr_deref_2979_load_2_req_1,
        ptr_deref_2979_load_2_ack_1,
        "ptr_deref_2979_load_2",
        "memory_space_5" ,
        ptr_deref_2979_data_2,
        ptr_deref_2979_word_address_2,
        "ptr_deref_2979_data_2",
        "ptr_deref_2979_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2979_load_3_req_0,
        ptr_deref_2979_load_3_ack_0,
        ptr_deref_2979_load_3_req_1,
        ptr_deref_2979_load_3_ack_1,
        "ptr_deref_2979_load_3",
        "memory_space_5" ,
        ptr_deref_2979_data_3,
        ptr_deref_2979_word_address_3,
        "ptr_deref_2979_data_3",
        "ptr_deref_2979_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2994_load_0_req_0,
        ptr_deref_2994_load_0_ack_0,
        ptr_deref_2994_load_0_req_1,
        ptr_deref_2994_load_0_ack_1,
        "ptr_deref_2994_load_0",
        "memory_space_5" ,
        ptr_deref_2994_data_0,
        ptr_deref_2994_word_address_0,
        "ptr_deref_2994_data_0",
        "ptr_deref_2994_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2994_load_1_req_0,
        ptr_deref_2994_load_1_ack_0,
        ptr_deref_2994_load_1_req_1,
        ptr_deref_2994_load_1_ack_1,
        "ptr_deref_2994_load_1",
        "memory_space_5" ,
        ptr_deref_2994_data_1,
        ptr_deref_2994_word_address_1,
        "ptr_deref_2994_data_1",
        "ptr_deref_2994_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2994_load_2_req_0,
        ptr_deref_2994_load_2_ack_0,
        ptr_deref_2994_load_2_req_1,
        ptr_deref_2994_load_2_ack_1,
        "ptr_deref_2994_load_2",
        "memory_space_5" ,
        ptr_deref_2994_data_2,
        ptr_deref_2994_word_address_2,
        "ptr_deref_2994_data_2",
        "ptr_deref_2994_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_2994_load_3_req_0,
        ptr_deref_2994_load_3_ack_0,
        ptr_deref_2994_load_3_req_1,
        ptr_deref_2994_load_3_ack_1,
        "ptr_deref_2994_load_3",
        "memory_space_5" ,
        ptr_deref_2994_data_3,
        ptr_deref_2994_word_address_3,
        "ptr_deref_2994_data_3",
        "ptr_deref_2994_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3064_load_0_req_0,
        ptr_deref_3064_load_0_ack_0,
        ptr_deref_3064_load_0_req_1,
        ptr_deref_3064_load_0_ack_1,
        "ptr_deref_3064_load_0",
        "memory_space_5" ,
        ptr_deref_3064_data_0,
        ptr_deref_3064_word_address_0,
        "ptr_deref_3064_data_0",
        "ptr_deref_3064_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3064_load_1_req_0,
        ptr_deref_3064_load_1_ack_0,
        ptr_deref_3064_load_1_req_1,
        ptr_deref_3064_load_1_ack_1,
        "ptr_deref_3064_load_1",
        "memory_space_5" ,
        ptr_deref_3064_data_1,
        ptr_deref_3064_word_address_1,
        "ptr_deref_3064_data_1",
        "ptr_deref_3064_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3064_load_2_req_0,
        ptr_deref_3064_load_2_ack_0,
        ptr_deref_3064_load_2_req_1,
        ptr_deref_3064_load_2_ack_1,
        "ptr_deref_3064_load_2",
        "memory_space_5" ,
        ptr_deref_3064_data_2,
        ptr_deref_3064_word_address_2,
        "ptr_deref_3064_data_2",
        "ptr_deref_3064_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3064_load_3_req_0,
        ptr_deref_3064_load_3_ack_0,
        ptr_deref_3064_load_3_req_1,
        ptr_deref_3064_load_3_ack_1,
        "ptr_deref_3064_load_3",
        "memory_space_5" ,
        ptr_deref_3064_data_3,
        ptr_deref_3064_word_address_3,
        "ptr_deref_3064_data_3",
        "ptr_deref_3064_word_address_3" -- 
      );
      reqL(11) <= ptr_deref_2979_load_0_req_0;
      reqL(10) <= ptr_deref_2979_load_1_req_0;
      reqL(9) <= ptr_deref_2979_load_2_req_0;
      reqL(8) <= ptr_deref_2979_load_3_req_0;
      reqL(7) <= ptr_deref_2994_load_0_req_0;
      reqL(6) <= ptr_deref_2994_load_1_req_0;
      reqL(5) <= ptr_deref_2994_load_2_req_0;
      reqL(4) <= ptr_deref_2994_load_3_req_0;
      reqL(3) <= ptr_deref_3064_load_0_req_0;
      reqL(2) <= ptr_deref_3064_load_1_req_0;
      reqL(1) <= ptr_deref_3064_load_2_req_0;
      reqL(0) <= ptr_deref_3064_load_3_req_0;
      ptr_deref_2979_load_0_ack_0 <= ackL(11);
      ptr_deref_2979_load_1_ack_0 <= ackL(10);
      ptr_deref_2979_load_2_ack_0 <= ackL(9);
      ptr_deref_2979_load_3_ack_0 <= ackL(8);
      ptr_deref_2994_load_0_ack_0 <= ackL(7);
      ptr_deref_2994_load_1_ack_0 <= ackL(6);
      ptr_deref_2994_load_2_ack_0 <= ackL(5);
      ptr_deref_2994_load_3_ack_0 <= ackL(4);
      ptr_deref_3064_load_0_ack_0 <= ackL(3);
      ptr_deref_3064_load_1_ack_0 <= ackL(2);
      ptr_deref_3064_load_2_ack_0 <= ackL(1);
      ptr_deref_3064_load_3_ack_0 <= ackL(0);
      reqR(11) <= ptr_deref_2979_load_0_req_1;
      reqR(10) <= ptr_deref_2979_load_1_req_1;
      reqR(9) <= ptr_deref_2979_load_2_req_1;
      reqR(8) <= ptr_deref_2979_load_3_req_1;
      reqR(7) <= ptr_deref_2994_load_0_req_1;
      reqR(6) <= ptr_deref_2994_load_1_req_1;
      reqR(5) <= ptr_deref_2994_load_2_req_1;
      reqR(4) <= ptr_deref_2994_load_3_req_1;
      reqR(3) <= ptr_deref_3064_load_0_req_1;
      reqR(2) <= ptr_deref_3064_load_1_req_1;
      reqR(1) <= ptr_deref_3064_load_2_req_1;
      reqR(0) <= ptr_deref_3064_load_3_req_1;
      ptr_deref_2979_load_0_ack_1 <= ackR(11);
      ptr_deref_2979_load_1_ack_1 <= ackR(10);
      ptr_deref_2979_load_2_ack_1 <= ackR(9);
      ptr_deref_2979_load_3_ack_1 <= ackR(8);
      ptr_deref_2994_load_0_ack_1 <= ackR(7);
      ptr_deref_2994_load_1_ack_1 <= ackR(6);
      ptr_deref_2994_load_2_ack_1 <= ackR(5);
      ptr_deref_2994_load_3_ack_1 <= ackR(4);
      ptr_deref_3064_load_0_ack_1 <= ackR(3);
      ptr_deref_3064_load_1_ack_1 <= ackR(2);
      ptr_deref_3064_load_2_ack_1 <= ackR(1);
      ptr_deref_3064_load_3_ack_1 <= ackR(0);
      data_in <= ptr_deref_2979_word_address_0 & ptr_deref_2979_word_address_1 & ptr_deref_2979_word_address_2 & ptr_deref_2979_word_address_3 & ptr_deref_2994_word_address_0 & ptr_deref_2994_word_address_1 & ptr_deref_2994_word_address_2 & ptr_deref_2994_word_address_3 & ptr_deref_3064_word_address_0 & ptr_deref_3064_word_address_1 & ptr_deref_3064_word_address_2 & ptr_deref_3064_word_address_3;
      ptr_deref_2979_data_0 <= data_out(95 downto 88);
      ptr_deref_2979_data_1 <= data_out(87 downto 80);
      ptr_deref_2979_data_2 <= data_out(79 downto 72);
      ptr_deref_2979_data_3 <= data_out(71 downto 64);
      ptr_deref_2994_data_0 <= data_out(63 downto 56);
      ptr_deref_2994_data_1 <= data_out(55 downto 48);
      ptr_deref_2994_data_2 <= data_out(47 downto 40);
      ptr_deref_2994_data_3 <= data_out(39 downto 32);
      ptr_deref_3064_data_0 <= data_out(31 downto 24);
      ptr_deref_3064_data_1 <= data_out(23 downto 16);
      ptr_deref_3064_data_2 <= data_out(15 downto 8);
      ptr_deref_3064_data_3 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 12,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 12,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_2947_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2947_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_2947_word_address_0) &  " data ptr_deref_2947_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_2947_data_0) severity note; --
        end if;
        if ptr_deref_2947_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_2947_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_2947_word_address_1) &  " data ptr_deref_2947_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_2947_data_1) severity note; --
        end if;
        if ptr_deref_3052_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3052_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3052_word_address_0) &  " data ptr_deref_3052_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3052_data_0) severity note; --
        end if;
        if ptr_deref_3052_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3052_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_3052_word_address_1) &  " data ptr_deref_3052_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_3052_data_1) severity note; --
        end if;
        if ptr_deref_3059_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3059_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3059_word_address_0) &  " data ptr_deref_3059_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3059_data_0) severity note; --
        end if;
        if ptr_deref_3059_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3059_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_3059_word_address_1) &  " data ptr_deref_3059_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_3059_data_1) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_2947_store_0 ptr_deref_2947_store_1 ptr_deref_3052_store_0 ptr_deref_3052_store_1 ptr_deref_3059_store_0 ptr_deref_3059_store_1 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(95 downto 0);
      signal data_in: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      -- 
    begin -- 
      reqL(5) <= ptr_deref_2947_store_0_req_0;
      reqL(4) <= ptr_deref_2947_store_1_req_0;
      reqL(3) <= ptr_deref_3052_store_0_req_0;
      reqL(2) <= ptr_deref_3052_store_1_req_0;
      reqL(1) <= ptr_deref_3059_store_0_req_0;
      reqL(0) <= ptr_deref_3059_store_1_req_0;
      ptr_deref_2947_store_0_ack_0 <= ackL(5);
      ptr_deref_2947_store_1_ack_0 <= ackL(4);
      ptr_deref_3052_store_0_ack_0 <= ackL(3);
      ptr_deref_3052_store_1_ack_0 <= ackL(2);
      ptr_deref_3059_store_0_ack_0 <= ackL(1);
      ptr_deref_3059_store_1_ack_0 <= ackL(0);
      reqR(5) <= ptr_deref_2947_store_0_req_1;
      reqR(4) <= ptr_deref_2947_store_1_req_1;
      reqR(3) <= ptr_deref_3052_store_0_req_1;
      reqR(2) <= ptr_deref_3052_store_1_req_1;
      reqR(1) <= ptr_deref_3059_store_0_req_1;
      reqR(0) <= ptr_deref_3059_store_1_req_1;
      ptr_deref_2947_store_0_ack_1 <= ackR(5);
      ptr_deref_2947_store_1_ack_1 <= ackR(4);
      ptr_deref_3052_store_0_ack_1 <= ackR(3);
      ptr_deref_3052_store_1_ack_1 <= ackR(2);
      ptr_deref_3059_store_0_ack_1 <= ackR(1);
      ptr_deref_3059_store_1_ack_1 <= ackR(0);
      addr_in <= ptr_deref_2947_word_address_0 & ptr_deref_2947_word_address_1 & ptr_deref_3052_word_address_0 & ptr_deref_3052_word_address_1 & ptr_deref_3059_word_address_0 & ptr_deref_3059_word_address_1;
      data_in <= ptr_deref_2947_data_0 & ptr_deref_2947_data_1 & ptr_deref_3052_data_0 & ptr_deref_3052_data_1 & ptr_deref_3059_data_0 & ptr_deref_3059_data_1;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 6,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 6,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_2925_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_2925_inst_ack_0 then -- 
            assert false report " ReadPipe to3_in0 to wire simple_obj_ref_2925_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_2925_inst_req_0;
      simple_obj_ref_2925_inst_ack_0 <= ack(0);
      simple_obj_ref_2925_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => to3_in0_pipe_read_req(0),
          oack => to3_in0_pipe_read_ack(0),
          odata => to3_in0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3070_inst_ack_0 then -- 
          assert false report " WritePipe tofpga_port_number from wire type_cast_3072_wire_constant value="  &  convert_slv_to_hex_string(type_cast_3072_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3070_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3070_inst_req_0;
      simple_obj_ref_3070_inst_ack_0 <= ack(0);
      data_in <= type_cast_3072_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga_port_number_pipe_write_req(0),
          oack => tofpga_port_number_pipe_write_ack(0),
          odata => tofpga_port_number_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3074_inst_ack_0 then -- 
          assert false report " WritePipe tofpga3_out0 from wire type_cast_3076_wire value="  &  convert_slv_to_hex_string(type_cast_3076_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_3074_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3074_inst_req_0;
      simple_obj_ref_3074_inst_ack_0 <= ack(0);
      data_in <= type_cast_3076_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => tofpga3_out0_pipe_write_req(0),
          oack => tofpga3_out0_pipe_write_ack(0),
          odata => tofpga3_out0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_2945_call call_stmt_3050_call call_stmt_3057_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(47 downto 0);
      signal data_out: std_logic_vector(47 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      reqL(2) <= call_stmt_2945_call_req_0;
      reqL(1) <= call_stmt_3050_call_req_0;
      reqL(0) <= call_stmt_3057_call_req_0;
      call_stmt_2945_call_ack_0 <= ackL(2);
      call_stmt_3050_call_ack_0 <= ackL(1);
      call_stmt_3057_call_ack_0 <= ackL(0);
      reqR(2) <= call_stmt_2945_call_req_1;
      reqR(1) <= call_stmt_3050_call_req_1;
      reqR(0) <= call_stmt_3057_call_req_1;
      call_stmt_2945_call_ack_1 <= ackR(2);
      call_stmt_3050_call_ack_1 <= ackR(1);
      call_stmt_3057_call_ack_1 <= ackR(0);
      data_in <= type_cast_2943_wire_constant & tmp16_3008 & tmp21_3047;
      tmp4_2945 <= data_out(47 downto 32);
      tmp22_3050 <= data_out(31 downto 16);
      tmp23_3057 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 48,
        owidth => 16,
        twidth => 2,
        nreqs => 3,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => ahir_glue_bswap_i16_call_reqs(0),
          ackR => ahir_glue_bswap_i16_call_acks(0),
          dataR => ahir_glue_bswap_i16_call_data(15 downto 0),
          tagR => ahir_glue_bswap_i16_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 16, owidth => 48, twidth => 2, nreqs => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => ahir_glue_bswap_i16_return_acks(0), -- cross-over
          ackL => ahir_glue_bswap_i16_return_reqs(0), -- cross-over
          dataL => ahir_glue_bswap_i16_return_data(15 downto 0),
          tagL => ahir_glue_bswap_i16_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity analyze_packet is -- 
  generic (tag_length : integer); 
  port ( -- 
    pkt : in  std_logic_vector(31 downto 0);
    buf : out  std_logic_vector(31 downto 0);
    wlen : out  std_logic_vector(15 downto 0);
    blen : out  std_logic_vector(15 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity analyze_packet;
architecture Default of analyze_packet is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal buf_buffer :  std_logic_vector(31 downto 0);
  signal wlen_buffer :  std_logic_vector(15 downto 0);
  signal blen_buffer :  std_logic_vector(15 downto 0);
  signal analyze_packet_CP_15576_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3115_addr_1_req_0 : boolean;
  signal type_cast_3099_inst_req_0 : boolean;
  signal type_cast_3099_inst_ack_0 : boolean;
  signal binary_3095_inst_req_0 : boolean;
  signal array_obj_ref_3111_root_address_inst_req_0 : boolean;
  signal binary_3095_inst_ack_0 : boolean;
  signal array_obj_ref_3111_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3111_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3111_root_address_inst_ack_1 : boolean;
  signal binary_3095_inst_req_1 : boolean;
  signal ptr_deref_3115_addr_0_ack_0 : boolean;
  signal ptr_deref_3115_addr_1_ack_1 : boolean;
  signal ptr_deref_3115_addr_0_req_0 : boolean;
  signal type_cast_3103_inst_req_0 : boolean;
  signal array_obj_ref_3111_final_reg_req_0 : boolean;
  signal binary_3095_inst_ack_1 : boolean;
  signal ptr_deref_3115_addr_0_req_1 : boolean;
  signal array_obj_ref_3111_final_reg_ack_0 : boolean;
  signal array_obj_ref_3111_base_resize_ack_0 : boolean;
  signal type_cast_3103_inst_ack_0 : boolean;
  signal ptr_deref_3115_load_0_req_0 : boolean;
  signal ptr_deref_3115_load_0_ack_0 : boolean;
  signal ptr_deref_3115_addr_1_ack_0 : boolean;
  signal ptr_deref_3115_addr_1_req_1 : boolean;
  signal simple_obj_ref_3105_inst_req_0 : boolean;
  signal ptr_deref_3115_addr_0_ack_1 : boolean;
  signal ptr_deref_3115_base_resize_req_0 : boolean;
  signal ptr_deref_3115_base_resize_ack_0 : boolean;
  signal type_cast_3089_inst_req_0 : boolean;
  signal ptr_deref_3115_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_3105_inst_ack_0 : boolean;
  signal ptr_deref_3115_root_address_inst_ack_0 : boolean;
  signal type_cast_3089_inst_ack_0 : boolean;
  signal array_obj_ref_3111_base_resize_req_0 : boolean;
  signal ptr_deref_3115_load_1_req_0 : boolean;
  signal ptr_deref_3115_load_1_ack_0 : boolean;
  signal ptr_deref_3115_load_0_req_1 : boolean;
  signal ptr_deref_3115_load_0_ack_1 : boolean;
  signal ptr_deref_3115_load_1_req_1 : boolean;
  signal ptr_deref_3115_load_1_ack_1 : boolean;
  signal ptr_deref_3115_gather_scatter_req_0 : boolean;
  signal ptr_deref_3115_gather_scatter_ack_0 : boolean;
  signal type_cast_3119_inst_req_0 : boolean;
  signal type_cast_3119_inst_ack_0 : boolean;
  signal array_obj_ref_3124_base_resize_req_0 : boolean;
  signal array_obj_ref_3124_base_resize_ack_0 : boolean;
  signal array_obj_ref_3124_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3124_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3124_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3124_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3124_final_reg_req_0 : boolean;
  signal array_obj_ref_3124_final_reg_ack_0 : boolean;
  signal ptr_deref_3128_base_resize_req_0 : boolean;
  signal ptr_deref_3128_base_resize_ack_0 : boolean;
  signal ptr_deref_3128_root_address_inst_req_0 : boolean;
  signal ptr_deref_3128_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3128_addr_0_req_0 : boolean;
  signal ptr_deref_3128_addr_0_ack_0 : boolean;
  signal ptr_deref_3128_addr_0_req_1 : boolean;
  signal ptr_deref_3128_addr_0_ack_1 : boolean;
  signal ptr_deref_3128_addr_1_req_0 : boolean;
  signal ptr_deref_3128_addr_1_ack_0 : boolean;
  signal ptr_deref_3128_addr_1_req_1 : boolean;
  signal ptr_deref_3128_addr_1_ack_1 : boolean;
  signal ptr_deref_3128_load_0_req_0 : boolean;
  signal ptr_deref_3128_load_0_ack_0 : boolean;
  signal ptr_deref_3128_load_1_req_0 : boolean;
  signal ptr_deref_3128_load_1_ack_0 : boolean;
  signal ptr_deref_3128_load_0_req_1 : boolean;
  signal ptr_deref_3128_load_0_ack_1 : boolean;
  signal ptr_deref_3128_load_1_req_1 : boolean;
  signal ptr_deref_3128_load_1_ack_1 : boolean;
  signal ptr_deref_3128_gather_scatter_req_0 : boolean;
  signal ptr_deref_3128_gather_scatter_ack_0 : boolean;
  signal type_cast_3132_inst_req_0 : boolean;
  signal type_cast_3132_inst_ack_0 : boolean;
  signal binary_3138_inst_req_0 : boolean;
  signal binary_3138_inst_ack_0 : boolean;
  signal binary_3138_inst_req_1 : boolean;
  signal binary_3138_inst_ack_1 : boolean;
  signal type_cast_3142_inst_req_0 : boolean;
  signal type_cast_3142_inst_ack_0 : boolean;
  signal type_cast_3146_inst_req_0 : boolean;
  signal type_cast_3146_inst_ack_0 : boolean;
  signal binary_3150_inst_req_0 : boolean;
  signal binary_3150_inst_ack_0 : boolean;
  signal binary_3150_inst_req_1 : boolean;
  signal binary_3150_inst_ack_1 : boolean;
  signal type_cast_3151_inst_req_0 : boolean;
  signal type_cast_3151_inst_ack_0 : boolean;
  signal binary_3156_inst_req_0 : boolean;
  signal binary_3156_inst_ack_0 : boolean;
  signal binary_3156_inst_req_1 : boolean;
  signal binary_3156_inst_ack_1 : boolean;
  signal type_cast_3160_inst_req_0 : boolean;
  signal type_cast_3160_inst_ack_0 : boolean;
  signal type_cast_3164_inst_req_0 : boolean;
  signal type_cast_3164_inst_ack_0 : boolean;
  signal array_obj_ref_3169_base_resize_req_0 : boolean;
  signal array_obj_ref_3169_base_resize_ack_0 : boolean;
  signal array_obj_ref_3169_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3169_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3169_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3169_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3169_final_reg_req_0 : boolean;
  signal array_obj_ref_3169_final_reg_ack_0 : boolean;
  signal ptr_deref_3173_base_resize_req_0 : boolean;
  signal ptr_deref_3173_base_resize_ack_0 : boolean;
  signal ptr_deref_3173_root_address_inst_req_0 : boolean;
  signal ptr_deref_3173_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3173_addr_0_req_0 : boolean;
  signal ptr_deref_3173_addr_0_ack_0 : boolean;
  signal ptr_deref_3173_addr_0_req_1 : boolean;
  signal ptr_deref_3173_addr_0_ack_1 : boolean;
  signal ptr_deref_3173_addr_1_req_0 : boolean;
  signal ptr_deref_3173_addr_1_ack_0 : boolean;
  signal ptr_deref_3173_addr_1_req_1 : boolean;
  signal ptr_deref_3173_addr_1_ack_1 : boolean;
  signal ptr_deref_3173_load_0_req_0 : boolean;
  signal ptr_deref_3173_load_0_ack_0 : boolean;
  signal ptr_deref_3173_load_1_req_0 : boolean;
  signal ptr_deref_3173_load_1_ack_0 : boolean;
  signal ptr_deref_3173_load_0_req_1 : boolean;
  signal ptr_deref_3173_load_0_ack_1 : boolean;
  signal ptr_deref_3173_load_1_req_1 : boolean;
  signal ptr_deref_3173_load_1_ack_1 : boolean;
  signal ptr_deref_3173_gather_scatter_req_0 : boolean;
  signal ptr_deref_3173_gather_scatter_ack_0 : boolean;
  signal type_cast_3177_inst_req_0 : boolean;
  signal type_cast_3177_inst_ack_0 : boolean;
  signal array_obj_ref_3182_base_resize_req_0 : boolean;
  signal array_obj_ref_3182_base_resize_ack_0 : boolean;
  signal array_obj_ref_3182_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3182_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3182_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3182_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3182_final_reg_req_0 : boolean;
  signal array_obj_ref_3182_final_reg_ack_0 : boolean;
  signal ptr_deref_3186_base_resize_req_0 : boolean;
  signal ptr_deref_3186_base_resize_ack_0 : boolean;
  signal ptr_deref_3186_root_address_inst_req_0 : boolean;
  signal ptr_deref_3186_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3186_addr_0_req_0 : boolean;
  signal ptr_deref_3186_addr_0_ack_0 : boolean;
  signal ptr_deref_3186_addr_0_req_1 : boolean;
  signal ptr_deref_3186_addr_0_ack_1 : boolean;
  signal ptr_deref_3186_addr_1_req_0 : boolean;
  signal ptr_deref_3186_addr_1_ack_0 : boolean;
  signal ptr_deref_3186_addr_1_req_1 : boolean;
  signal ptr_deref_3186_addr_1_ack_1 : boolean;
  signal ptr_deref_3186_load_0_req_0 : boolean;
  signal ptr_deref_3186_load_0_ack_0 : boolean;
  signal ptr_deref_3186_load_1_req_0 : boolean;
  signal ptr_deref_3186_load_1_ack_0 : boolean;
  signal ptr_deref_3186_load_0_req_1 : boolean;
  signal ptr_deref_3186_load_0_ack_1 : boolean;
  signal ptr_deref_3186_load_1_req_1 : boolean;
  signal ptr_deref_3186_load_1_ack_1 : boolean;
  signal ptr_deref_3186_gather_scatter_req_0 : boolean;
  signal ptr_deref_3186_gather_scatter_ack_0 : boolean;
  signal type_cast_3190_inst_req_0 : boolean;
  signal type_cast_3190_inst_ack_0 : boolean;
  signal binary_3196_inst_req_0 : boolean;
  signal binary_3196_inst_ack_0 : boolean;
  signal binary_3196_inst_req_1 : boolean;
  signal binary_3196_inst_ack_1 : boolean;
  signal type_cast_3200_inst_req_0 : boolean;
  signal type_cast_3200_inst_ack_0 : boolean;
  signal type_cast_3204_inst_req_0 : boolean;
  signal type_cast_3204_inst_ack_0 : boolean;
  signal binary_3208_inst_req_0 : boolean;
  signal binary_3208_inst_ack_0 : boolean;
  signal binary_3208_inst_req_1 : boolean;
  signal binary_3208_inst_ack_1 : boolean;
  signal type_cast_3209_inst_req_0 : boolean;
  signal type_cast_3209_inst_ack_0 : boolean;
  signal binary_3214_inst_req_0 : boolean;
  signal binary_3214_inst_ack_0 : boolean;
  signal binary_3214_inst_req_1 : boolean;
  signal binary_3214_inst_ack_1 : boolean;
  signal type_cast_3218_inst_req_0 : boolean;
  signal type_cast_3218_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  buf <= buf_buffer; 
  wlen <= wlen_buffer; 
  blen <= blen_buffer; 
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  analyze_packet_CP_15576: Block -- control-path 
    signal cp_elements: BooleanArray(190 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(190);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(190), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cpelement_group_1 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(3));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => type_cast_3089_inst_req_0); -- 
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(0);
    ack_15591_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3089_inst_ack_0, ack => cp_elements(4)); -- 
    cpelement_group_5 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(4) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(5),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => binary_3095_inst_req_0); -- 
    cp_elements(6) <= cp_elements(0);
    ra_15601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3095_inst_ack_0, ack => cp_elements(7)); -- 
    cr_15602_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => binary_3095_inst_req_1); -- 
    cp_elements(8) <= binary_3095_inst_ack_1;
    cpelement_group_9 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(10) & cp_elements(11));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(9),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15612_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => type_cast_3099_inst_req_0); -- 
    cp_elements(10) <= cp_elements(0);
    cp_elements(11) <= cp_elements(8);
    cp_elements(12) <= type_cast_3099_inst_ack_0;
    cpelement_group_13 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(15));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(13),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15622_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => type_cast_3103_inst_req_0); -- 
    cp_elements(14) <= cp_elements(0);
    cp_elements(15) <= cp_elements(8);
    ack_15623_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3103_inst_ack_0, ack => cp_elements(16)); -- 
    base_resize_req_15642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_3111_base_resize_req_0); -- 
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(12) & cp_elements(19));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(18) <= cp_elements(12);
    req_15630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => simple_obj_ref_3105_inst_req_0); -- 
    ack_15631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3105_inst_ack_0, ack => cp_elements(19)); -- 
    cp_elements(20) <= cp_elements(0);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(20) & cp_elements(24));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15655_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => array_obj_ref_3111_final_reg_req_0); -- 
    base_resize_ack_15643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3111_base_resize_ack_0, ack => cp_elements(22)); -- 
    plus_base_rr_15648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => array_obj_ref_3111_root_address_inst_req_0); -- 
    plus_base_ra_15649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3111_root_address_inst_ack_0, ack => cp_elements(23)); -- 
    plus_base_cr_15650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => array_obj_ref_3111_root_address_inst_req_1); -- 
    plus_base_ca_15651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3111_root_address_inst_ack_1, ack => cp_elements(24)); -- 
    final_reg_ack_15656_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3111_final_reg_ack_0, ack => cp_elements(25)); -- 
    base_resize_req_15669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(25), ack => ptr_deref_3115_base_resize_req_0); -- 
    base_resize_ack_15670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_base_resize_ack_0, ack => cp_elements(26)); -- 
    sum_rename_req_15674_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => ptr_deref_3115_root_address_inst_req_0); -- 
    cp_elements(27) <= ptr_deref_3115_root_address_inst_ack_0;
    cp_elements(28) <= cp_elements(27);
    rr_15682_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_3115_addr_0_req_0); -- 
    ra_15683_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_addr_0_ack_0, ack => cp_elements(29)); -- 
    cr_15684_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => ptr_deref_3115_addr_0_req_1); -- 
    ca_15685_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_addr_0_ack_1, ack => cp_elements(30)); -- 
    cp_elements(31) <= cp_elements(27);
    rr_15689_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_3115_addr_1_req_0); -- 
    ra_15690_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_addr_1_ack_0, ack => cp_elements(32)); -- 
    cr_15691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => ptr_deref_3115_addr_1_req_1); -- 
    ca_15692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_addr_1_ack_1, ack => cp_elements(33)); -- 
    cpelement_group_34 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(30) & cp_elements(33));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(34),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(35) <= cp_elements(34);
    rr_15702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => ptr_deref_3115_load_0_req_0); -- 
    ra_15703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_load_0_ack_0, ack => cp_elements(36)); -- 
    cp_elements(37) <= cp_elements(34);
    rr_15707_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_3115_load_1_req_0); -- 
    ra_15708_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_load_1_ack_0, ack => cp_elements(38)); -- 
    cpelement_group_39 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(36) & cp_elements(38));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(39),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(40) <= cp_elements(39);
    cr_15718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_3115_load_0_req_1); -- 
    ca_15719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_load_0_ack_1, ack => cp_elements(41)); -- 
    cp_elements(42) <= cp_elements(39);
    cr_15723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_3115_load_1_req_1); -- 
    ca_15724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_load_1_ack_1, ack => cp_elements(43)); -- 
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(41) & cp_elements(43));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_15725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => ptr_deref_3115_gather_scatter_req_0); -- 
    merge_ack_15726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3115_gather_scatter_ack_0, ack => cp_elements(45)); -- 
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(47) & cp_elements(48));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15735_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => type_cast_3119_inst_req_0); -- 
    cp_elements(47) <= cp_elements(0);
    cp_elements(48) <= cp_elements(17);
    ack_15736_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3119_inst_ack_0, ack => cp_elements(49)); -- 
    base_resize_req_15747_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => array_obj_ref_3124_base_resize_req_0); -- 
    cp_elements(50) <= cp_elements(0);
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(54));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => array_obj_ref_3124_final_reg_req_0); -- 
    base_resize_ack_15748_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3124_base_resize_ack_0, ack => cp_elements(52)); -- 
    plus_base_rr_15753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_3124_root_address_inst_req_0); -- 
    plus_base_ra_15754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3124_root_address_inst_ack_0, ack => cp_elements(53)); -- 
    plus_base_cr_15755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_3124_root_address_inst_req_1); -- 
    plus_base_ca_15756_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3124_root_address_inst_ack_1, ack => cp_elements(54)); -- 
    final_reg_ack_15761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3124_final_reg_ack_0, ack => cp_elements(55)); -- 
    base_resize_req_15774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => ptr_deref_3128_base_resize_req_0); -- 
    base_resize_ack_15775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_base_resize_ack_0, ack => cp_elements(56)); -- 
    sum_rename_req_15779_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(56), ack => ptr_deref_3128_root_address_inst_req_0); -- 
    cp_elements(57) <= ptr_deref_3128_root_address_inst_ack_0;
    cp_elements(58) <= cp_elements(57);
    rr_15787_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => ptr_deref_3128_addr_0_req_0); -- 
    ra_15788_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_addr_0_ack_0, ack => cp_elements(59)); -- 
    cr_15789_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => ptr_deref_3128_addr_0_req_1); -- 
    ca_15790_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_addr_0_ack_1, ack => cp_elements(60)); -- 
    cp_elements(61) <= cp_elements(57);
    rr_15794_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => ptr_deref_3128_addr_1_req_0); -- 
    ra_15795_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_addr_1_ack_0, ack => cp_elements(62)); -- 
    cr_15796_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_3128_addr_1_req_1); -- 
    ca_15797_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_addr_1_ack_1, ack => cp_elements(63)); -- 
    cpelement_group_64 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(60) & cp_elements(63));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(64),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(65) <= cp_elements(64);
    rr_15807_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_3128_load_0_req_0); -- 
    ra_15808_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_load_0_ack_0, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(64);
    rr_15812_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => ptr_deref_3128_load_1_req_0); -- 
    ra_15813_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_load_1_ack_0, ack => cp_elements(68)); -- 
    cpelement_group_69 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(66) & cp_elements(68));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(69),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(70) <= cp_elements(69);
    cr_15823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_3128_load_0_req_1); -- 
    ca_15824_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_load_0_ack_1, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(69);
    cr_15828_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_3128_load_1_req_1); -- 
    ca_15829_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_load_1_ack_1, ack => cp_elements(73)); -- 
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(73));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_15830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => ptr_deref_3128_gather_scatter_req_0); -- 
    merge_ack_15831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3128_gather_scatter_ack_0, ack => cp_elements(75)); -- 
    cpelement_group_76 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(77));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(76),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => type_cast_3132_inst_req_0); -- 
    cp_elements(77) <= cp_elements(0);
    ack_15841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3132_inst_ack_0, ack => cp_elements(78)); -- 
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(80));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => binary_3138_inst_req_0); -- 
    cp_elements(80) <= cp_elements(0);
    ra_15851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3138_inst_ack_0, ack => cp_elements(81)); -- 
    cr_15852_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => binary_3138_inst_req_1); -- 
    ca_15853_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3138_inst_ack_1, ack => cp_elements(82)); -- 
    cpelement_group_83 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(45) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(83),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => type_cast_3142_inst_req_0); -- 
    cp_elements(84) <= cp_elements(0);
    ack_15863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3142_inst_ack_0, ack => cp_elements(85)); -- 
    cpelement_group_86 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(87) & cp_elements(94));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(86),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => type_cast_3151_inst_req_0); -- 
    cp_elements(87) <= cp_elements(0);
    cpelement_group_88 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(92));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(88),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => binary_3150_inst_req_0); -- 
    cp_elements(89) <= cp_elements(0);
    cpelement_group_90 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(85) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(90),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => type_cast_3146_inst_req_0); -- 
    cp_elements(91) <= cp_elements(0);
    ack_15877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3146_inst_ack_0, ack => cp_elements(92)); -- 
    ra_15882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3150_inst_ack_0, ack => cp_elements(93)); -- 
    cr_15883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => binary_3150_inst_req_1); -- 
    ca_15884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3150_inst_ack_1, ack => cp_elements(94)); -- 
    ack_15889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3151_inst_ack_0, ack => cp_elements(95)); -- 
    cpelement_group_96 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(82) & cp_elements(95) & cp_elements(97));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(96),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_15899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => binary_3156_inst_req_0); -- 
    cp_elements(97) <= cp_elements(0);
    ra_15900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3156_inst_ack_0, ack => cp_elements(98)); -- 
    cr_15901_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => binary_3156_inst_req_1); -- 
    ca_15902_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3156_inst_ack_1, ack => cp_elements(99)); -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(99) & cp_elements(101));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(100), ack => type_cast_3160_inst_req_0); -- 
    cp_elements(101) <= cp_elements(0);
    ack_15912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3160_inst_ack_0, ack => cp_elements(102)); -- 
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(104) & cp_elements(105));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_15921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => type_cast_3164_inst_req_0); -- 
    cp_elements(104) <= cp_elements(0);
    cp_elements(105) <= cp_elements(17);
    ack_15922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3164_inst_ack_0, ack => cp_elements(106)); -- 
    base_resize_req_15933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => array_obj_ref_3169_base_resize_req_0); -- 
    cp_elements(107) <= cp_elements(0);
    cpelement_group_108 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(107) & cp_elements(111));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(108),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_15946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => array_obj_ref_3169_final_reg_req_0); -- 
    base_resize_ack_15934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3169_base_resize_ack_0, ack => cp_elements(109)); -- 
    plus_base_rr_15939_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => array_obj_ref_3169_root_address_inst_req_0); -- 
    plus_base_ra_15940_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3169_root_address_inst_ack_0, ack => cp_elements(110)); -- 
    plus_base_cr_15941_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => array_obj_ref_3169_root_address_inst_req_1); -- 
    plus_base_ca_15942_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3169_root_address_inst_ack_1, ack => cp_elements(111)); -- 
    final_reg_ack_15947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3169_final_reg_ack_0, ack => cp_elements(112)); -- 
    base_resize_req_15960_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => ptr_deref_3173_base_resize_req_0); -- 
    base_resize_ack_15961_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_base_resize_ack_0, ack => cp_elements(113)); -- 
    sum_rename_req_15965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_3173_root_address_inst_req_0); -- 
    cp_elements(114) <= ptr_deref_3173_root_address_inst_ack_0;
    cp_elements(115) <= cp_elements(114);
    rr_15973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(115), ack => ptr_deref_3173_addr_0_req_0); -- 
    ra_15974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_addr_0_ack_0, ack => cp_elements(116)); -- 
    cr_15975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(116), ack => ptr_deref_3173_addr_0_req_1); -- 
    ca_15976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_addr_0_ack_1, ack => cp_elements(117)); -- 
    cp_elements(118) <= cp_elements(114);
    rr_15980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => ptr_deref_3173_addr_1_req_0); -- 
    ra_15981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_addr_1_ack_0, ack => cp_elements(119)); -- 
    cr_15982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_3173_addr_1_req_1); -- 
    ca_15983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_addr_1_ack_1, ack => cp_elements(120)); -- 
    cpelement_group_121 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(117) & cp_elements(120));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(121),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(122) <= cp_elements(121);
    rr_15993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_3173_load_0_req_0); -- 
    ra_15994_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_load_0_ack_0, ack => cp_elements(123)); -- 
    cp_elements(124) <= cp_elements(121);
    rr_15998_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => ptr_deref_3173_load_1_req_0); -- 
    ra_15999_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_load_1_ack_0, ack => cp_elements(125)); -- 
    cpelement_group_126 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(125));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(127) <= cp_elements(126);
    cr_16009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(127), ack => ptr_deref_3173_load_0_req_1); -- 
    ca_16010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_load_0_ack_1, ack => cp_elements(128)); -- 
    cp_elements(129) <= cp_elements(126);
    cr_16014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => ptr_deref_3173_load_1_req_1); -- 
    ca_16015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_load_1_ack_1, ack => cp_elements(130)); -- 
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(128) & cp_elements(130));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_16016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => ptr_deref_3173_gather_scatter_req_0); -- 
    merge_ack_16017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3173_gather_scatter_ack_0, ack => cp_elements(132)); -- 
    cpelement_group_133 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(133),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => type_cast_3177_inst_req_0); -- 
    cp_elements(134) <= cp_elements(0);
    cp_elements(135) <= cp_elements(17);
    ack_16027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3177_inst_ack_0, ack => cp_elements(136)); -- 
    base_resize_req_16038_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => array_obj_ref_3182_base_resize_req_0); -- 
    cp_elements(137) <= cp_elements(0);
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(137) & cp_elements(141));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_16051_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => array_obj_ref_3182_final_reg_req_0); -- 
    base_resize_ack_16039_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3182_base_resize_ack_0, ack => cp_elements(139)); -- 
    plus_base_rr_16044_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(139), ack => array_obj_ref_3182_root_address_inst_req_0); -- 
    plus_base_ra_16045_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3182_root_address_inst_ack_0, ack => cp_elements(140)); -- 
    plus_base_cr_16046_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => array_obj_ref_3182_root_address_inst_req_1); -- 
    plus_base_ca_16047_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3182_root_address_inst_ack_1, ack => cp_elements(141)); -- 
    final_reg_ack_16052_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3182_final_reg_ack_0, ack => cp_elements(142)); -- 
    base_resize_req_16065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => ptr_deref_3186_base_resize_req_0); -- 
    base_resize_ack_16066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_base_resize_ack_0, ack => cp_elements(143)); -- 
    sum_rename_req_16070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(143), ack => ptr_deref_3186_root_address_inst_req_0); -- 
    cp_elements(144) <= ptr_deref_3186_root_address_inst_ack_0;
    cp_elements(145) <= cp_elements(144);
    rr_16078_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(145), ack => ptr_deref_3186_addr_0_req_0); -- 
    ra_16079_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_addr_0_ack_0, ack => cp_elements(146)); -- 
    cr_16080_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => ptr_deref_3186_addr_0_req_1); -- 
    ca_16081_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_addr_0_ack_1, ack => cp_elements(147)); -- 
    cp_elements(148) <= cp_elements(144);
    rr_16085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => ptr_deref_3186_addr_1_req_0); -- 
    ra_16086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_addr_1_ack_0, ack => cp_elements(149)); -- 
    cr_16087_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(149), ack => ptr_deref_3186_addr_1_req_1); -- 
    ca_16088_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_addr_1_ack_1, ack => cp_elements(150)); -- 
    cpelement_group_151 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(147) & cp_elements(150));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(151),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(152) <= cp_elements(151);
    rr_16098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(152), ack => ptr_deref_3186_load_0_req_0); -- 
    ra_16099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_load_0_ack_0, ack => cp_elements(153)); -- 
    cp_elements(154) <= cp_elements(151);
    rr_16103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => ptr_deref_3186_load_1_req_0); -- 
    ra_16104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_load_1_ack_0, ack => cp_elements(155)); -- 
    cpelement_group_156 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(153) & cp_elements(155));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(156),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(157) <= cp_elements(156);
    cr_16114_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => ptr_deref_3186_load_0_req_1); -- 
    ca_16115_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_load_0_ack_1, ack => cp_elements(158)); -- 
    cp_elements(159) <= cp_elements(156);
    cr_16119_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(159), ack => ptr_deref_3186_load_1_req_1); -- 
    ca_16120_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_load_1_ack_1, ack => cp_elements(160)); -- 
    cpelement_group_161 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(158) & cp_elements(160));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(161),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_16121_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => ptr_deref_3186_gather_scatter_req_0); -- 
    merge_ack_16122_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3186_gather_scatter_ack_0, ack => cp_elements(162)); -- 
    cpelement_group_163 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(162) & cp_elements(164));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(163),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16131_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => type_cast_3190_inst_req_0); -- 
    cp_elements(164) <= cp_elements(0);
    ack_16132_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3190_inst_ack_0, ack => cp_elements(165)); -- 
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(165) & cp_elements(167));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => binary_3196_inst_req_0); -- 
    cp_elements(167) <= cp_elements(0);
    ra_16142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3196_inst_ack_0, ack => cp_elements(168)); -- 
    cr_16143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(168), ack => binary_3196_inst_req_1); -- 
    ca_16144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3196_inst_ack_1, ack => cp_elements(169)); -- 
    cpelement_group_170 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(171));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(170),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16153_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(170), ack => type_cast_3200_inst_req_0); -- 
    cp_elements(171) <= cp_elements(0);
    ack_16154_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3200_inst_ack_0, ack => cp_elements(172)); -- 
    cpelement_group_173 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(174) & cp_elements(181));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(173),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16179_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => type_cast_3209_inst_req_0); -- 
    cp_elements(174) <= cp_elements(0);
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(176) & cp_elements(179));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(175), ack => binary_3208_inst_req_0); -- 
    cp_elements(176) <= cp_elements(0);
    cpelement_group_177 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(172) & cp_elements(178));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(177), ack => type_cast_3204_inst_req_0); -- 
    cp_elements(178) <= cp_elements(0);
    ack_16168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3204_inst_ack_0, ack => cp_elements(179)); -- 
    ra_16173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3208_inst_ack_0, ack => cp_elements(180)); -- 
    cr_16174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_3208_inst_req_1); -- 
    ca_16175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3208_inst_ack_1, ack => cp_elements(181)); -- 
    ack_16180_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3209_inst_ack_0, ack => cp_elements(182)); -- 
    cpelement_group_183 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(169) & cp_elements(182) & cp_elements(184));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(183),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => binary_3214_inst_req_0); -- 
    cp_elements(184) <= cp_elements(0);
    ra_16191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3214_inst_ack_0, ack => cp_elements(185)); -- 
    cr_16192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => binary_3214_inst_req_1); -- 
    ca_16193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3214_inst_ack_1, ack => cp_elements(186)); -- 
    cpelement_group_187 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(186) & cp_elements(188));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(187),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16202_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => type_cast_3218_inst_req_0); -- 
    cp_elements(188) <= cp_elements(0);
    ack_16203_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3218_inst_ack_0, ack => cp_elements(189)); -- 
    cpelement_group_190 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(102) & cp_elements(189));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(190),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal addx_xptr16_3125 : std_logic_vector(31 downto 0);
    signal addx_xptr25_3170 : std_logic_vector(31 downto 0);
    signal addx_xptr29_3183 : std_logic_vector(31 downto 0);
    signal addx_xptr_3112 : std_logic_vector(31 downto 0);
    signal and_3096 : std_logic_vector(31 downto 0);
    signal array_obj_ref_3111_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3111_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3111_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3124_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3124_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3124_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3169_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3169_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3169_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3182_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3182_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3182_root_address : std_logic_vector(15 downto 0);
    signal binary_3150_wire : std_logic_vector(31 downto 0);
    signal binary_3208_wire : std_logic_vector(31 downto 0);
    signal blen_h_3174 : std_logic_vector(15 downto 0);
    signal blen_l_3187 : std_logic_vector(15 downto 0);
    signal conv21_3143 : std_logic_vector(31 downto 0);
    signal conv33_3191 : std_logic_vector(31 downto 0);
    signal conv36_3201 : std_logic_vector(31 downto 0);
    signal conv_3133 : std_logic_vector(31 downto 0);
    signal iNsTr_11_3120 : std_logic_vector(31 downto 0);
    signal iNsTr_14_3165 : std_logic_vector(31 downto 0);
    signal iNsTr_16_3178 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3090 : std_logic_vector(31 downto 0);
    signal iNsTr_7_3100 : std_logic_vector(31 downto 0);
    signal iNsTr_9_3104 : std_logic_vector(31 downto 0);
    signal or38_3215 : std_logic_vector(31 downto 0);
    signal or_3157 : std_logic_vector(31 downto 0);
    signal ptr_deref_3115_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3115_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3115_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3115_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3115_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3115_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3115_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3115_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3128_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3128_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3128_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3173_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3173_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3173_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3186_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3186_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3186_word_offset_1 : std_logic_vector(15 downto 0);
    signal shl34_3197 : std_logic_vector(31 downto 0);
    signal shl_3139 : std_logic_vector(31 downto 0);
    signal shr37_3210 : std_logic_vector(31 downto 0);
    signal shr_3152 : std_logic_vector(31 downto 0);
    signal type_cast_3094_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3137_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3146_wire : std_logic_vector(31 downto 0);
    signal type_cast_3149_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3195_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3204_wire : std_logic_vector(31 downto 0);
    signal type_cast_3207_wire_constant : std_logic_vector(31 downto 0);
    signal wlen_h_3116 : std_logic_vector(15 downto 0);
    signal wlen_l_3129 : std_logic_vector(15 downto 0);
    -- 
  begin -- 
    array_obj_ref_3111_final_offset <= "0000000000000010";
    array_obj_ref_3124_final_offset <= "0000000000000010";
    array_obj_ref_3169_final_offset <= "0000000000000110";
    array_obj_ref_3182_final_offset <= "0000000000000110";
    ptr_deref_3115_word_offset_0 <= "0000000000000000";
    ptr_deref_3115_word_offset_1 <= "0000000000000001";
    ptr_deref_3128_word_offset_0 <= "0000000000000000";
    ptr_deref_3128_word_offset_1 <= "0000000000000001";
    ptr_deref_3173_word_offset_0 <= "0000000000000000";
    ptr_deref_3173_word_offset_1 <= "0000000000000001";
    ptr_deref_3186_word_offset_0 <= "0000000000000000";
    ptr_deref_3186_word_offset_1 <= "0000000000000001";
    type_cast_3094_wire_constant <= "11111111111111111111100000000000";
    type_cast_3137_wire_constant <= "00000000000000000000000000001000";
    type_cast_3149_wire_constant <= "00000000000000000000000000001000";
    type_cast_3195_wire_constant <= "00000000000000000000000000001000";
    type_cast_3207_wire_constant <= "00000000000000000000000000001000";
    array_obj_ref_3111_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_9_3104, dout => array_obj_ref_3111_resized_base_address, req => array_obj_ref_3111_base_resize_req_0, ack => array_obj_ref_3111_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3111_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3111_root_address, dout => addx_xptr_3112, req => array_obj_ref_3111_final_reg_req_0, ack => array_obj_ref_3111_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3124_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_11_3120, dout => array_obj_ref_3124_resized_base_address, req => array_obj_ref_3124_base_resize_req_0, ack => array_obj_ref_3124_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3124_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3124_root_address, dout => addx_xptr16_3125, req => array_obj_ref_3124_final_reg_req_0, ack => array_obj_ref_3124_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3169_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_14_3165, dout => array_obj_ref_3169_resized_base_address, req => array_obj_ref_3169_base_resize_req_0, ack => array_obj_ref_3169_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3169_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3169_root_address, dout => addx_xptr25_3170, req => array_obj_ref_3169_final_reg_req_0, ack => array_obj_ref_3169_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3182_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_16_3178, dout => array_obj_ref_3182_resized_base_address, req => array_obj_ref_3182_base_resize_req_0, ack => array_obj_ref_3182_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3182_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3182_root_address, dout => addx_xptr29_3183, req => array_obj_ref_3182_final_reg_req_0, ack => array_obj_ref_3182_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3115_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr_3112, dout => ptr_deref_3115_resized_base_address, req => ptr_deref_3115_base_resize_req_0, ack => ptr_deref_3115_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3128_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr16_3125, dout => ptr_deref_3128_resized_base_address, req => ptr_deref_3128_base_resize_req_0, ack => ptr_deref_3128_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3173_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr25_3170, dout => ptr_deref_3173_resized_base_address, req => ptr_deref_3173_base_resize_req_0, ack => ptr_deref_3173_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3186_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => addx_xptr29_3183, dout => ptr_deref_3186_resized_base_address, req => ptr_deref_3186_base_resize_req_0, ack => ptr_deref_3186_base_resize_ack_0, clk => clk, reset => reset); -- 
    simple_obj_ref_3105_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_7_3100, dout => buf_buffer, req => simple_obj_ref_3105_inst_req_0, ack => simple_obj_ref_3105_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3089_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => pkt, dout => iNsTr_6_3090, req => type_cast_3089_inst_req_0, ack => type_cast_3089_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3099_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => and_3096, dout => iNsTr_7_3100, req => type_cast_3099_inst_req_0, ack => type_cast_3099_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3103_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => and_3096, dout => iNsTr_9_3104, req => type_cast_3103_inst_req_0, ack => type_cast_3103_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3119_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_11_3120, req => type_cast_3119_inst_req_0, ack => type_cast_3119_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3132_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => wlen_l_3129, dout => conv_3133, req => type_cast_3132_inst_req_0, ack => type_cast_3132_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3142_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => wlen_h_3116, dout => conv21_3143, req => type_cast_3142_inst_req_0, ack => type_cast_3142_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3146_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => conv21_3143, dout => type_cast_3146_wire, req => type_cast_3146_inst_req_0, ack => type_cast_3146_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3151_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => binary_3150_wire, dout => shr_3152, req => type_cast_3151_inst_req_0, ack => type_cast_3151_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3160_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => or_3157, dout => wlen_buffer, req => type_cast_3160_inst_req_0, ack => type_cast_3160_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3164_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_14_3165, req => type_cast_3164_inst_req_0, ack => type_cast_3164_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3177_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_buffer, dout => iNsTr_16_3178, req => type_cast_3177_inst_req_0, ack => type_cast_3177_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3190_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => blen_l_3187, dout => conv33_3191, req => type_cast_3190_inst_req_0, ack => type_cast_3190_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3200_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => blen_h_3174, dout => conv36_3201, req => type_cast_3200_inst_req_0, ack => type_cast_3200_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3204_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => conv36_3201, dout => type_cast_3204_wire, req => type_cast_3204_inst_req_0, ack => type_cast_3204_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3209_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => binary_3208_wire, dout => shr37_3210, req => type_cast_3209_inst_req_0, ack => type_cast_3209_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3218_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => false ) 
      port map( din => or38_3215, dout => blen_buffer, req => type_cast_3218_inst_req_0, ack => type_cast_3218_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3115_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3115_gather_scatter_ack_0 <= ptr_deref_3115_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3115_data_1 & ptr_deref_3115_data_0;
      wlen_h_3116 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3115_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3115_root_address_inst_ack_0 <= ptr_deref_3115_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3115_resized_base_address;
      ptr_deref_3115_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3128_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3128_gather_scatter_ack_0 <= ptr_deref_3128_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3128_data_1 & ptr_deref_3128_data_0;
      wlen_l_3129 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3128_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3128_root_address_inst_ack_0 <= ptr_deref_3128_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3128_resized_base_address;
      ptr_deref_3128_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3173_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3173_gather_scatter_ack_0 <= ptr_deref_3173_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3173_data_1 & ptr_deref_3173_data_0;
      blen_h_3174 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3173_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3173_root_address_inst_ack_0 <= ptr_deref_3173_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3173_resized_base_address;
      ptr_deref_3173_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3186_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3186_gather_scatter_ack_0 <= ptr_deref_3186_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3186_data_1 & ptr_deref_3186_data_0;
      blen_l_3187 <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3186_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3186_root_address_inst_ack_0 <= ptr_deref_3186_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3186_resized_base_address;
      ptr_deref_3186_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    -- shared split operator group (0) : array_obj_ref_3111_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3111_resized_base_address;
      array_obj_ref_3111_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3111_root_address_inst_req_0,
          ackL => array_obj_ref_3111_root_address_inst_ack_0,
          reqR => array_obj_ref_3111_root_address_inst_req_1,
          ackR => array_obj_ref_3111_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_3124_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3124_resized_base_address;
      array_obj_ref_3124_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3124_root_address_inst_req_0,
          ackL => array_obj_ref_3124_root_address_inst_ack_0,
          reqR => array_obj_ref_3124_root_address_inst_req_1,
          ackR => array_obj_ref_3124_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_3169_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3169_resized_base_address;
      array_obj_ref_3169_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3169_root_address_inst_req_0,
          ackL => array_obj_ref_3169_root_address_inst_ack_0,
          reqR => array_obj_ref_3169_root_address_inst_req_1,
          ackR => array_obj_ref_3169_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : array_obj_ref_3182_root_address_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3182_resized_base_address;
      array_obj_ref_3182_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3182_root_address_inst_req_0,
          ackL => array_obj_ref_3182_root_address_inst_ack_0,
          reqR => array_obj_ref_3182_root_address_inst_req_1,
          ackR => array_obj_ref_3182_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_3095_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_6_3090;
      and_3096 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3095_inst_req_0,
          ackL => binary_3095_inst_ack_0,
          reqR => binary_3095_inst_req_1,
          ackR => binary_3095_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_3138_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= conv_3133;
      shl_3139 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3138_inst_req_0,
          ackL => binary_3138_inst_ack_0,
          reqR => binary_3138_inst_req_1,
          ackR => binary_3138_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_3150_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3146_wire;
      binary_3150_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntASHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3150_inst_req_0,
          ackL => binary_3150_inst_ack_0,
          reqR => binary_3150_inst_req_1,
          ackR => binary_3150_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_3156_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= shl_3139 & shr_3152;
      or_3157 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3156_inst_req_0,
          ackL => binary_3156_inst_ack_0,
          reqR => binary_3156_inst_req_1,
          ackR => binary_3156_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_3196_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= conv33_3191;
      shl34_3197 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3196_inst_req_0,
          ackL => binary_3196_inst_ack_0,
          reqR => binary_3196_inst_req_1,
          ackR => binary_3196_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_3208_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3204_wire;
      binary_3208_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntASHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3208_inst_req_0,
          ackL => binary_3208_inst_ack_0,
          reqR => binary_3208_inst_req_1,
          ackR => binary_3208_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_3214_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= shl34_3197 & shr37_3210;
      or38_3215 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3214_inst_req_0,
          ackL => binary_3214_inst_ack_0,
          reqR => binary_3214_inst_req_1,
          ackR => binary_3214_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : ptr_deref_3115_addr_0 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3115_root_address;
      ptr_deref_3115_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3115_addr_0_req_0,
          ackL => ptr_deref_3115_addr_0_ack_0,
          reqR => ptr_deref_3115_addr_0_req_1,
          ackR => ptr_deref_3115_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : ptr_deref_3115_addr_1 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3115_root_address;
      ptr_deref_3115_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3115_addr_1_req_0,
          ackL => ptr_deref_3115_addr_1_ack_0,
          reqR => ptr_deref_3115_addr_1_req_1,
          ackR => ptr_deref_3115_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : ptr_deref_3128_addr_0 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3128_root_address;
      ptr_deref_3128_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3128_addr_0_req_0,
          ackL => ptr_deref_3128_addr_0_ack_0,
          reqR => ptr_deref_3128_addr_0_req_1,
          ackR => ptr_deref_3128_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : ptr_deref_3128_addr_1 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3128_root_address;
      ptr_deref_3128_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3128_addr_1_req_0,
          ackL => ptr_deref_3128_addr_1_ack_0,
          reqR => ptr_deref_3128_addr_1_req_1,
          ackR => ptr_deref_3128_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : ptr_deref_3173_addr_0 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3173_root_address;
      ptr_deref_3173_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3173_addr_0_req_0,
          ackL => ptr_deref_3173_addr_0_ack_0,
          reqR => ptr_deref_3173_addr_0_req_1,
          ackR => ptr_deref_3173_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : ptr_deref_3173_addr_1 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3173_root_address;
      ptr_deref_3173_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3173_addr_1_req_0,
          ackL => ptr_deref_3173_addr_1_ack_0,
          reqR => ptr_deref_3173_addr_1_req_1,
          ackR => ptr_deref_3173_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : ptr_deref_3186_addr_0 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3186_root_address;
      ptr_deref_3186_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3186_addr_0_req_0,
          ackL => ptr_deref_3186_addr_0_ack_0,
          reqR => ptr_deref_3186_addr_0_req_1,
          ackR => ptr_deref_3186_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : ptr_deref_3186_addr_1 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3186_root_address;
      ptr_deref_3186_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3186_addr_1_req_0,
          ackL => ptr_deref_3186_addr_1_ack_0,
          reqR => ptr_deref_3186_addr_1_req_1,
          ackR => ptr_deref_3186_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared load operator group (0) : ptr_deref_3128_load_1 ptr_deref_3115_load_0 ptr_deref_3115_load_1 ptr_deref_3186_load_0 ptr_deref_3128_load_0 ptr_deref_3173_load_0 ptr_deref_3173_load_1 ptr_deref_3186_load_1 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3128_load_1_req_0,
        ptr_deref_3128_load_1_ack_0,
        ptr_deref_3128_load_1_req_1,
        ptr_deref_3128_load_1_ack_1,
        "ptr_deref_3128_load_1",
        "memory_space_5" ,
        ptr_deref_3128_data_1,
        ptr_deref_3128_word_address_1,
        "ptr_deref_3128_data_1",
        "ptr_deref_3128_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3115_load_0_req_0,
        ptr_deref_3115_load_0_ack_0,
        ptr_deref_3115_load_0_req_1,
        ptr_deref_3115_load_0_ack_1,
        "ptr_deref_3115_load_0",
        "memory_space_5" ,
        ptr_deref_3115_data_0,
        ptr_deref_3115_word_address_0,
        "ptr_deref_3115_data_0",
        "ptr_deref_3115_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3115_load_1_req_0,
        ptr_deref_3115_load_1_ack_0,
        ptr_deref_3115_load_1_req_1,
        ptr_deref_3115_load_1_ack_1,
        "ptr_deref_3115_load_1",
        "memory_space_5" ,
        ptr_deref_3115_data_1,
        ptr_deref_3115_word_address_1,
        "ptr_deref_3115_data_1",
        "ptr_deref_3115_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3186_load_0_req_0,
        ptr_deref_3186_load_0_ack_0,
        ptr_deref_3186_load_0_req_1,
        ptr_deref_3186_load_0_ack_1,
        "ptr_deref_3186_load_0",
        "memory_space_5" ,
        ptr_deref_3186_data_0,
        ptr_deref_3186_word_address_0,
        "ptr_deref_3186_data_0",
        "ptr_deref_3186_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3128_load_0_req_0,
        ptr_deref_3128_load_0_ack_0,
        ptr_deref_3128_load_0_req_1,
        ptr_deref_3128_load_0_ack_1,
        "ptr_deref_3128_load_0",
        "memory_space_5" ,
        ptr_deref_3128_data_0,
        ptr_deref_3128_word_address_0,
        "ptr_deref_3128_data_0",
        "ptr_deref_3128_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3173_load_0_req_0,
        ptr_deref_3173_load_0_ack_0,
        ptr_deref_3173_load_0_req_1,
        ptr_deref_3173_load_0_ack_1,
        "ptr_deref_3173_load_0",
        "memory_space_5" ,
        ptr_deref_3173_data_0,
        ptr_deref_3173_word_address_0,
        "ptr_deref_3173_data_0",
        "ptr_deref_3173_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3173_load_1_req_0,
        ptr_deref_3173_load_1_ack_0,
        ptr_deref_3173_load_1_req_1,
        ptr_deref_3173_load_1_ack_1,
        "ptr_deref_3173_load_1",
        "memory_space_5" ,
        ptr_deref_3173_data_1,
        ptr_deref_3173_word_address_1,
        "ptr_deref_3173_data_1",
        "ptr_deref_3173_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3186_load_1_req_0,
        ptr_deref_3186_load_1_ack_0,
        ptr_deref_3186_load_1_req_1,
        ptr_deref_3186_load_1_ack_1,
        "ptr_deref_3186_load_1",
        "memory_space_5" ,
        ptr_deref_3186_data_1,
        ptr_deref_3186_word_address_1,
        "ptr_deref_3186_data_1",
        "ptr_deref_3186_word_address_1" -- 
      );
      reqL(7) <= ptr_deref_3128_load_1_req_0;
      reqL(6) <= ptr_deref_3115_load_0_req_0;
      reqL(5) <= ptr_deref_3115_load_1_req_0;
      reqL(4) <= ptr_deref_3186_load_0_req_0;
      reqL(3) <= ptr_deref_3128_load_0_req_0;
      reqL(2) <= ptr_deref_3173_load_0_req_0;
      reqL(1) <= ptr_deref_3173_load_1_req_0;
      reqL(0) <= ptr_deref_3186_load_1_req_0;
      ptr_deref_3128_load_1_ack_0 <= ackL(7);
      ptr_deref_3115_load_0_ack_0 <= ackL(6);
      ptr_deref_3115_load_1_ack_0 <= ackL(5);
      ptr_deref_3186_load_0_ack_0 <= ackL(4);
      ptr_deref_3128_load_0_ack_0 <= ackL(3);
      ptr_deref_3173_load_0_ack_0 <= ackL(2);
      ptr_deref_3173_load_1_ack_0 <= ackL(1);
      ptr_deref_3186_load_1_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_3128_load_1_req_1;
      reqR(6) <= ptr_deref_3115_load_0_req_1;
      reqR(5) <= ptr_deref_3115_load_1_req_1;
      reqR(4) <= ptr_deref_3186_load_0_req_1;
      reqR(3) <= ptr_deref_3128_load_0_req_1;
      reqR(2) <= ptr_deref_3173_load_0_req_1;
      reqR(1) <= ptr_deref_3173_load_1_req_1;
      reqR(0) <= ptr_deref_3186_load_1_req_1;
      ptr_deref_3128_load_1_ack_1 <= ackR(7);
      ptr_deref_3115_load_0_ack_1 <= ackR(6);
      ptr_deref_3115_load_1_ack_1 <= ackR(5);
      ptr_deref_3186_load_0_ack_1 <= ackR(4);
      ptr_deref_3128_load_0_ack_1 <= ackR(3);
      ptr_deref_3173_load_0_ack_1 <= ackR(2);
      ptr_deref_3173_load_1_ack_1 <= ackR(1);
      ptr_deref_3186_load_1_ack_1 <= ackR(0);
      data_in <= ptr_deref_3128_word_address_1 & ptr_deref_3115_word_address_0 & ptr_deref_3115_word_address_1 & ptr_deref_3186_word_address_0 & ptr_deref_3128_word_address_0 & ptr_deref_3173_word_address_0 & ptr_deref_3173_word_address_1 & ptr_deref_3186_word_address_1;
      ptr_deref_3128_data_1 <= data_out(63 downto 56);
      ptr_deref_3115_data_0 <= data_out(55 downto 48);
      ptr_deref_3115_data_1 <= data_out(47 downto 40);
      ptr_deref_3186_data_0 <= data_out(39 downto 32);
      ptr_deref_3128_data_0 <= data_out(31 downto 24);
      ptr_deref_3173_data_0 <= data_out(23 downto 16);
      ptr_deref_3173_data_1 <= data_out(15 downto 8);
      ptr_deref_3186_data_1 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 8,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity click_bc_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    GV_15_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
    GV_15_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
    GV_16_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity click_bc_storage_initializer_x;
architecture Default of click_bc_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal click_bc_storage_initializer_x_xCP_16204_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_3223_call_req_0 : boolean;
  signal call_stmt_3223_call_ack_0 : boolean;
  signal call_stmt_3223_call_req_1 : boolean;
  signal call_stmt_3223_call_ack_1 : boolean;
  signal call_stmt_3224_call_req_0 : boolean;
  signal call_stmt_3224_call_ack_0 : boolean;
  signal call_stmt_3224_call_req_1 : boolean;
  signal call_stmt_3224_call_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  click_bc_storage_initializer_x_xCP_16204: Block -- control-path 
    signal cp_elements: BooleanArray(7 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(7);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(7), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    crr_16218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_3223_call_req_0); -- 
    cra_16219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3223_call_ack_0, ack => cp_elements(2)); -- 
    ccr_16223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => call_stmt_3223_call_req_1); -- 
    cca_16224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3223_call_ack_1, ack => cp_elements(3)); -- 
    cp_elements(4) <= cp_elements(0);
    crr_16235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_3224_call_req_0); -- 
    cra_16236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3224_call_ack_0, ack => cp_elements(5)); -- 
    ccr_16240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_3224_call_req_1); -- 
    cca_16241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3224_call_ack_1, ack => cp_elements(6)); -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(6));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_3223_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3223_call_req_0;
      call_stmt_3223_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3223_call_req_1;
      call_stmt_3223_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => GV_15_initializer_in_click_bc_call_reqs(0),
          ackR => GV_15_initializer_in_click_bc_call_acks(0),
          tagR => GV_15_initializer_in_click_bc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => GV_15_initializer_in_click_bc_return_acks(0), -- cross-over
          ackL => GV_15_initializer_in_click_bc_return_reqs(0), -- cross-over
          tagL => GV_15_initializer_in_click_bc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_3224_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3224_call_req_0;
      call_stmt_3224_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3224_call_req_1;
      call_stmt_3224_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => GV_16_initializer_in_click_bc_call_reqs(0),
          ackR => GV_16_initializer_in_click_bc_call_acks(0),
          tagR => GV_16_initializer_in_click_bc_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => GV_16_initializer_in_click_bc_return_acks(0), -- cross-over
          ackL => GV_16_initializer_in_click_bc_return_reqs(0), -- cross-over
          tagL => GV_16_initializer_in_click_bc_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity free_queue_init is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity free_queue_init;
architecture Default of free_queue_init is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal free_queue_init_CP_16244_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3235_base_resize_req_0 : boolean;
  signal ptr_deref_3235_base_resize_ack_0 : boolean;
  signal ptr_deref_3235_root_address_inst_req_0 : boolean;
  signal ptr_deref_3235_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3235_addr_0_req_0 : boolean;
  signal ptr_deref_3235_addr_0_ack_0 : boolean;
  signal ptr_deref_3235_gather_scatter_req_0 : boolean;
  signal ptr_deref_3235_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3235_store_0_req_0 : boolean;
  signal ptr_deref_3235_store_0_ack_0 : boolean;
  signal ptr_deref_3235_store_0_req_1 : boolean;
  signal ptr_deref_3235_store_0_ack_1 : boolean;
  signal ptr_deref_3243_base_resize_req_0 : boolean;
  signal ptr_deref_3243_base_resize_ack_0 : boolean;
  signal ptr_deref_3243_root_address_inst_req_0 : boolean;
  signal ptr_deref_3243_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3243_addr_0_req_0 : boolean;
  signal ptr_deref_3243_addr_0_ack_0 : boolean;
  signal ptr_deref_3243_load_0_req_0 : boolean;
  signal ptr_deref_3243_load_0_ack_0 : boolean;
  signal ptr_deref_3243_load_0_req_1 : boolean;
  signal ptr_deref_3243_load_0_ack_1 : boolean;
  signal ptr_deref_3243_gather_scatter_req_0 : boolean;
  signal ptr_deref_3243_gather_scatter_ack_0 : boolean;
  signal type_cast_3247_inst_req_0 : boolean;
  signal type_cast_3247_inst_ack_0 : boolean;
  signal binary_3251_inst_req_0 : boolean;
  signal binary_3251_inst_ack_0 : boolean;
  signal binary_3251_inst_req_1 : boolean;
  signal binary_3251_inst_ack_1 : boolean;
  signal if_stmt_3253_branch_req_0 : boolean;
  signal if_stmt_3253_branch_ack_1 : boolean;
  signal if_stmt_3253_branch_ack_0 : boolean;
  signal ptr_deref_3262_base_resize_req_0 : boolean;
  signal ptr_deref_3262_base_resize_ack_0 : boolean;
  signal ptr_deref_3262_root_address_inst_req_0 : boolean;
  signal ptr_deref_3262_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3262_addr_0_req_0 : boolean;
  signal ptr_deref_3262_addr_0_ack_0 : boolean;
  signal ptr_deref_3262_load_0_req_0 : boolean;
  signal ptr_deref_3262_load_0_ack_0 : boolean;
  signal ptr_deref_3262_load_0_req_1 : boolean;
  signal ptr_deref_3262_load_0_ack_1 : boolean;
  signal ptr_deref_3262_gather_scatter_req_0 : boolean;
  signal ptr_deref_3262_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_3266_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3266_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_3266_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3266_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3266_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3266_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_3266_offset_inst_req_0 : boolean;
  signal array_obj_ref_3266_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3266_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3266_root_address_inst_ack_0 : boolean;
  signal addr_of_3267_final_reg_req_0 : boolean;
  signal addr_of_3267_final_reg_ack_0 : boolean;
  signal array_obj_ref_3274_base_resize_req_0 : boolean;
  signal array_obj_ref_3274_base_resize_ack_0 : boolean;
  signal array_obj_ref_3274_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3274_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3274_final_reg_req_0 : boolean;
  signal array_obj_ref_3274_final_reg_ack_0 : boolean;
  signal array_obj_ref_3281_base_resize_req_0 : boolean;
  signal array_obj_ref_3281_base_resize_ack_0 : boolean;
  signal array_obj_ref_3281_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3281_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3281_final_reg_req_0 : boolean;
  signal array_obj_ref_3281_final_reg_ack_0 : boolean;
  signal type_cast_3285_inst_req_0 : boolean;
  signal type_cast_3285_inst_ack_0 : boolean;
  signal simple_obj_ref_3287_inst_req_0 : boolean;
  signal simple_obj_ref_3287_inst_ack_0 : boolean;
  signal ptr_deref_3294_base_resize_req_0 : boolean;
  signal ptr_deref_3294_base_resize_ack_0 : boolean;
  signal ptr_deref_3294_root_address_inst_req_0 : boolean;
  signal ptr_deref_3294_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3294_addr_0_req_0 : boolean;
  signal ptr_deref_3294_addr_0_ack_0 : boolean;
  signal ptr_deref_3294_load_0_req_0 : boolean;
  signal ptr_deref_3294_load_0_ack_0 : boolean;
  signal ptr_deref_3294_load_0_req_1 : boolean;
  signal ptr_deref_3294_load_0_ack_1 : boolean;
  signal ptr_deref_3294_gather_scatter_req_0 : boolean;
  signal ptr_deref_3294_gather_scatter_ack_0 : boolean;
  signal binary_3300_inst_req_0 : boolean;
  signal binary_3300_inst_ack_0 : boolean;
  signal binary_3300_inst_req_1 : boolean;
  signal binary_3300_inst_ack_1 : boolean;
  signal ptr_deref_3303_base_resize_req_0 : boolean;
  signal ptr_deref_3303_base_resize_ack_0 : boolean;
  signal ptr_deref_3303_root_address_inst_req_0 : boolean;
  signal ptr_deref_3303_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3303_addr_0_req_0 : boolean;
  signal ptr_deref_3303_addr_0_ack_0 : boolean;
  signal ptr_deref_3303_gather_scatter_req_0 : boolean;
  signal ptr_deref_3303_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3303_store_0_req_0 : boolean;
  signal ptr_deref_3303_store_0_ack_0 : boolean;
  signal ptr_deref_3303_store_0_req_1 : boolean;
  signal ptr_deref_3303_store_0_ack_1 : boolean;
  signal memory_space_6_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_lr_tag : std_logic_vector(4 downto 0);
  signal memory_space_6_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_6_lc_tag :  std_logic_vector(1 downto 0);
  signal memory_space_6_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_6_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_6_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_6_sr_tag : std_logic_vector(4 downto 0);
  signal memory_space_6_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_6_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_6_sc_tag :  std_logic_vector(1 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  free_queue_init_CP_16244: Block -- control-path 
    signal cp_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(36);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(36), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= OrReduce(cp_elements(34) & cp_elements(91));
    cp_elements(2) <= cp_elements(0);
    cp_elements(3) <= cp_elements(2);
    cpelement_group_4 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(3) & cp_elements(5) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(4),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => ptr_deref_3235_gather_scatter_req_0); -- 
    cp_elements(5) <= cp_elements(2);
    cp_elements(6) <= cp_elements(5);
    base_resize_req_16289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => ptr_deref_3235_base_resize_req_0); -- 
    base_resize_ack_16290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_base_resize_ack_0, ack => cp_elements(7)); -- 
    sum_rename_req_16294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_3235_root_address_inst_req_0); -- 
    sum_rename_ack_16295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_root_address_inst_ack_0, ack => cp_elements(8)); -- 
    root_rename_req_16299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => ptr_deref_3235_addr_0_req_0); -- 
    root_rename_ack_16300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_addr_0_ack_0, ack => cp_elements(9)); -- 
    split_ack_16305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_gather_scatter_ack_0, ack => cp_elements(10)); -- 
    rr_16312_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_3235_store_0_req_0); -- 
    ra_16313_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_store_0_ack_0, ack => cp_elements(11)); -- 
    cr_16323_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => ptr_deref_3235_store_0_req_1); -- 
    ca_16324_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3235_store_0_ack_1, ack => cp_elements(12)); -- 
    cp_elements(13) <= cp_elements(89);
    cp_elements(14) <= cp_elements(13);
    base_resize_req_16340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => ptr_deref_3243_base_resize_req_0); -- 
    base_resize_ack_16341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_base_resize_ack_0, ack => cp_elements(15)); -- 
    sum_rename_req_16345_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => ptr_deref_3243_root_address_inst_req_0); -- 
    sum_rename_ack_16346_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_root_address_inst_ack_0, ack => cp_elements(16)); -- 
    root_rename_req_16350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_3243_addr_0_req_0); -- 
    root_rename_ack_16351_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_addr_0_ack_0, ack => cp_elements(17)); -- 
    rr_16361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_3243_load_0_req_0); -- 
    ra_16362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_load_0_ack_0, ack => cp_elements(18)); -- 
    cr_16372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_3243_load_0_req_1); -- 
    ca_16373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_load_0_ack_1, ack => cp_elements(19)); -- 
    merge_req_16374_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_3243_gather_scatter_req_0); -- 
    merge_ack_16375_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3243_gather_scatter_ack_0, ack => cp_elements(20)); -- 
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(25));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => binary_3251_inst_req_0); -- 
    cp_elements(22) <= cp_elements(13);
    cpelement_group_23 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(20) & cp_elements(24));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(23),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16386_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => type_cast_3247_inst_req_0); -- 
    cp_elements(24) <= cp_elements(13);
    ack_16387_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3247_inst_ack_0, ack => cp_elements(25)); -- 
    ra_16392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3251_inst_ack_0, ack => cp_elements(26)); -- 
    cr_16393_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_3251_inst_req_1); -- 
    ca_16394_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3251_inst_ack_1, ack => cp_elements(27)); -- 
    cp_elements(28) <= cp_elements(27);
    cp_elements(29) <= false;
    cp_elements(30) <= cp_elements(29);
    cp_elements(31) <= cp_elements(27);
    branch_req_16402_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => if_stmt_3253_branch_req_0); -- 
    cp_elements(32) <= cp_elements(31);
    cp_elements(33) <= cp_elements(32);
    if_choice_transition_16407_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3253_branch_ack_1, ack => cp_elements(34)); -- 
    cp_elements(35) <= cp_elements(32);
    else_choice_transition_16411_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3253_branch_ack_0, ack => cp_elements(36)); -- 
    cp_elements(37) <= cp_elements(1);
    cp_elements(38) <= cp_elements(37);
    base_resize_req_16429_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => ptr_deref_3262_base_resize_req_0); -- 
    base_resize_ack_16430_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_base_resize_ack_0, ack => cp_elements(39)); -- 
    sum_rename_req_16434_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => ptr_deref_3262_root_address_inst_req_0); -- 
    sum_rename_ack_16435_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_root_address_inst_ack_0, ack => cp_elements(40)); -- 
    root_rename_req_16439_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_3262_addr_0_req_0); -- 
    root_rename_ack_16440_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_addr_0_ack_0, ack => cp_elements(41)); -- 
    rr_16450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_3262_load_0_req_0); -- 
    ra_16451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_load_0_ack_0, ack => cp_elements(42)); -- 
    cr_16461_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => ptr_deref_3262_load_0_req_1); -- 
    ca_16462_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_load_0_ack_1, ack => cp_elements(43)); -- 
    merge_req_16463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => ptr_deref_3262_gather_scatter_req_0); -- 
    merge_ack_16464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3262_gather_scatter_ack_0, ack => cp_elements(44)); -- 
    index_resize_req_16478_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => array_obj_ref_3266_index_0_resize_req_0); -- 
    cpelement_group_45 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(46) & cp_elements(51));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(45),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_16500_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => addr_of_3267_final_reg_req_0); -- 
    cp_elements(46) <= cp_elements(37);
    index_resize_ack_16479_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3266_index_0_resize_ack_0, ack => cp_elements(47)); -- 
    scale_rr_16483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(47), ack => array_obj_ref_3266_index_0_scale_req_0); -- 
    scale_ra_16484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3266_index_0_scale_ack_0, ack => cp_elements(48)); -- 
    scale_cr_16485_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => array_obj_ref_3266_index_0_scale_req_1); -- 
    scale_ca_16486_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3266_index_0_scale_ack_1, ack => cp_elements(49)); -- 
    final_index_req_16490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => array_obj_ref_3266_offset_inst_req_0); -- 
    final_index_ack_16491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3266_offset_inst_ack_0, ack => cp_elements(50)); -- 
    sum_rename_req_16495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => array_obj_ref_3266_root_address_inst_req_0); -- 
    sum_rename_ack_16496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3266_root_address_inst_ack_0, ack => cp_elements(51)); -- 
    final_reg_ack_16501_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_3267_final_reg_ack_0, ack => cp_elements(52)); -- 
    base_resize_req_16512_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => array_obj_ref_3274_base_resize_req_0); -- 
    cp_elements(53) <= cp_elements(37);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_16522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => array_obj_ref_3274_final_reg_req_0); -- 
    base_resize_ack_16513_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3274_base_resize_ack_0, ack => cp_elements(55)); -- 
    sum_rename_req_16517_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => array_obj_ref_3274_root_address_inst_req_0); -- 
    sum_rename_ack_16518_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3274_root_address_inst_ack_0, ack => cp_elements(56)); -- 
    final_reg_ack_16523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3274_final_reg_ack_0, ack => cp_elements(57)); -- 
    base_resize_req_16534_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => array_obj_ref_3281_base_resize_req_0); -- 
    cp_elements(58) <= cp_elements(37);
    cpelement_group_59 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(58) & cp_elements(61));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(59),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_16544_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => array_obj_ref_3281_final_reg_req_0); -- 
    base_resize_ack_16535_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3281_base_resize_ack_0, ack => cp_elements(60)); -- 
    sum_rename_req_16539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => array_obj_ref_3281_root_address_inst_req_0); -- 
    sum_rename_ack_16540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3281_root_address_inst_ack_0, ack => cp_elements(61)); -- 
    final_reg_ack_16545_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3281_final_reg_ack_0, ack => cp_elements(62)); -- 
    cpelement_group_63 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(62) & cp_elements(64));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(63),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => type_cast_3285_inst_req_0); -- 
    cp_elements(64) <= cp_elements(37);
    ack_16555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3285_inst_ack_0, ack => cp_elements(65)); -- 
    pipe_wreq_16566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => simple_obj_ref_3287_inst_req_0); -- 
    pipe_wack_16567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3287_inst_ack_0, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(66);
    cp_elements(68) <= cp_elements(67);
    base_resize_req_16583_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_3294_base_resize_req_0); -- 
    base_resize_ack_16584_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_base_resize_ack_0, ack => cp_elements(69)); -- 
    sum_rename_req_16588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_3294_root_address_inst_req_0); -- 
    sum_rename_ack_16589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_root_address_inst_ack_0, ack => cp_elements(70)); -- 
    root_rename_req_16593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => ptr_deref_3294_addr_0_req_0); -- 
    root_rename_ack_16594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_addr_0_ack_0, ack => cp_elements(71)); -- 
    rr_16604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => ptr_deref_3294_load_0_req_0); -- 
    ra_16605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_load_0_ack_0, ack => cp_elements(72)); -- 
    cr_16615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => ptr_deref_3294_load_0_req_1); -- 
    ca_16616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_load_0_ack_1, ack => cp_elements(73)); -- 
    merge_req_16617_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => ptr_deref_3294_gather_scatter_req_0); -- 
    merge_ack_16618_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3294_gather_scatter_ack_0, ack => cp_elements(74)); -- 
    cpelement_group_75 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(75),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16627_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => binary_3300_inst_req_0); -- 
    cp_elements(76) <= cp_elements(67);
    ra_16628_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3300_inst_ack_0, ack => cp_elements(77)); -- 
    cr_16629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => binary_3300_inst_req_1); -- 
    ca_16630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3300_inst_ack_1, ack => cp_elements(78)); -- 
    cpelement_group_79 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(78) & cp_elements(80) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(79),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_16659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_3303_gather_scatter_req_0); -- 
    cp_elements(80) <= cp_elements(67);
    cp_elements(81) <= cp_elements(80);
    base_resize_req_16644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_3303_base_resize_req_0); -- 
    base_resize_ack_16645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_base_resize_ack_0, ack => cp_elements(82)); -- 
    sum_rename_req_16649_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => ptr_deref_3303_root_address_inst_req_0); -- 
    sum_rename_ack_16650_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_root_address_inst_ack_0, ack => cp_elements(83)); -- 
    root_rename_req_16654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_3303_addr_0_req_0); -- 
    root_rename_ack_16655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_addr_0_ack_0, ack => cp_elements(84)); -- 
    split_ack_16660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_gather_scatter_ack_0, ack => cp_elements(85)); -- 
    rr_16667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => ptr_deref_3303_store_0_req_0); -- 
    ra_16668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_store_0_ack_0, ack => cp_elements(86)); -- 
    cr_16678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(86), ack => ptr_deref_3303_store_0_req_1); -- 
    ca_16679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3303_store_0_ack_1, ack => cp_elements(87)); -- 
    cp_elements(88) <= OrReduce(cp_elements(12) & cp_elements(87));
    cp_elements(89) <= cp_elements(88);
    cp_elements(90) <= false;
    cp_elements(91) <= cp_elements(90);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_3266_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3266_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3266_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3266_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3274_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3274_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3281_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3281_root_address : std_logic_vector(15 downto 0);
    signal iNsTr_14_3295 : std_logic_vector(31 downto 0);
    signal iNsTr_15_3301 : std_logic_vector(31 downto 0);
    signal iNsTr_2_3244 : std_logic_vector(31 downto 0);
    signal iNsTr_3_3252 : std_logic_vector(0 downto 0);
    signal iNsTr_5_3263 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3268 : std_logic_vector(31 downto 0);
    signal iNsTr_7_3275 : std_logic_vector(31 downto 0);
    signal iNsTr_8_3282 : std_logic_vector(31 downto 0);
    signal iNsTr_9_3286 : std_logic_vector(31 downto 0);
    signal i_3233 : std_logic_vector(31 downto 0);
    signal ptr_deref_3235_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3235_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3235_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3235_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3235_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3235_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3243_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3243_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3243_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3243_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3243_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3262_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3262_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3262_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3262_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3262_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3294_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3294_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3294_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3294_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3294_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3303_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3303_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3303_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3303_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3303_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3303_word_offset_0 : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3265_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3265_scaled : std_logic_vector(15 downto 0);
    signal type_cast_3237_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3247_wire : std_logic_vector(31 downto 0);
    signal type_cast_3250_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_3299_wire_constant : std_logic_vector(31 downto 0);
    signal xxfree_queue_initxxbodyxxi_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_3266_offset_scale_factor_0 <= "0000100000000000";
    array_obj_ref_3266_resized_base_address <= "0000000000000000";
    i_3233 <= "00000000000000000000000000000000";
    ptr_deref_3235_word_offset_0 <= "0";
    ptr_deref_3243_word_offset_0 <= "0";
    ptr_deref_3262_word_offset_0 <= "0";
    ptr_deref_3294_word_offset_0 <= "0";
    ptr_deref_3303_word_offset_0 <= "0";
    type_cast_3237_wire_constant <= "00000000000000000000000000000000";
    type_cast_3250_wire_constant <= "00000000000000000000000000010000";
    type_cast_3299_wire_constant <= "00000000000000000000000000000001";
    xxfree_queue_initxxbodyxxi_alloc_base_address <= "0";
    addr_of_3267_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3266_root_address, dout => iNsTr_6_3268, req => addr_of_3267_final_reg_req_0, ack => addr_of_3267_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3266_index_0_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_5_3263, dout => simple_obj_ref_3265_resized, req => array_obj_ref_3266_index_0_resize_req_0, ack => array_obj_ref_3266_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3266_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3265_scaled, dout => array_obj_ref_3266_final_offset, req => array_obj_ref_3266_offset_inst_req_0, ack => array_obj_ref_3266_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3274_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_6_3268, dout => array_obj_ref_3274_resized_base_address, req => array_obj_ref_3274_base_resize_req_0, ack => array_obj_ref_3274_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3274_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3274_root_address, dout => iNsTr_7_3275, req => array_obj_ref_3274_final_reg_req_0, ack => array_obj_ref_3274_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3281_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => iNsTr_7_3275, dout => array_obj_ref_3281_resized_base_address, req => array_obj_ref_3281_base_resize_req_0, ack => array_obj_ref_3281_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3281_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3281_root_address, dout => iNsTr_8_3282, req => array_obj_ref_3281_final_reg_req_0, ack => array_obj_ref_3281_final_reg_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3235_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_3233, dout => ptr_deref_3235_resized_base_address, req => ptr_deref_3235_base_resize_req_0, ack => ptr_deref_3235_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3243_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_3233, dout => ptr_deref_3243_resized_base_address, req => ptr_deref_3243_base_resize_req_0, ack => ptr_deref_3243_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3262_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_3233, dout => ptr_deref_3262_resized_base_address, req => ptr_deref_3262_base_resize_req_0, ack => ptr_deref_3262_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3294_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_3233, dout => ptr_deref_3294_resized_base_address, req => ptr_deref_3294_base_resize_req_0, ack => ptr_deref_3294_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3303_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => i_3233, dout => ptr_deref_3303_resized_base_address, req => ptr_deref_3303_base_resize_req_0, ack => ptr_deref_3303_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_3247_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => iNsTr_2_3244, dout => type_cast_3247_wire, req => type_cast_3247_inst_req_0, ack => type_cast_3247_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3285_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_8_3282, dout => iNsTr_9_3286, req => type_cast_3285_inst_req_0, ack => type_cast_3285_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3266_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_3266_root_address_inst_ack_0 <= array_obj_ref_3266_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_3266_final_offset;
      array_obj_ref_3266_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_3274_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_3274_root_address_inst_ack_0 <= array_obj_ref_3274_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_3274_resized_base_address;
      array_obj_ref_3274_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    array_obj_ref_3281_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      array_obj_ref_3281_root_address_inst_ack_0 <= array_obj_ref_3281_root_address_inst_req_0;
      aggregated_sig <= array_obj_ref_3281_resized_base_address;
      array_obj_ref_3281_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    ptr_deref_3235_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3235_addr_0_ack_0 <= ptr_deref_3235_addr_0_req_0;
      aggregated_sig <= ptr_deref_3235_root_address;
      ptr_deref_3235_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3235_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3235_gather_scatter_ack_0 <= ptr_deref_3235_gather_scatter_req_0;
      aggregated_sig <= type_cast_3237_wire_constant;
      ptr_deref_3235_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3235_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3235_root_address_inst_ack_0 <= ptr_deref_3235_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3235_resized_base_address;
      ptr_deref_3235_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3243_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3243_addr_0_ack_0 <= ptr_deref_3243_addr_0_req_0;
      aggregated_sig <= ptr_deref_3243_root_address;
      ptr_deref_3243_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3243_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3243_gather_scatter_ack_0 <= ptr_deref_3243_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3243_data_0;
      iNsTr_2_3244 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3243_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3243_root_address_inst_ack_0 <= ptr_deref_3243_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3243_resized_base_address;
      ptr_deref_3243_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3262_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3262_addr_0_ack_0 <= ptr_deref_3262_addr_0_req_0;
      aggregated_sig <= ptr_deref_3262_root_address;
      ptr_deref_3262_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3262_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3262_gather_scatter_ack_0 <= ptr_deref_3262_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3262_data_0;
      iNsTr_5_3263 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3262_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3262_root_address_inst_ack_0 <= ptr_deref_3262_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3262_resized_base_address;
      ptr_deref_3262_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3294_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3294_addr_0_ack_0 <= ptr_deref_3294_addr_0_req_0;
      aggregated_sig <= ptr_deref_3294_root_address;
      ptr_deref_3294_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3294_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3294_gather_scatter_ack_0 <= ptr_deref_3294_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3294_data_0;
      iNsTr_14_3295 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3294_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3294_root_address_inst_ack_0 <= ptr_deref_3294_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3294_resized_base_address;
      ptr_deref_3294_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3303_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3303_addr_0_ack_0 <= ptr_deref_3303_addr_0_req_0;
      aggregated_sig <= ptr_deref_3303_root_address;
      ptr_deref_3303_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3303_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3303_gather_scatter_ack_0 <= ptr_deref_3303_gather_scatter_req_0;
      aggregated_sig <= iNsTr_15_3301;
      ptr_deref_3303_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3303_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3303_root_address_inst_ack_0 <= ptr_deref_3303_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3303_resized_base_address;
      ptr_deref_3303_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    if_stmt_3253_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= iNsTr_3_3252;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3253_branch_req_0,
          ack0 => if_stmt_3253_branch_ack_0,
          ack1 => if_stmt_3253_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_3266_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3265_resized;
      simple_obj_ref_3265_scaled <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000100000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3266_index_0_scale_req_0,
          ackL => array_obj_ref_3266_index_0_scale_ack_0,
          reqR => array_obj_ref_3266_index_0_scale_req_1,
          ackR => array_obj_ref_3266_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : binary_3251_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3247_wire;
      iNsTr_3_3252 <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000010000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3251_inst_req_0,
          ackL => binary_3251_inst_ack_0,
          reqR => binary_3251_inst_req_1,
          ackR => binary_3251_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : binary_3300_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_14_3295;
      iNsTr_15_3301 <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3300_inst_req_0,
          ackL => binary_3300_inst_ack_0,
          reqR => binary_3300_inst_req_1,
          ackR => binary_3300_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared load operator group (0) : ptr_deref_3294_load_0 ptr_deref_3243_load_0 ptr_deref_3262_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal data_out: std_logic_vector(95 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3294_load_0_req_0,
        ptr_deref_3294_load_0_ack_0,
        ptr_deref_3294_load_0_req_1,
        ptr_deref_3294_load_0_ack_1,
        "ptr_deref_3294_load_0",
        "memory_space_6" ,
        ptr_deref_3294_data_0,
        ptr_deref_3294_word_address_0,
        "ptr_deref_3294_data_0",
        "ptr_deref_3294_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3243_load_0_req_0,
        ptr_deref_3243_load_0_ack_0,
        ptr_deref_3243_load_0_req_1,
        ptr_deref_3243_load_0_ack_1,
        "ptr_deref_3243_load_0",
        "memory_space_6" ,
        ptr_deref_3243_data_0,
        ptr_deref_3243_word_address_0,
        "ptr_deref_3243_data_0",
        "ptr_deref_3243_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3262_load_0_req_0,
        ptr_deref_3262_load_0_ack_0,
        ptr_deref_3262_load_0_req_1,
        ptr_deref_3262_load_0_ack_1,
        "ptr_deref_3262_load_0",
        "memory_space_6" ,
        ptr_deref_3262_data_0,
        ptr_deref_3262_word_address_0,
        "ptr_deref_3262_data_0",
        "ptr_deref_3262_word_address_0" -- 
      );
      reqL(2) <= ptr_deref_3294_load_0_req_0;
      reqL(1) <= ptr_deref_3243_load_0_req_0;
      reqL(0) <= ptr_deref_3262_load_0_req_0;
      ptr_deref_3294_load_0_ack_0 <= ackL(2);
      ptr_deref_3243_load_0_ack_0 <= ackL(1);
      ptr_deref_3262_load_0_ack_0 <= ackL(0);
      reqR(2) <= ptr_deref_3294_load_0_req_1;
      reqR(1) <= ptr_deref_3243_load_0_req_1;
      reqR(0) <= ptr_deref_3262_load_0_req_1;
      ptr_deref_3294_load_0_ack_1 <= ackR(2);
      ptr_deref_3243_load_0_ack_1 <= ackR(1);
      ptr_deref_3262_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3294_word_address_0 & ptr_deref_3243_word_address_0 & ptr_deref_3262_word_address_0;
      ptr_deref_3294_data_0 <= data_out(95 downto 64);
      ptr_deref_3243_data_0 <= data_out(63 downto 32);
      ptr_deref_3262_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 3,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_6_lr_req(0),
          mack => memory_space_6_lr_ack(0),
          maddr => memory_space_6_lr_addr(0 downto 0),
          mtag => memory_space_6_lr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 3,  tag_length => 2,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_6_lc_req(0),
          mack => memory_space_6_lc_ack(0),
          mdata => memory_space_6_lc_data(31 downto 0),
          mtag => memory_space_6_lc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3303_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_6 address ptr_deref_3303_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3303_word_address_0) &  " data ptr_deref_3303_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3303_data_0) severity note; --
        end if;
        if ptr_deref_3235_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_6 address ptr_deref_3235_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3235_word_address_0) &  " data ptr_deref_3235_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3235_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3303_store_0 ptr_deref_3235_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(1 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      reqL(1) <= ptr_deref_3303_store_0_req_0;
      reqL(0) <= ptr_deref_3235_store_0_req_0;
      ptr_deref_3303_store_0_ack_0 <= ackL(1);
      ptr_deref_3235_store_0_ack_0 <= ackL(0);
      reqR(1) <= ptr_deref_3303_store_0_req_1;
      reqR(0) <= ptr_deref_3235_store_0_req_1;
      ptr_deref_3303_store_0_ack_1 <= ackR(1);
      ptr_deref_3235_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3303_word_address_0 & ptr_deref_3235_word_address_0;
      data_in <= ptr_deref_3303_data_0 & ptr_deref_3235_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 2,
        tag_length => 2,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_6_sr_req(0),
          mack => memory_space_6_sr_ack(0),
          maddr => memory_space_6_sr_addr(0 downto 0),
          mdata => memory_space_6_sr_data(31 downto 0),
          mtag => memory_space_6_sr_tag(4 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 2,
          tag_length => 2 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_6_sc_req(0),
          mack => memory_space_6_sc_ack(0),
          mtag => memory_space_6_sc_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3287_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire iNsTr_9_3286 value="  &  convert_slv_to_hex_string(iNsTr_9_3286) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3287_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3287_inst_req_0;
      simple_obj_ref_3287_inst_ack_0 <= ack(0);
      data_in <= iNsTr_9_3286;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_6: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 2,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_6_lr_addr,
      lr_req_in => memory_space_6_lr_req,
      lr_ack_out => memory_space_6_lr_ack,
      lr_tag_in => memory_space_6_lr_tag,
      lc_req_in => memory_space_6_lc_req,
      lc_ack_out => memory_space_6_lc_ack,
      lc_data_out => memory_space_6_lc_data,
      lc_tag_out => memory_space_6_lc_tag,
      sr_addr_in => memory_space_6_sr_addr,
      sr_data_in => memory_space_6_sr_data,
      sr_req_in => memory_space_6_sr_req,
      sr_ack_out => memory_space_6_sr_ack,
      sr_tag_in => memory_space_6_sr_tag,
      sc_req_in=> memory_space_6_sc_req,
      sc_ack_out => memory_space_6_sc_ack,
      sc_tag_out => memory_space_6_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity global_storage_initializer_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    click_bc_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    click_bc_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity global_storage_initializer_x;
architecture Default of global_storage_initializer_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal global_storage_initializer_x_xCP_16727_start: Boolean;
  -- links between control-path and data-path
  signal call_stmt_3314_call_req_1 : boolean;
  signal call_stmt_3314_call_ack_1 : boolean;
  signal call_stmt_3314_call_req_0 : boolean;
  signal call_stmt_3314_call_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  global_storage_initializer_x_xCP_16727: Block -- control-path 
    signal cp_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    crr_16741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => call_stmt_3314_call_req_0); -- 
    cra_16742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3314_call_ack_0, ack => cp_elements(1)); -- 
    ccr_16746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => call_stmt_3314_call_req_1); -- 
    cca_16747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3314_call_ack_1, ack => cp_elements(2)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- shared call operator group (0) : call_stmt_3314_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3314_call_req_0;
      call_stmt_3314_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3314_call_req_1;
      call_stmt_3314_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => click_bc_storage_initializer_x_call_reqs(0),
          ackR => click_bc_storage_initializer_x_call_acks(0),
          tagR => click_bc_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => click_bc_storage_initializer_x_return_acks(0), -- cross-over
          ackL => click_bc_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => click_bc_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity receive_packet_pipeline is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
    memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
    free_queue_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
    in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    receive_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
    swapped_in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    swapped_in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    swapped_in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
    receive_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
    receive_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
    swapped_in_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    swapped_in_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    swapped_in_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    receive_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity receive_packet_pipeline;
architecture Default of receive_packet_pipeline is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal receive_packet_pipeline_CP_16919_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_3425_inst_ack_0 : boolean;
  signal binary_3348_inst_req_0 : boolean;
  signal type_cast_3343_inst_ack_0 : boolean;
  signal type_cast_3347_inst_req_0 : boolean;
  signal binary_3352_inst_req_1 : boolean;
  signal simple_obj_ref_3330_inst_req_0 : boolean;
  signal type_cast_3347_inst_ack_0 : boolean;
  signal binary_3346_inst_ack_0 : boolean;
  signal binary_3346_inst_ack_1 : boolean;
  signal simple_obj_ref_3416_inst_req_0 : boolean;
  signal binary_3346_inst_req_0 : boolean;
  signal simple_obj_ref_3377_inst_req_0 : boolean;
  signal simple_obj_ref_3430_inst_req_0 : boolean;
  signal binary_3339_inst_req_0 : boolean;
  signal simple_obj_ref_3332_inst_req_0 : boolean;
  signal binary_3348_inst_ack_1 : boolean;
  signal simple_obj_ref_3416_inst_ack_0 : boolean;
  signal binary_3365_inst_req_1 : boolean;
  signal binary_3365_inst_ack_1 : boolean;
  signal simple_obj_ref_3402_inst_req_0 : boolean;
  signal binary_3339_inst_req_1 : boolean;
  signal binary_3339_inst_ack_0 : boolean;
  signal binary_3365_inst_ack_0 : boolean;
  signal array_obj_ref_3390_root_address_inst_req_0 : boolean;
  signal binary_3365_inst_req_0 : boolean;
  signal binary_3348_inst_ack_0 : boolean;
  signal type_cast_3343_inst_req_0 : boolean;
  signal simple_obj_ref_3406_inst_req_0 : boolean;
  signal array_obj_ref_3390_base_resize_ack_0 : boolean;
  signal type_cast_3362_inst_ack_0 : boolean;
  signal binary_3348_inst_req_1 : boolean;
  signal array_obj_ref_3390_root_address_inst_ack_1 : boolean;
  signal simple_obj_ref_3431_inst_ack_0 : boolean;
  signal type_cast_3386_inst_req_0 : boolean;
  signal array_obj_ref_3390_root_address_inst_req_1 : boolean;
  signal binary_3342_inst_ack_1 : boolean;
  signal simple_obj_ref_3332_inst_ack_0 : boolean;
  signal type_cast_3362_inst_req_0 : boolean;
  signal type_cast_3404_inst_ack_0 : boolean;
  signal type_cast_3386_inst_ack_0 : boolean;
  signal simple_obj_ref_3406_inst_ack_0 : boolean;
  signal binary_3349_inst_req_0 : boolean;
  signal type_cast_3404_inst_req_0 : boolean;
  signal binary_3339_inst_ack_1 : boolean;
  signal simple_obj_ref_3330_inst_ack_0 : boolean;
  signal binary_3346_inst_req_1 : boolean;
  signal type_cast_3366_inst_req_0 : boolean;
  signal type_cast_3366_inst_ack_0 : boolean;
  signal binary_3349_inst_ack_0 : boolean;
  signal binary_3349_inst_req_1 : boolean;
  signal simple_obj_ref_3431_inst_req_0 : boolean;
  signal binary_3349_inst_ack_1 : boolean;
  signal binary_3361_inst_ack_1 : boolean;
  signal type_cast_3353_inst_ack_0 : boolean;
  signal binary_3361_inst_req_1 : boolean;
  signal simple_obj_ref_3377_inst_ack_0 : boolean;
  signal binary_3352_inst_ack_1 : boolean;
  signal binary_3361_inst_ack_0 : boolean;
  signal type_cast_3353_inst_req_0 : boolean;
  signal binary_3361_inst_req_0 : boolean;
  signal binary_3352_inst_ack_0 : boolean;
  signal binary_3367_inst_req_0 : boolean;
  signal binary_3367_inst_ack_0 : boolean;
  signal binary_3367_inst_req_1 : boolean;
  signal binary_3367_inst_ack_1 : boolean;
  signal binary_3368_inst_req_0 : boolean;
  signal binary_3368_inst_ack_0 : boolean;
  signal array_obj_ref_3390_root_address_inst_ack_0 : boolean;
  signal type_cast_3334_inst_req_0 : boolean;
  signal type_cast_3334_inst_ack_0 : boolean;
  signal binary_3368_inst_req_1 : boolean;
  signal simple_obj_ref_3422_inst_req_0 : boolean;
  signal binary_3368_inst_ack_1 : boolean;
  signal simple_obj_ref_3399_inst_req_0 : boolean;
  signal simple_obj_ref_3399_inst_ack_0 : boolean;
  signal binary_3369_inst_req_0 : boolean;
  signal type_cast_3338_inst_req_0 : boolean;
  signal simple_obj_ref_3425_inst_req_0 : boolean;
  signal binary_3369_inst_ack_0 : boolean;
  signal simple_obj_ref_3422_inst_ack_0 : boolean;
  signal binary_3337_inst_req_0 : boolean;
  signal binary_3369_inst_req_1 : boolean;
  signal binary_3369_inst_ack_1 : boolean;
  signal type_cast_3338_inst_ack_0 : boolean;
  signal binary_3337_inst_ack_0 : boolean;
  signal binary_3337_inst_req_1 : boolean;
  signal binary_3337_inst_ack_1 : boolean;
  signal array_obj_ref_3390_base_resize_req_0 : boolean;
  signal binary_3352_inst_req_0 : boolean;
  signal simple_obj_ref_3440_inst_req_0 : boolean;
  signal binary_3342_inst_req_1 : boolean;
  signal simple_obj_ref_3436_inst_ack_0 : boolean;
  signal binary_3342_inst_ack_0 : boolean;
  signal type_cast_3382_inst_ack_0 : boolean;
  signal binary_3342_inst_req_0 : boolean;
  signal simple_obj_ref_3396_inst_ack_0 : boolean;
  signal binary_3358_inst_ack_1 : boolean;
  signal simple_obj_ref_3396_inst_req_0 : boolean;
  signal binary_3358_inst_req_1 : boolean;
  signal simple_obj_ref_3433_inst_ack_0 : boolean;
  signal if_stmt_3443_branch_req_0 : boolean;
  signal if_stmt_3443_branch_ack_0 : boolean;
  signal binary_3358_inst_ack_0 : boolean;
  signal if_stmt_3443_branch_ack_1 : boolean;
  signal binary_3446_inst_req_0 : boolean;
  signal simple_obj_ref_3402_inst_ack_0 : boolean;
  signal binary_3446_inst_ack_0 : boolean;
  signal binary_3446_inst_req_1 : boolean;
  signal binary_3446_inst_ack_1 : boolean;
  signal simple_obj_ref_3457_inst_req_0 : boolean;
  signal simple_obj_ref_3457_inst_ack_0 : boolean;
  signal simple_obj_ref_3458_inst_req_0 : boolean;
  signal simple_obj_ref_3458_inst_ack_0 : boolean;
  signal binary_3358_inst_req_0 : boolean;
  signal type_cast_3382_inst_req_0 : boolean;
  signal type_cast_3357_inst_ack_0 : boolean;
  signal type_cast_3357_inst_req_0 : boolean;
  signal binary_3356_inst_ack_1 : boolean;
  signal simple_obj_ref_3430_inst_ack_0 : boolean;
  signal binary_3356_inst_req_1 : boolean;
  signal simple_obj_ref_3419_inst_ack_0 : boolean;
  signal binary_3356_inst_ack_0 : boolean;
  signal simple_obj_ref_3393_inst_ack_0 : boolean;
  signal simple_obj_ref_3419_inst_req_0 : boolean;
  signal simple_obj_ref_3393_inst_req_0 : boolean;
  signal simple_obj_ref_3440_inst_ack_0 : boolean;
  signal simple_obj_ref_3433_inst_req_0 : boolean;
  signal simple_obj_ref_3436_inst_req_0 : boolean;
  signal binary_3356_inst_req_0 : boolean;
  signal array_obj_ref_3390_final_reg_ack_0 : boolean;
  signal array_obj_ref_3390_final_reg_req_0 : boolean;
  signal array_obj_ref_3462_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3462_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_3462_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3462_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3462_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3462_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_3462_offset_inst_req_0 : boolean;
  signal array_obj_ref_3462_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3462_base_resize_req_0 : boolean;
  signal array_obj_ref_3462_base_resize_ack_0 : boolean;
  signal array_obj_ref_3462_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3462_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3462_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3462_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3462_final_reg_req_0 : boolean;
  signal array_obj_ref_3462_final_reg_ack_0 : boolean;
  signal simple_obj_ref_3460_inst_req_0 : boolean;
  signal simple_obj_ref_3460_inst_ack_0 : boolean;
  signal simple_obj_ref_3465_inst_req_0 : boolean;
  signal simple_obj_ref_3465_inst_ack_0 : boolean;
  signal binary_3470_inst_req_0 : boolean;
  signal binary_3470_inst_ack_0 : boolean;
  signal binary_3470_inst_req_1 : boolean;
  signal binary_3470_inst_ack_1 : boolean;
  signal binary_3476_inst_req_0 : boolean;
  signal binary_3476_inst_ack_0 : boolean;
  signal binary_3476_inst_req_1 : boolean;
  signal binary_3476_inst_ack_1 : boolean;
  signal ternary_3479_inst_req_0 : boolean;
  signal ternary_3479_inst_ack_0 : boolean;
  signal simple_obj_ref_3473_inst_req_0 : boolean;
  signal simple_obj_ref_3473_inst_ack_0 : boolean;
  signal binary_3484_inst_req_0 : boolean;
  signal binary_3484_inst_ack_0 : boolean;
  signal binary_3484_inst_req_1 : boolean;
  signal binary_3484_inst_ack_1 : boolean;
  signal if_stmt_3481_branch_req_0 : boolean;
  signal if_stmt_3481_branch_ack_1 : boolean;
  signal if_stmt_3481_branch_ack_0 : boolean;
  signal phi_stmt_3450_req_0 : boolean;
  signal phi_stmt_3450_req_1 : boolean;
  signal phi_stmt_3450_ack_0 : boolean;
  signal simple_obj_ref_3493_inst_req_0 : boolean;
  signal simple_obj_ref_3493_inst_ack_0 : boolean;
  signal simple_obj_ref_3491_inst_req_0 : boolean;
  signal simple_obj_ref_3491_inst_ack_0 : boolean;
  signal ptr_deref_3492_base_resize_req_0 : boolean;
  signal ptr_deref_3492_base_resize_ack_0 : boolean;
  signal ptr_deref_3492_root_address_inst_req_0 : boolean;
  signal ptr_deref_3492_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3492_addr_0_req_0 : boolean;
  signal ptr_deref_3492_addr_0_ack_0 : boolean;
  signal ptr_deref_3492_addr_0_req_1 : boolean;
  signal ptr_deref_3492_addr_0_ack_1 : boolean;
  signal ptr_deref_3492_addr_1_req_0 : boolean;
  signal ptr_deref_3492_addr_1_ack_0 : boolean;
  signal ptr_deref_3492_addr_1_req_1 : boolean;
  signal ptr_deref_3492_addr_1_ack_1 : boolean;
  signal ptr_deref_3492_addr_2_req_0 : boolean;
  signal ptr_deref_3492_addr_2_ack_0 : boolean;
  signal ptr_deref_3492_addr_2_req_1 : boolean;
  signal ptr_deref_3492_addr_2_ack_1 : boolean;
  signal ptr_deref_3492_addr_3_req_0 : boolean;
  signal ptr_deref_3492_addr_3_ack_0 : boolean;
  signal ptr_deref_3492_addr_3_req_1 : boolean;
  signal ptr_deref_3492_addr_3_ack_1 : boolean;
  signal ptr_deref_3492_addr_4_req_0 : boolean;
  signal ptr_deref_3492_addr_4_ack_0 : boolean;
  signal ptr_deref_3492_addr_4_req_1 : boolean;
  signal ptr_deref_3492_addr_4_ack_1 : boolean;
  signal ptr_deref_3492_addr_5_req_0 : boolean;
  signal ptr_deref_3492_addr_5_ack_0 : boolean;
  signal ptr_deref_3492_addr_5_req_1 : boolean;
  signal ptr_deref_3492_addr_5_ack_1 : boolean;
  signal ptr_deref_3492_addr_6_req_0 : boolean;
  signal ptr_deref_3492_addr_6_ack_0 : boolean;
  signal ptr_deref_3492_addr_6_req_1 : boolean;
  signal ptr_deref_3492_addr_6_ack_1 : boolean;
  signal ptr_deref_3492_addr_7_req_0 : boolean;
  signal ptr_deref_3492_addr_7_ack_0 : boolean;
  signal ptr_deref_3492_addr_7_req_1 : boolean;
  signal ptr_deref_3492_addr_7_ack_1 : boolean;
  signal ptr_deref_3492_gather_scatter_req_0 : boolean;
  signal ptr_deref_3492_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3492_store_0_req_0 : boolean;
  signal ptr_deref_3492_store_0_ack_0 : boolean;
  signal ptr_deref_3492_store_1_req_0 : boolean;
  signal ptr_deref_3492_store_1_ack_0 : boolean;
  signal ptr_deref_3492_store_2_req_0 : boolean;
  signal ptr_deref_3492_store_2_ack_0 : boolean;
  signal ptr_deref_3492_store_3_req_0 : boolean;
  signal ptr_deref_3492_store_3_ack_0 : boolean;
  signal ptr_deref_3492_store_4_req_0 : boolean;
  signal ptr_deref_3492_store_4_ack_0 : boolean;
  signal ptr_deref_3492_store_5_req_0 : boolean;
  signal ptr_deref_3492_store_5_ack_0 : boolean;
  signal ptr_deref_3492_store_6_req_0 : boolean;
  signal ptr_deref_3492_store_6_ack_0 : boolean;
  signal ptr_deref_3492_store_7_req_0 : boolean;
  signal ptr_deref_3492_store_7_ack_0 : boolean;
  signal ptr_deref_3492_store_0_req_1 : boolean;
  signal ptr_deref_3492_store_0_ack_1 : boolean;
  signal ptr_deref_3492_store_1_req_1 : boolean;
  signal ptr_deref_3492_store_1_ack_1 : boolean;
  signal ptr_deref_3492_store_2_req_1 : boolean;
  signal ptr_deref_3492_store_2_ack_1 : boolean;
  signal ptr_deref_3492_store_3_req_1 : boolean;
  signal ptr_deref_3492_store_3_ack_1 : boolean;
  signal ptr_deref_3492_store_4_req_1 : boolean;
  signal ptr_deref_3492_store_4_ack_1 : boolean;
  signal ptr_deref_3492_store_5_req_1 : boolean;
  signal ptr_deref_3492_store_5_ack_1 : boolean;
  signal ptr_deref_3492_store_6_req_1 : boolean;
  signal ptr_deref_3492_store_6_ack_1 : boolean;
  signal ptr_deref_3492_store_7_req_1 : boolean;
  signal ptr_deref_3492_store_7_ack_1 : boolean;
  signal simple_obj_ref_3496_inst_req_0 : boolean;
  signal simple_obj_ref_3496_inst_ack_0 : boolean;
  signal binary_3498_inst_req_0 : boolean;
  signal binary_3498_inst_ack_0 : boolean;
  signal binary_3498_inst_req_1 : boolean;
  signal binary_3498_inst_ack_1 : boolean;
  signal if_stmt_3495_branch_req_0 : boolean;
  signal if_stmt_3495_branch_ack_1 : boolean;
  signal if_stmt_3495_branch_ack_0 : boolean;
  signal simple_obj_ref_3500_inst_req_0 : boolean;
  signal simple_obj_ref_3500_inst_ack_0 : boolean;
  signal type_cast_3501_inst_req_0 : boolean;
  signal type_cast_3501_inst_ack_0 : boolean;
  signal simple_obj_ref_3499_inst_req_0 : boolean;
  signal simple_obj_ref_3499_inst_ack_0 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  receive_packet_pipeline_CP_16919: Block -- control-path 
    signal cp_elements: BooleanArray(353 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(353);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(353), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cp_elements(2) <= false; 
    cp_elements(3) <= OrReduce(cp_elements(97) & cp_elements(100));
    req_16946_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_3330_inst_req_0); -- 
    ack_16947_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3330_inst_ack_0, ack => cp_elements(4)); -- 
    cp_elements(5) <= cp_elements(4);
    cpelement_group_6 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(7) & cp_elements(47) & cp_elements(91));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(6),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17139_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(6), ack => binary_3369_inst_req_0); -- 
    cp_elements(7) <= cp_elements(5);
    cpelement_group_8 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(9) & cp_elements(25) & cp_elements(45));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(8),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => binary_3349_inst_req_0); -- 
    cp_elements(9) <= cp_elements(5);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(11) & cp_elements(15) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16987_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => binary_3339_inst_req_0); -- 
    cp_elements(11) <= cp_elements(5);
    cpelement_group_12 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(13) & cp_elements(14));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(12),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16965_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => type_cast_3334_inst_req_0); -- 
    cp_elements(13) <= cp_elements(5);
    cp_elements(14) <= cp_elements(5);
    ack_16966_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3334_inst_ack_0, ack => cp_elements(15)); -- 
    cpelement_group_16 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(17) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(16),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_16982_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => type_cast_3338_inst_req_0); -- 
    cp_elements(17) <= cp_elements(5);
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(20));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_16975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => binary_3337_inst_req_0); -- 
    cp_elements(19) <= cp_elements(5);
    cp_elements(20) <= cp_elements(5);
    ra_16976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3337_inst_ack_0, ack => cp_elements(21)); -- 
    cr_16977_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => binary_3337_inst_req_1); -- 
    ca_16978_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3337_inst_ack_1, ack => cp_elements(22)); -- 
    ack_16983_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3338_inst_ack_0, ack => cp_elements(23)); -- 
    ra_16988_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3339_inst_ack_0, ack => cp_elements(24)); -- 
    cr_16989_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => binary_3339_inst_req_1); -- 
    ca_16990_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3339_inst_ack_1, ack => cp_elements(25)); -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(27) & cp_elements(35) & cp_elements(43));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => binary_3348_inst_req_0); -- 
    cp_elements(27) <= cp_elements(5);
    cpelement_group_28 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(29) & cp_elements(34));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(28),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => type_cast_3343_inst_req_0); -- 
    cp_elements(29) <= cp_elements(5);
    cpelement_group_30 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(31) & cp_elements(32));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(30),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17001_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => binary_3342_inst_req_0); -- 
    cp_elements(31) <= cp_elements(5);
    cp_elements(32) <= cp_elements(5);
    ra_17002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3342_inst_ack_0, ack => cp_elements(33)); -- 
    cr_17003_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => binary_3342_inst_req_1); -- 
    ca_17004_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3342_inst_ack_1, ack => cp_elements(34)); -- 
    ack_17009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3343_inst_ack_0, ack => cp_elements(35)); -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(37) & cp_elements(42));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17025_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => type_cast_3347_inst_req_0); -- 
    cp_elements(37) <= cp_elements(5);
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(39) & cp_elements(40));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => binary_3346_inst_req_0); -- 
    cp_elements(39) <= cp_elements(5);
    cp_elements(40) <= cp_elements(5);
    ra_17019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3346_inst_ack_0, ack => cp_elements(41)); -- 
    cr_17020_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => binary_3346_inst_req_1); -- 
    ca_17021_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3346_inst_ack_1, ack => cp_elements(42)); -- 
    ack_17026_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3347_inst_ack_0, ack => cp_elements(43)); -- 
    ra_17031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3348_inst_ack_0, ack => cp_elements(44)); -- 
    cr_17032_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => binary_3348_inst_req_1); -- 
    ca_17033_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3348_inst_ack_1, ack => cp_elements(45)); -- 
    ra_17038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3349_inst_ack_0, ack => cp_elements(46)); -- 
    cr_17039_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => binary_3349_inst_req_1); -- 
    ca_17040_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3349_inst_ack_1, ack => cp_elements(47)); -- 
    cpelement_group_48 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(49) & cp_elements(69) & cp_elements(89));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(48),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17132_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(48), ack => binary_3368_inst_req_0); -- 
    cp_elements(49) <= cp_elements(5);
    cpelement_group_50 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(51) & cp_elements(59) & cp_elements(67));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(50),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(50), ack => binary_3358_inst_req_0); -- 
    cp_elements(51) <= cp_elements(5);
    cpelement_group_52 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(53) & cp_elements(58));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(52),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => type_cast_3353_inst_req_0); -- 
    cp_elements(53) <= cp_elements(5);
    cpelement_group_54 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(55) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(54),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(54), ack => binary_3352_inst_req_0); -- 
    cp_elements(55) <= cp_elements(5);
    cp_elements(56) <= cp_elements(5);
    ra_17054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3352_inst_ack_0, ack => cp_elements(57)); -- 
    cr_17055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => binary_3352_inst_req_1); -- 
    ca_17056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3352_inst_ack_1, ack => cp_elements(58)); -- 
    ack_17061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3353_inst_ack_0, ack => cp_elements(59)); -- 
    cpelement_group_60 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(66));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(60),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => type_cast_3357_inst_req_0); -- 
    cp_elements(61) <= cp_elements(5);
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(63) & cp_elements(64));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => binary_3356_inst_req_0); -- 
    cp_elements(63) <= cp_elements(5);
    cp_elements(64) <= cp_elements(5);
    ra_17071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3356_inst_ack_0, ack => cp_elements(65)); -- 
    cr_17072_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => binary_3356_inst_req_1); -- 
    ca_17073_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3356_inst_ack_1, ack => cp_elements(66)); -- 
    ack_17078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3357_inst_ack_0, ack => cp_elements(67)); -- 
    ra_17083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3358_inst_ack_0, ack => cp_elements(68)); -- 
    cr_17084_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => binary_3358_inst_req_1); -- 
    ca_17085_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3358_inst_ack_1, ack => cp_elements(69)); -- 
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(71) & cp_elements(79) & cp_elements(87));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => binary_3367_inst_req_0); -- 
    cp_elements(71) <= cp_elements(5);
    cpelement_group_72 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(73) & cp_elements(78));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(72),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17103_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => type_cast_3362_inst_req_0); -- 
    cp_elements(73) <= cp_elements(5);
    cpelement_group_74 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(75) & cp_elements(76));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(74),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => binary_3361_inst_req_0); -- 
    cp_elements(75) <= cp_elements(5);
    cp_elements(76) <= cp_elements(5);
    ra_17097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3361_inst_ack_0, ack => cp_elements(77)); -- 
    cr_17098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => binary_3361_inst_req_1); -- 
    ca_17099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3361_inst_ack_1, ack => cp_elements(78)); -- 
    ack_17104_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3362_inst_ack_0, ack => cp_elements(79)); -- 
    cpelement_group_80 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(81) & cp_elements(86));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(80),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => type_cast_3366_inst_req_0); -- 
    cp_elements(81) <= cp_elements(5);
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17113_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => binary_3365_inst_req_0); -- 
    cp_elements(83) <= cp_elements(5);
    cp_elements(84) <= cp_elements(5);
    ra_17114_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3365_inst_ack_0, ack => cp_elements(85)); -- 
    cr_17115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => binary_3365_inst_req_1); -- 
    ca_17116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3365_inst_ack_1, ack => cp_elements(86)); -- 
    ack_17121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3366_inst_ack_0, ack => cp_elements(87)); -- 
    ra_17126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3367_inst_ack_0, ack => cp_elements(88)); -- 
    cr_17127_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => binary_3367_inst_req_1); -- 
    ca_17128_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3367_inst_ack_1, ack => cp_elements(89)); -- 
    ra_17133_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3368_inst_ack_0, ack => cp_elements(90)); -- 
    cr_17134_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(90), ack => binary_3368_inst_req_1); -- 
    ca_17135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3368_inst_ack_1, ack => cp_elements(91)); -- 
    ra_17140_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3369_inst_ack_0, ack => cp_elements(92)); -- 
    cr_17141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => binary_3369_inst_req_1); -- 
    ca_17142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3369_inst_ack_1, ack => cp_elements(93)); -- 
    pipe_wreq_17147_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => simple_obj_ref_3332_inst_req_0); -- 
    pipe_wack_17148_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3332_inst_ack_0, ack => cp_elements(94)); -- 
    cp_elements(95) <= cp_elements(1);
    cp_elements(96) <= false;
    cp_elements(97) <= cp_elements(96);
    cp_elements(98) <= cp_elements(1);
    cp_elements(99) <= OrReduce(cp_elements(94) & cp_elements(98));
    cp_elements(100) <= cp_elements(99);
    cp_elements(101) <= cp_elements(0);
    cp_elements(102) <= false; 
    cp_elements(103) <= OrReduce(cp_elements(141) & cp_elements(144));
    req_17190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => simple_obj_ref_3377_inst_req_0); -- 
    cp_elements(104) <= cp_elements(122);
    cp_elements(105) <= cp_elements(138);
    ack_17191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3377_inst_ack_0, ack => cp_elements(106)); -- 
    cp_elements(107) <= cp_elements(106);
    cpelement_group_108 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(109) & cp_elements(110));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(108),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => type_cast_3382_inst_req_0); -- 
    cp_elements(109) <= cp_elements(107);
    cp_elements(110) <= cp_elements(107);
    ack_17204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3382_inst_ack_0, ack => cp_elements(111)); -- 
    base_resize_req_17225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => array_obj_ref_3390_base_resize_req_0); -- 
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(113) & cp_elements(114));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => type_cast_3386_inst_req_0); -- 
    cp_elements(113) <= cp_elements(107);
    cp_elements(114) <= cp_elements(107);
    ack_17214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3386_inst_ack_0, ack => cp_elements(115)); -- 
    cp_elements(116) <= cp_elements(107);
    cpelement_group_117 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(116) & cp_elements(120));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_17238_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => array_obj_ref_3390_final_reg_req_0); -- 
    base_resize_ack_17226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3390_base_resize_ack_0, ack => cp_elements(118)); -- 
    plus_base_rr_17231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_3390_root_address_inst_req_0); -- 
    plus_base_ra_17232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3390_root_address_inst_ack_0, ack => cp_elements(119)); -- 
    plus_base_cr_17233_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => array_obj_ref_3390_root_address_inst_req_1); -- 
    plus_base_ca_17234_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3390_root_address_inst_ack_1, ack => cp_elements(120)); -- 
    final_reg_ack_17239_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3390_final_reg_ack_0, ack => cp_elements(121)); -- 
    cpelement_group_122 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(115) & cp_elements(121));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(122),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(123) <= cp_elements(104);
    cp_elements(124) <= cp_elements(123);
    pipe_wreq_17253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => simple_obj_ref_3393_inst_req_0); -- 
    pipe_wack_17254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3393_inst_ack_0, ack => cp_elements(125)); -- 
    cp_elements(126) <= cp_elements(123);
    pipe_wreq_17265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => simple_obj_ref_3396_inst_req_0); -- 
    pipe_wack_17266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3396_inst_ack_0, ack => cp_elements(127)); -- 
    cp_elements(128) <= cp_elements(123);
    pipe_wreq_17277_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => simple_obj_ref_3399_inst_req_0); -- 
    pipe_wack_17278_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3399_inst_ack_0, ack => cp_elements(129)); -- 
    cp_elements(130) <= cp_elements(123);
    cpelement_group_131 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(132) & cp_elements(133));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(131),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17290_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => type_cast_3404_inst_req_0); -- 
    cp_elements(132) <= cp_elements(130);
    cp_elements(133) <= cp_elements(130);
    ack_17291_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3404_inst_ack_0, ack => cp_elements(134)); -- 
    pipe_wreq_17296_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(134), ack => simple_obj_ref_3402_inst_req_0); -- 
    pipe_wack_17297_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3402_inst_ack_0, ack => cp_elements(135)); -- 
    cp_elements(136) <= cp_elements(123);
    pipe_wreq_17308_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => simple_obj_ref_3406_inst_req_0); -- 
    pipe_wack_17309_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3406_inst_ack_0, ack => cp_elements(137)); -- 
    cpelement_group_138 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(125) & cp_elements(127) & cp_elements(129) & cp_elements(135) & cp_elements(137));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(138),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(139) <= cp_elements(101);
    cp_elements(140) <= false;
    cp_elements(141) <= cp_elements(140);
    cp_elements(142) <= cp_elements(101);
    cp_elements(143) <= OrReduce(cp_elements(105) & cp_elements(142));
    cp_elements(144) <= cp_elements(143);
    cp_elements(145) <= cp_elements(0);
    cp_elements(146) <= false; 
    cp_elements(147) <= OrReduce(cp_elements(238) & cp_elements(241));
    cp_elements(148) <= cp_elements(164);
    cp_elements(149) <= OrReduce(cp_elements(244) & cp_elements(247));
    cp_elements(150) <= cp_elements(175);
    cp_elements(151) <= OrReduce(cp_elements(178) & cp_elements(186));
    cp_elements(152) <= OrReduce(cp_elements(250) & cp_elements(254));
    cp_elements(153) <= cp_elements(214);
    cp_elements(154) <= OrReduce(cp_elements(227) & cp_elements(235));
    cp_elements(155) <= cp_elements(147);
    cp_elements(156) <= cp_elements(155);
    req_17361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => simple_obj_ref_3416_inst_req_0); -- 
    ack_17362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3416_inst_ack_0, ack => cp_elements(157)); -- 
    cp_elements(158) <= cp_elements(155);
    req_17372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => simple_obj_ref_3419_inst_req_0); -- 
    ack_17373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3419_inst_ack_0, ack => cp_elements(159)); -- 
    cp_elements(160) <= cp_elements(155);
    req_17383_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => simple_obj_ref_3422_inst_req_0); -- 
    ack_17384_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3422_inst_ack_0, ack => cp_elements(161)); -- 
    cp_elements(162) <= cp_elements(155);
    req_17394_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => simple_obj_ref_3425_inst_req_0); -- 
    ack_17395_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3425_inst_ack_0, ack => cp_elements(163)); -- 
    cpelement_group_164 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(157) & cp_elements(159) & cp_elements(161) & cp_elements(163));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(164),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(165) <= cp_elements(149);
    cp_elements(166) <= cp_elements(165);
    req_17408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(166), ack => simple_obj_ref_3431_inst_req_0); -- 
    ack_17409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3431_inst_ack_0, ack => cp_elements(167)); -- 
    pipe_wreq_17414_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(167), ack => simple_obj_ref_3430_inst_req_0); -- 
    pipe_wack_17415_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3430_inst_ack_0, ack => cp_elements(168)); -- 
    cp_elements(169) <= cp_elements(165);
    pipe_wreq_17425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(169), ack => simple_obj_ref_3433_inst_req_0); -- 
    pipe_wack_17426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3433_inst_ack_0, ack => cp_elements(170)); -- 
    cp_elements(171) <= cp_elements(165);
    pipe_wreq_17437_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => simple_obj_ref_3436_inst_req_0); -- 
    pipe_wack_17438_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3436_inst_ack_0, ack => cp_elements(172)); -- 
    cp_elements(173) <= cp_elements(165);
    req_17448_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => simple_obj_ref_3440_inst_req_0); -- 
    ack_17449_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3440_inst_ack_0, ack => cp_elements(174)); -- 
    cpelement_group_175 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(168) & cp_elements(170) & cp_elements(172) & cp_elements(174));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(176) <= cp_elements(150);
    cp_elements(177) <= false;
    cp_elements(178) <= cp_elements(177);
    cp_elements(179) <= cp_elements(150);
    rr_17463_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(179), ack => binary_3446_inst_req_0); -- 
    ra_17464_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3446_inst_ack_0, ack => cp_elements(180)); -- 
    cr_17465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(180), ack => binary_3446_inst_req_1); -- 
    ca_17466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3446_inst_ack_1, ack => cp_elements(181)); -- 
    branch_req_17467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(181), ack => if_stmt_3443_branch_req_0); -- 
    cp_elements(182) <= cp_elements(181);
    cp_elements(183) <= cp_elements(182);
    if_choice_transition_17472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3443_branch_ack_1, ack => cp_elements(184)); -- 
    cp_elements(185) <= cp_elements(182);
    else_choice_transition_17476_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3443_branch_ack_0, ack => cp_elements(186)); -- 
    cp_elements(187) <= cp_elements(152);
    cp_elements(188) <= cp_elements(187);
    req_17490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => simple_obj_ref_3458_inst_req_0); -- 
    ack_17491_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3458_inst_ack_0, ack => cp_elements(189)); -- 
    pipe_wreq_17496_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => simple_obj_ref_3457_inst_req_0); -- 
    pipe_wack_17497_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3457_inst_ack_0, ack => cp_elements(190)); -- 
    cp_elements(191) <= cp_elements(187);
    cp_elements(192) <= cp_elements(191);
    cpelement_group_193 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(192) & cp_elements(203));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(193),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_17546_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => array_obj_ref_3462_final_reg_req_0); -- 
    cp_elements(194) <= cp_elements(191);
    base_resize_req_17533_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => array_obj_ref_3462_base_resize_req_0); -- 
    cp_elements(195) <= cp_elements(191);
    index_resize_req_17515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(195), ack => array_obj_ref_3462_index_0_resize_req_0); -- 
    index_resize_ack_17516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_index_0_resize_ack_0, ack => cp_elements(196)); -- 
    scale_rr_17520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => array_obj_ref_3462_index_0_scale_req_0); -- 
    scale_ra_17521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_index_0_scale_ack_0, ack => cp_elements(197)); -- 
    scale_cr_17522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => array_obj_ref_3462_index_0_scale_req_1); -- 
    scale_ca_17523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_index_0_scale_ack_1, ack => cp_elements(198)); -- 
    final_index_req_17527_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(198), ack => array_obj_ref_3462_offset_inst_req_0); -- 
    final_index_ack_17528_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_offset_inst_ack_0, ack => cp_elements(199)); -- 
    base_resize_ack_17534_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_base_resize_ack_0, ack => cp_elements(200)); -- 
    cpelement_group_201 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(199) & cp_elements(200));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(201),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_17539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => array_obj_ref_3462_root_address_inst_req_0); -- 
    plus_base_ra_17540_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_root_address_inst_ack_0, ack => cp_elements(202)); -- 
    plus_base_cr_17541_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(202), ack => array_obj_ref_3462_root_address_inst_req_1); -- 
    plus_base_ca_17542_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_root_address_inst_ack_1, ack => cp_elements(203)); -- 
    final_reg_ack_17547_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3462_final_reg_ack_0, ack => cp_elements(204)); -- 
    pipe_wreq_17552_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(204), ack => simple_obj_ref_3460_inst_req_0); -- 
    pipe_wack_17553_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3460_inst_ack_0, ack => cp_elements(205)); -- 
    cp_elements(206) <= cp_elements(187);
    req_17563_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => simple_obj_ref_3465_inst_req_0); -- 
    ack_17564_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3465_inst_ack_0, ack => cp_elements(207)); -- 
    cp_elements(208) <= cp_elements(187);
    cpelement_group_209 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(210) & cp_elements(211));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(209),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => binary_3470_inst_req_0); -- 
    cp_elements(210) <= cp_elements(208);
    cp_elements(211) <= cp_elements(208);
    ra_17577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3470_inst_ack_0, ack => cp_elements(212)); -- 
    cr_17578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => binary_3470_inst_req_1); -- 
    ca_17579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3470_inst_ack_1, ack => cp_elements(213)); -- 
    cpelement_group_214 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(190) & cp_elements(205) & cp_elements(207) & cp_elements(213));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(214),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(215) <= cp_elements(153);
    cp_elements(216) <= cp_elements(215);
    cpelement_group_217 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(216) & cp_elements(222));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(217),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ternary_3479_inst_req_0); -- 
    cpelement_group_218 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(219) & cp_elements(220));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(218),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_17593_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(218), ack => binary_3476_inst_req_0); -- 
    cp_elements(219) <= cp_elements(215);
    cp_elements(220) <= cp_elements(215);
    ra_17594_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3476_inst_ack_0, ack => cp_elements(221)); -- 
    cr_17595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => binary_3476_inst_req_1); -- 
    ca_17596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3476_inst_ack_1, ack => cp_elements(222)); -- 
    ack_17601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ternary_3479_inst_ack_0, ack => cp_elements(223)); -- 
    pipe_wreq_17606_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => simple_obj_ref_3473_inst_req_0); -- 
    pipe_wack_17607_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3473_inst_ack_0, ack => cp_elements(224)); -- 
    cp_elements(225) <= cp_elements(224);
    cp_elements(226) <= false;
    cp_elements(227) <= cp_elements(226);
    cp_elements(228) <= cp_elements(224);
    rr_17621_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(228), ack => binary_3484_inst_req_0); -- 
    ra_17622_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3484_inst_ack_0, ack => cp_elements(229)); -- 
    cr_17623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => binary_3484_inst_req_1); -- 
    ca_17624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3484_inst_ack_1, ack => cp_elements(230)); -- 
    branch_req_17625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(230), ack => if_stmt_3481_branch_req_0); -- 
    cp_elements(231) <= cp_elements(230);
    cp_elements(232) <= cp_elements(231);
    if_choice_transition_17630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3481_branch_ack_1, ack => cp_elements(233)); -- 
    phi_stmt_3450_req_17689_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(233), ack => phi_stmt_3450_req_1); -- 
    cp_elements(234) <= cp_elements(231);
    else_choice_transition_17634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3481_branch_ack_0, ack => cp_elements(235)); -- 
    cp_elements(236) <= cp_elements(145);
    cp_elements(237) <= false;
    cp_elements(238) <= cp_elements(237);
    cp_elements(239) <= cp_elements(145);
    cp_elements(240) <= OrReduce(cp_elements(154) & cp_elements(239));
    cp_elements(241) <= cp_elements(240);
    cp_elements(242) <= cp_elements(148);
    cp_elements(243) <= false;
    cp_elements(244) <= cp_elements(243);
    cp_elements(245) <= cp_elements(148);
    cp_elements(246) <= OrReduce(cp_elements(184) & cp_elements(245));
    cp_elements(247) <= cp_elements(246);
    cp_elements(248) <= cp_elements(151);
    cp_elements(249) <= false;
    cp_elements(250) <= cp_elements(249);
    cp_elements(251) <= cp_elements(151);
    phi_stmt_3450_req_17679_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => phi_stmt_3450_req_0); -- 
    cp_elements(252) <= OrReduce(cp_elements(233) & cp_elements(251));
    cp_elements(253) <= cp_elements(252);
    phi_stmt_3450_ack_17694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3450_ack_0, ack => cp_elements(254)); -- 
    cp_elements(255) <= cp_elements(0);
    cp_elements(256) <= false; 
    cp_elements(257) <= OrReduce(cp_elements(349) & cp_elements(352));
    cp_elements(258) <= OrReduce(cp_elements(330) & cp_elements(339) & cp_elements(346));
    cp_elements(259) <= cp_elements(257);
    cp_elements(260) <= cp_elements(259);
    req_17716_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(260), ack => simple_obj_ref_3493_inst_req_0); -- 
    ack_17717_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3493_inst_ack_0, ack => cp_elements(261)); -- 
    cpelement_group_262 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(261) & cp_elements(264) & cp_elements(292));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(262),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_17802_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(262), ack => ptr_deref_3492_gather_scatter_req_0); -- 
    cp_elements(263) <= cp_elements(259);
    req_17725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(263), ack => simple_obj_ref_3491_inst_req_0); -- 
    cp_elements(264) <= simple_obj_ref_3491_inst_ack_0;
    cp_elements(265) <= cp_elements(264);
    base_resize_req_17733_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(265), ack => ptr_deref_3492_base_resize_req_0); -- 
    base_resize_ack_17734_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_base_resize_ack_0, ack => cp_elements(266)); -- 
    sum_rename_req_17738_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => ptr_deref_3492_root_address_inst_req_0); -- 
    cp_elements(267) <= ptr_deref_3492_root_address_inst_ack_0;
    cp_elements(268) <= cp_elements(267);
    rr_17746_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => ptr_deref_3492_addr_0_req_0); -- 
    ra_17747_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_0_ack_0, ack => cp_elements(269)); -- 
    cr_17748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(269), ack => ptr_deref_3492_addr_0_req_1); -- 
    ca_17749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_0_ack_1, ack => cp_elements(270)); -- 
    cp_elements(271) <= cp_elements(267);
    rr_17753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => ptr_deref_3492_addr_1_req_0); -- 
    ra_17754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_1_ack_0, ack => cp_elements(272)); -- 
    cr_17755_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(272), ack => ptr_deref_3492_addr_1_req_1); -- 
    ca_17756_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_1_ack_1, ack => cp_elements(273)); -- 
    cp_elements(274) <= cp_elements(267);
    rr_17760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => ptr_deref_3492_addr_2_req_0); -- 
    ra_17761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_2_ack_0, ack => cp_elements(275)); -- 
    cr_17762_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => ptr_deref_3492_addr_2_req_1); -- 
    ca_17763_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_2_ack_1, ack => cp_elements(276)); -- 
    cp_elements(277) <= cp_elements(267);
    rr_17767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => ptr_deref_3492_addr_3_req_0); -- 
    ra_17768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_3_ack_0, ack => cp_elements(278)); -- 
    cr_17769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(278), ack => ptr_deref_3492_addr_3_req_1); -- 
    ca_17770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_3_ack_1, ack => cp_elements(279)); -- 
    cp_elements(280) <= cp_elements(267);
    rr_17774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(280), ack => ptr_deref_3492_addr_4_req_0); -- 
    ra_17775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_4_ack_0, ack => cp_elements(281)); -- 
    cr_17776_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => ptr_deref_3492_addr_4_req_1); -- 
    ca_17777_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_4_ack_1, ack => cp_elements(282)); -- 
    cp_elements(283) <= cp_elements(267);
    rr_17781_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => ptr_deref_3492_addr_5_req_0); -- 
    ra_17782_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_5_ack_0, ack => cp_elements(284)); -- 
    cr_17783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => ptr_deref_3492_addr_5_req_1); -- 
    ca_17784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_5_ack_1, ack => cp_elements(285)); -- 
    cp_elements(286) <= cp_elements(267);
    rr_17788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => ptr_deref_3492_addr_6_req_0); -- 
    ra_17789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_6_ack_0, ack => cp_elements(287)); -- 
    cr_17790_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(287), ack => ptr_deref_3492_addr_6_req_1); -- 
    ca_17791_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_6_ack_1, ack => cp_elements(288)); -- 
    cp_elements(289) <= cp_elements(267);
    rr_17795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => ptr_deref_3492_addr_7_req_0); -- 
    ra_17796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_7_ack_0, ack => cp_elements(290)); -- 
    cr_17797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => ptr_deref_3492_addr_7_req_1); -- 
    ca_17798_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_addr_7_ack_1, ack => cp_elements(291)); -- 
    cpelement_group_292 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(270) & cp_elements(273) & cp_elements(276) & cp_elements(279) & cp_elements(282) & cp_elements(285) & cp_elements(288) & cp_elements(291));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(292),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(293) <= ptr_deref_3492_gather_scatter_ack_0;
    cp_elements(294) <= cp_elements(293);
    rr_17810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(294), ack => ptr_deref_3492_store_0_req_0); -- 
    ra_17811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_0_ack_0, ack => cp_elements(295)); -- 
    cp_elements(296) <= cp_elements(293);
    rr_17815_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(296), ack => ptr_deref_3492_store_1_req_0); -- 
    ra_17816_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_1_ack_0, ack => cp_elements(297)); -- 
    cp_elements(298) <= cp_elements(293);
    rr_17820_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => ptr_deref_3492_store_2_req_0); -- 
    ra_17821_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_2_ack_0, ack => cp_elements(299)); -- 
    cp_elements(300) <= cp_elements(293);
    rr_17825_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(300), ack => ptr_deref_3492_store_3_req_0); -- 
    ra_17826_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_3_ack_0, ack => cp_elements(301)); -- 
    cp_elements(302) <= cp_elements(293);
    rr_17830_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(302), ack => ptr_deref_3492_store_4_req_0); -- 
    ra_17831_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_4_ack_0, ack => cp_elements(303)); -- 
    cp_elements(304) <= cp_elements(293);
    rr_17835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(304), ack => ptr_deref_3492_store_5_req_0); -- 
    ra_17836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_5_ack_0, ack => cp_elements(305)); -- 
    cp_elements(306) <= cp_elements(293);
    rr_17840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => ptr_deref_3492_store_6_req_0); -- 
    ra_17841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_6_ack_0, ack => cp_elements(307)); -- 
    cp_elements(308) <= cp_elements(293);
    rr_17845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(308), ack => ptr_deref_3492_store_7_req_0); -- 
    ra_17846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_7_ack_0, ack => cp_elements(309)); -- 
    cpelement_group_310 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(295) & cp_elements(297) & cp_elements(299) & cp_elements(301) & cp_elements(303) & cp_elements(305) & cp_elements(307) & cp_elements(309));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(310),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(311) <= cp_elements(310);
    cr_17856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => ptr_deref_3492_store_0_req_1); -- 
    ca_17857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_0_ack_1, ack => cp_elements(312)); -- 
    cp_elements(313) <= cp_elements(310);
    cr_17861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => ptr_deref_3492_store_1_req_1); -- 
    ca_17862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_1_ack_1, ack => cp_elements(314)); -- 
    cp_elements(315) <= cp_elements(310);
    cr_17866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => ptr_deref_3492_store_2_req_1); -- 
    ca_17867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_2_ack_1, ack => cp_elements(316)); -- 
    cp_elements(317) <= cp_elements(310);
    cr_17871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(317), ack => ptr_deref_3492_store_3_req_1); -- 
    ca_17872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_3_ack_1, ack => cp_elements(318)); -- 
    cp_elements(319) <= cp_elements(310);
    cr_17876_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => ptr_deref_3492_store_4_req_1); -- 
    ca_17877_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_4_ack_1, ack => cp_elements(320)); -- 
    cp_elements(321) <= cp_elements(310);
    cr_17881_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => ptr_deref_3492_store_5_req_1); -- 
    ca_17882_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_5_ack_1, ack => cp_elements(322)); -- 
    cp_elements(323) <= cp_elements(310);
    cr_17886_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(323), ack => ptr_deref_3492_store_6_req_1); -- 
    ca_17887_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_6_ack_1, ack => cp_elements(324)); -- 
    cp_elements(325) <= cp_elements(310);
    cr_17891_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => ptr_deref_3492_store_7_req_1); -- 
    ca_17892_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3492_store_7_ack_1, ack => cp_elements(326)); -- 
    cpelement_group_327 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(312) & cp_elements(314) & cp_elements(316) & cp_elements(318) & cp_elements(320) & cp_elements(322) & cp_elements(324) & cp_elements(326));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(327),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(328) <= cp_elements(327);
    cp_elements(329) <= false;
    cp_elements(330) <= cp_elements(329);
    cp_elements(331) <= cp_elements(327);
    req_17909_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => simple_obj_ref_3496_inst_req_0); -- 
    ack_17910_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3496_inst_ack_0, ack => cp_elements(332)); -- 
    rr_17911_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(332), ack => binary_3498_inst_req_0); -- 
    ra_17912_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3498_inst_ack_0, ack => cp_elements(333)); -- 
    cr_17913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => binary_3498_inst_req_1); -- 
    ca_17914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3498_inst_ack_1, ack => cp_elements(334)); -- 
    branch_req_17915_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(334), ack => if_stmt_3495_branch_req_0); -- 
    cp_elements(335) <= cp_elements(334);
    cp_elements(336) <= cp_elements(335);
    if_choice_transition_17920_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3495_branch_ack_1, ack => cp_elements(337)); -- 
    cp_elements(338) <= cp_elements(335);
    else_choice_transition_17924_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3495_branch_ack_0, ack => cp_elements(339)); -- 
    cp_elements(340) <= cp_elements(337);
    cpelement_group_341 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(342) & cp_elements(344));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(341),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_17943_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(341), ack => type_cast_3501_inst_req_0); -- 
    cp_elements(342) <= cp_elements(340);
    cp_elements(343) <= cp_elements(340);
    req_17938_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(343), ack => simple_obj_ref_3500_inst_req_0); -- 
    ack_17939_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3500_inst_ack_0, ack => cp_elements(344)); -- 
    ack_17944_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3501_inst_ack_0, ack => cp_elements(345)); -- 
    pipe_wreq_17949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => simple_obj_ref_3499_inst_req_0); -- 
    pipe_wack_17950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3499_inst_ack_0, ack => cp_elements(346)); -- 
    cp_elements(347) <= cp_elements(255);
    cp_elements(348) <= false;
    cp_elements(349) <= cp_elements(348);
    cp_elements(350) <= cp_elements(255);
    cp_elements(351) <= OrReduce(cp_elements(258) & cp_elements(350));
    cp_elements(352) <= cp_elements(351);
    cpelement_group_353 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(102) & cp_elements(146) & cp_elements(256));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(353),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_3450 : std_logic_vector(7 downto 0);
    signal NI_3471 : std_logic_vector(7 downto 0);
    signal a_3331 : std_logic_vector(63 downto 0);
    signal array_obj_ref_3390_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3390_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3390_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3462_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3462_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3462_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3462_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3462_wire : std_logic_vector(31 downto 0);
    signal binary_3337_wire : std_logic_vector(63 downto 0);
    signal binary_3339_wire : std_logic_vector(15 downto 0);
    signal binary_3342_wire : std_logic_vector(63 downto 0);
    signal binary_3346_wire : std_logic_vector(63 downto 0);
    signal binary_3348_wire : std_logic_vector(15 downto 0);
    signal binary_3349_wire : std_logic_vector(31 downto 0);
    signal binary_3352_wire : std_logic_vector(63 downto 0);
    signal binary_3356_wire : std_logic_vector(63 downto 0);
    signal binary_3358_wire : std_logic_vector(15 downto 0);
    signal binary_3361_wire : std_logic_vector(63 downto 0);
    signal binary_3365_wire : std_logic_vector(63 downto 0);
    signal binary_3367_wire : std_logic_vector(15 downto 0);
    signal binary_3368_wire : std_logic_vector(31 downto 0);
    signal binary_3369_wire : std_logic_vector(63 downto 0);
    signal binary_3446_wire : std_logic_vector(0 downto 0);
    signal binary_3476_wire : std_logic_vector(0 downto 0);
    signal binary_3484_wire : std_logic_vector(0 downto 0);
    signal binary_3498_wire : std_logic_vector(0 downto 0);
    signal buf64_ptr_3387 : std_logic_vector(31 downto 0);
    signal buf64_ptr_3420 : std_logic_vector(31 downto 0);
    signal buf8_ptr_3383 : std_logic_vector(31 downto 0);
    signal buf8_ptr_3417 : std_logic_vector(31 downto 0);
    signal buf_3378 : std_logic_vector(31 downto 0);
    signal expr_3336_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3341_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3345_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3351_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3355_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3360_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3364_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3434_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3445_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3469_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3475_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3477_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3478_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3483_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3497_wire_constant : std_logic_vector(0 downto 0);
    signal hdr_in_ctrl_3441 : std_logic_vector(7 downto 0);
    signal pkt64_ptr_3426 : std_logic_vector(31 downto 0);
    signal pkt8_ptr_3391 : std_logic_vector(31 downto 0);
    signal pkt8_ptr_3423 : std_logic_vector(31 downto 0);
    signal pkt_in_ctrl_3466 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_4 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_5 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_6 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_data_7 : std_logic_vector(7 downto 0);
    signal ptr_deref_3492_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3492_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_address_7 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3492_word_offset_7 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3431_wire : std_logic_vector(63 downto 0);
    signal simple_obj_ref_3458_wire : std_logic_vector(63 downto 0);
    signal simple_obj_ref_3461_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3461_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3491_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_3493_wire : std_logic_vector(63 downto 0);
    signal simple_obj_ref_3496_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3500_wire : std_logic_vector(31 downto 0);
    signal ternary_3479_wire : std_logic_vector(0 downto 0);
    signal type_cast_3334_wire : std_logic_vector(7 downto 0);
    signal type_cast_3338_wire : std_logic_vector(7 downto 0);
    signal type_cast_3343_wire : std_logic_vector(7 downto 0);
    signal type_cast_3347_wire : std_logic_vector(7 downto 0);
    signal type_cast_3353_wire : std_logic_vector(7 downto 0);
    signal type_cast_3357_wire : std_logic_vector(7 downto 0);
    signal type_cast_3362_wire : std_logic_vector(7 downto 0);
    signal type_cast_3366_wire : std_logic_vector(7 downto 0);
    signal type_cast_3404_wire : std_logic_vector(31 downto 0);
    signal type_cast_3453_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3501_wire : std_logic_vector(31 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxbuf64_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxbuf64_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxbuf8_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxbuf8_ptr_pipe
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxpkt64_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxpkt64_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxpkt8_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxpkt8_ptr_pipe
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data_last_word_flag
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data_last_word_flag
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxreceive_packet_pipelinexxwrite_data_wptr
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxreceive_packet_pipelinexxwrite_data_wptr
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_3390_final_offset <= "0000000010110100";
    array_obj_ref_3462_offset_scale_factor_0 <= "0000000000001000";
    expr_3336_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    expr_3341_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    expr_3345_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    expr_3351_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    expr_3355_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    expr_3360_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    expr_3364_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    expr_3434_wire_constant <= "0";
    expr_3445_wire_constant <= "11111111";
    expr_3469_wire_constant <= "00000001";
    expr_3475_wire_constant <= "00000000";
    expr_3477_wire_constant <= "0";
    expr_3478_wire_constant <= "1";
    expr_3483_wire_constant <= "00000000";
    expr_3497_wire_constant <= "0";
    ptr_deref_3492_word_offset_0 <= "0000000000000000";
    ptr_deref_3492_word_offset_1 <= "0000000000000001";
    ptr_deref_3492_word_offset_2 <= "0000000000000010";
    ptr_deref_3492_word_offset_3 <= "0000000000000011";
    ptr_deref_3492_word_offset_4 <= "0000000000000100";
    ptr_deref_3492_word_offset_5 <= "0000000000000101";
    ptr_deref_3492_word_offset_6 <= "0000000000000110";
    ptr_deref_3492_word_offset_7 <= "0000000000000111";
    type_cast_3453_wire_constant <= "00000000";
    phi_stmt_3450: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3453_wire_constant & NI_3471;
      req <= phi_stmt_3450_req_0 & phi_stmt_3450_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3450_ack_0,
          idata => idata,
          odata => I_3450,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3450
    ternary_3479_inst: SelectBase generic map(data_width => 1) -- 
      port map( x => expr_3477_wire_constant, y => expr_3478_wire_constant, sel => binary_3476_wire, z => ternary_3479_wire, req => ternary_3479_inst_req_0, ack => ternary_3479_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3390_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => buf8_ptr_3383, dout => array_obj_ref_3390_resized_base_address, req => array_obj_ref_3390_base_resize_req_0, ack => array_obj_ref_3390_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3390_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3390_root_address, dout => pkt8_ptr_3391, req => array_obj_ref_3390_final_reg_req_0, ack => array_obj_ref_3390_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3462_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_ptr_3426, dout => array_obj_ref_3462_resized_base_address, req => array_obj_ref_3462_base_resize_req_0, ack => array_obj_ref_3462_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3462_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3462_root_address, dout => array_obj_ref_3462_wire, req => array_obj_ref_3462_final_reg_req_0, ack => array_obj_ref_3462_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3462_index_0_resize: RegisterBase --
      generic map(in_data_width => 8,out_data_width => 16, flow_through => true ) 
      port map( din => I_3450, dout => simple_obj_ref_3461_resized, req => array_obj_ref_3462_index_0_resize_req_0, ack => array_obj_ref_3462_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3462_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3461_scaled, dout => array_obj_ref_3462_final_offset, req => array_obj_ref_3462_offset_inst_req_0, ack => array_obj_ref_3462_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3492_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3491_wire, dout => ptr_deref_3492_resized_base_address, req => ptr_deref_3492_base_resize_req_0, ack => ptr_deref_3492_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_3334_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => a_3331, dout => type_cast_3334_wire, req => type_cast_3334_inst_req_0, ack => type_cast_3334_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3338_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3337_wire, dout => type_cast_3338_wire, req => type_cast_3338_inst_req_0, ack => type_cast_3338_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3343_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3342_wire, dout => type_cast_3343_wire, req => type_cast_3343_inst_req_0, ack => type_cast_3343_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3347_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3346_wire, dout => type_cast_3347_wire, req => type_cast_3347_inst_req_0, ack => type_cast_3347_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3353_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3352_wire, dout => type_cast_3353_wire, req => type_cast_3353_inst_req_0, ack => type_cast_3353_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3357_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3356_wire, dout => type_cast_3357_wire, req => type_cast_3357_inst_req_0, ack => type_cast_3357_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3362_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3361_wire, dout => type_cast_3362_wire, req => type_cast_3362_inst_req_0, ack => type_cast_3362_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3366_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3365_wire, dout => type_cast_3366_wire, req => type_cast_3366_inst_req_0, ack => type_cast_3366_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3382_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_3378, dout => buf8_ptr_3383, req => type_cast_3382_inst_req_0, ack => type_cast_3382_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3386_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => buf_3378, dout => buf64_ptr_3387, req => type_cast_3386_inst_req_0, ack => type_cast_3386_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3404_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt8_ptr_3391, dout => type_cast_3404_wire, req => type_cast_3404_inst_req_0, ack => type_cast_3404_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3501_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => simple_obj_ref_3500_wire, dout => type_cast_3501_wire, req => type_cast_3501_inst_req_0, ack => type_cast_3501_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3492_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(63 downto 0); --
    begin -- 
      ptr_deref_3492_gather_scatter_ack_0 <= ptr_deref_3492_gather_scatter_req_0;
      aggregated_sig <= simple_obj_ref_3493_wire;
      ptr_deref_3492_data_7 <= aggregated_sig(63 downto 56);
      ptr_deref_3492_data_6 <= aggregated_sig(55 downto 48);
      ptr_deref_3492_data_5 <= aggregated_sig(47 downto 40);
      ptr_deref_3492_data_4 <= aggregated_sig(39 downto 32);
      ptr_deref_3492_data_3 <= aggregated_sig(31 downto 24);
      ptr_deref_3492_data_2 <= aggregated_sig(23 downto 16);
      ptr_deref_3492_data_1 <= aggregated_sig(15 downto 8);
      ptr_deref_3492_data_0 <= aggregated_sig(7 downto 0);
      --
    end Block;
    ptr_deref_3492_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3492_root_address_inst_ack_0 <= ptr_deref_3492_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3492_resized_base_address;
      ptr_deref_3492_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_3443_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3446_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3443_branch_req_0,
          ack0 => if_stmt_3443_branch_ack_0,
          ack1 => if_stmt_3443_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3481_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3484_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3481_branch_req_0,
          ack0 => if_stmt_3481_branch_ack_0,
          ack1 => if_stmt_3481_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3495_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3498_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3495_branch_req_0,
          ack0 => if_stmt_3495_branch_ack_0,
          ack1 => if_stmt_3495_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_3390_root_address_inst 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3390_resized_base_address;
      array_obj_ref_3390_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000010110100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3390_root_address_inst_req_0,
          ackL => array_obj_ref_3390_root_address_inst_ack_0,
          reqR => array_obj_ref_3390_root_address_inst_req_1,
          ackR => array_obj_ref_3390_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_3462_index_0_scale 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3461_resized;
      simple_obj_ref_3461_scaled <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3462_index_0_scale_req_0,
          ackL => array_obj_ref_3462_index_0_scale_ack_0,
          reqR => array_obj_ref_3462_index_0_scale_req_1,
          ackR => array_obj_ref_3462_index_0_scale_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_3462_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3462_final_offset & array_obj_ref_3462_resized_base_address;
      array_obj_ref_3462_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3462_root_address_inst_req_0,
          ackL => array_obj_ref_3462_root_address_inst_ack_0,
          reqR => array_obj_ref_3462_root_address_inst_req_1,
          ackR => array_obj_ref_3462_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_3337_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3337_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3337_inst_req_0,
          ackL => binary_3337_inst_ack_0,
          reqR => binary_3337_inst_req_1,
          ackR => binary_3337_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_3339_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3334_wire & type_cast_3338_wire;
      binary_3339_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3339_inst_req_0,
          ackL => binary_3339_inst_ack_0,
          reqR => binary_3339_inst_req_1,
          ackR => binary_3339_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_3342_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3342_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3342_inst_req_0,
          ackL => binary_3342_inst_ack_0,
          reqR => binary_3342_inst_req_1,
          ackR => binary_3342_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_3346_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3346_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3346_inst_req_0,
          ackL => binary_3346_inst_ack_0,
          reqR => binary_3346_inst_req_1,
          ackR => binary_3346_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_3348_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3343_wire & type_cast_3347_wire;
      binary_3348_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3348_inst_req_0,
          ackL => binary_3348_inst_ack_0,
          reqR => binary_3348_inst_req_1,
          ackR => binary_3348_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_3349_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3339_wire & binary_3348_wire;
      binary_3349_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3349_inst_req_0,
          ackL => binary_3349_inst_ack_0,
          reqR => binary_3349_inst_req_1,
          ackR => binary_3349_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_3352_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3352_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3352_inst_req_0,
          ackL => binary_3352_inst_ack_0,
          reqR => binary_3352_inst_req_1,
          ackR => binary_3352_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_3356_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3356_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3356_inst_req_0,
          ackL => binary_3356_inst_ack_0,
          reqR => binary_3356_inst_req_1,
          ackR => binary_3356_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_3358_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3353_wire & type_cast_3357_wire;
      binary_3358_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3358_inst_req_0,
          ackL => binary_3358_inst_ack_0,
          reqR => binary_3358_inst_req_1,
          ackR => binary_3358_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_3361_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3361_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3361_inst_req_0,
          ackL => binary_3361_inst_ack_0,
          reqR => binary_3361_inst_req_1,
          ackR => binary_3361_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_3365_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3331;
      binary_3365_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3365_inst_req_0,
          ackL => binary_3365_inst_ack_0,
          reqR => binary_3365_inst_req_1,
          ackR => binary_3365_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_3367_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3362_wire & type_cast_3366_wire;
      binary_3367_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3367_inst_req_0,
          ackL => binary_3367_inst_ack_0,
          reqR => binary_3367_inst_req_1,
          ackR => binary_3367_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_3368_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3358_wire & binary_3367_wire;
      binary_3368_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3368_inst_req_0,
          ackL => binary_3368_inst_ack_0,
          reqR => binary_3368_inst_req_1,
          ackR => binary_3368_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_3369_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3349_wire & binary_3368_wire;
      binary_3369_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3369_inst_req_0,
          ackL => binary_3369_inst_ack_0,
          reqR => binary_3369_inst_req_1,
          ackR => binary_3369_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_3446_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= hdr_in_ctrl_3441;
      binary_3446_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "11111111",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3446_inst_req_0,
          ackL => binary_3446_inst_ack_0,
          reqR => binary_3446_inst_req_1,
          ackR => binary_3446_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_3470_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_3450;
      NI_3471 <= data_out(7 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "00000001",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3470_inst_req_0,
          ackL => binary_3470_inst_ack_0,
          reqR => binary_3470_inst_req_1,
          ackR => binary_3470_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_3484_inst binary_3476_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(1 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= pkt_in_ctrl_3466 & pkt_in_ctrl_3466;
      binary_3484_wire <= data_out(1 downto 1);
      binary_3476_wire <= data_out(0 downto 0);
      reqL(1) <= binary_3484_inst_req_0;
      reqL(0) <= binary_3476_inst_req_0;
      binary_3484_inst_ack_0 <= ackL(1);
      binary_3476_inst_ack_0 <= ackL(0);
      reqR(1) <= binary_3484_inst_req_1;
      reqR(0) <= binary_3476_inst_req_1;
      binary_3484_inst_ack_1 <= ackR(1);
      binary_3476_inst_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000",
          constant_width => 8,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_3498_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3496_wire;
      binary_3498_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3498_inst_req_0,
          ackL => binary_3498_inst_ack_0,
          reqR => binary_3498_inst_req_1,
          ackR => binary_3498_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : ptr_deref_3492_addr_0 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_0_req_0,
          ackL => ptr_deref_3492_addr_0_ack_0,
          reqR => ptr_deref_3492_addr_0_req_1,
          ackR => ptr_deref_3492_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : ptr_deref_3492_addr_1 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_1_req_0,
          ackL => ptr_deref_3492_addr_1_ack_0,
          reqR => ptr_deref_3492_addr_1_req_1,
          ackR => ptr_deref_3492_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : ptr_deref_3492_addr_2 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_2_req_0,
          ackL => ptr_deref_3492_addr_2_ack_0,
          reqR => ptr_deref_3492_addr_2_req_1,
          ackR => ptr_deref_3492_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : ptr_deref_3492_addr_3 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_3_req_0,
          ackL => ptr_deref_3492_addr_3_ack_0,
          reqR => ptr_deref_3492_addr_3_req_1,
          ackR => ptr_deref_3492_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : ptr_deref_3492_addr_4 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_4 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_4_req_0,
          ackL => ptr_deref_3492_addr_4_ack_0,
          reqR => ptr_deref_3492_addr_4_req_1,
          ackR => ptr_deref_3492_addr_4_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : ptr_deref_3492_addr_5 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_5 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000101",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_5_req_0,
          ackL => ptr_deref_3492_addr_5_ack_0,
          reqR => ptr_deref_3492_addr_5_req_1,
          ackR => ptr_deref_3492_addr_5_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_3492_addr_6 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_6 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_6_req_0,
          ackL => ptr_deref_3492_addr_6_ack_0,
          reqR => ptr_deref_3492_addr_6_req_1,
          ackR => ptr_deref_3492_addr_6_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_3492_addr_7 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3492_root_address;
      ptr_deref_3492_word_address_7 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3492_addr_7_req_0,
          ackL => ptr_deref_3492_addr_7_ack_0,
          reqR => ptr_deref_3492_addr_7_req_1,
          ackR => ptr_deref_3492_addr_7_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3492_store_1_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_1 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_1) &  " data ptr_deref_3492_data_1 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_1) severity note; --
        end if;
        if ptr_deref_3492_store_6_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_6 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_6) &  " data ptr_deref_3492_data_6 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_6) severity note; --
        end if;
        if ptr_deref_3492_store_2_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_2 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_2) &  " data ptr_deref_3492_data_2 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_2) severity note; --
        end if;
        if ptr_deref_3492_store_5_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_5 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_5) &  " data ptr_deref_3492_data_5 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_5) severity note; --
        end if;
        if ptr_deref_3492_store_7_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_7 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_7) &  " data ptr_deref_3492_data_7 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_7) severity note; --
        end if;
        if ptr_deref_3492_store_4_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_4 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_4) &  " data ptr_deref_3492_data_4 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_4) severity note; --
        end if;
        if ptr_deref_3492_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_0) &  " data ptr_deref_3492_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_0) severity note; --
        end if;
        if ptr_deref_3492_store_3_ack_1 then -- 
          assert false report " WriteMem  memory_space_5 address ptr_deref_3492_word_address_3 ="  &  convert_slv_to_hex_string(ptr_deref_3492_word_address_3) &  " data ptr_deref_3492_data_3 ="  &  convert_slv_to_hex_string(ptr_deref_3492_data_3) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3492_store_1 ptr_deref_3492_store_6 ptr_deref_3492_store_2 ptr_deref_3492_store_5 ptr_deref_3492_store_7 ptr_deref_3492_store_4 ptr_deref_3492_store_0 ptr_deref_3492_store_3 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(127 downto 0);
      signal data_in: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      reqL(7) <= ptr_deref_3492_store_1_req_0;
      reqL(6) <= ptr_deref_3492_store_6_req_0;
      reqL(5) <= ptr_deref_3492_store_2_req_0;
      reqL(4) <= ptr_deref_3492_store_5_req_0;
      reqL(3) <= ptr_deref_3492_store_7_req_0;
      reqL(2) <= ptr_deref_3492_store_4_req_0;
      reqL(1) <= ptr_deref_3492_store_0_req_0;
      reqL(0) <= ptr_deref_3492_store_3_req_0;
      ptr_deref_3492_store_1_ack_0 <= ackL(7);
      ptr_deref_3492_store_6_ack_0 <= ackL(6);
      ptr_deref_3492_store_2_ack_0 <= ackL(5);
      ptr_deref_3492_store_5_ack_0 <= ackL(4);
      ptr_deref_3492_store_7_ack_0 <= ackL(3);
      ptr_deref_3492_store_4_ack_0 <= ackL(2);
      ptr_deref_3492_store_0_ack_0 <= ackL(1);
      ptr_deref_3492_store_3_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_3492_store_1_req_1;
      reqR(6) <= ptr_deref_3492_store_6_req_1;
      reqR(5) <= ptr_deref_3492_store_2_req_1;
      reqR(4) <= ptr_deref_3492_store_5_req_1;
      reqR(3) <= ptr_deref_3492_store_7_req_1;
      reqR(2) <= ptr_deref_3492_store_4_req_1;
      reqR(1) <= ptr_deref_3492_store_0_req_1;
      reqR(0) <= ptr_deref_3492_store_3_req_1;
      ptr_deref_3492_store_1_ack_1 <= ackR(7);
      ptr_deref_3492_store_6_ack_1 <= ackR(6);
      ptr_deref_3492_store_2_ack_1 <= ackR(5);
      ptr_deref_3492_store_5_ack_1 <= ackR(4);
      ptr_deref_3492_store_7_ack_1 <= ackR(3);
      ptr_deref_3492_store_4_ack_1 <= ackR(2);
      ptr_deref_3492_store_0_ack_1 <= ackR(1);
      ptr_deref_3492_store_3_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3492_word_address_1 & ptr_deref_3492_word_address_6 & ptr_deref_3492_word_address_2 & ptr_deref_3492_word_address_5 & ptr_deref_3492_word_address_7 & ptr_deref_3492_word_address_4 & ptr_deref_3492_word_address_0 & ptr_deref_3492_word_address_3;
      data_in <= ptr_deref_3492_data_1 & ptr_deref_3492_data_6 & ptr_deref_3492_data_2 & ptr_deref_3492_data_5 & ptr_deref_3492_data_7 & ptr_deref_3492_data_4 & ptr_deref_3492_data_0 & ptr_deref_3492_data_3;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 16,
        data_width => 8,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_5_sr_req(0),
          mack => memory_space_5_sr_ack(0),
          maddr => memory_space_5_sr_addr(15 downto 0),
          mdata => memory_space_5_sr_data(7 downto 0),
          mtag => memory_space_5_sr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 5 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_5_sc_req(0),
          mack => memory_space_5_sc_ack(0),
          mtag => memory_space_5_sc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    xxreceive_packet_pipelinexxbuf64_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxbuf8_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxpkt64_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxpkt8_ptr_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_last_word_flag_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 4 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxreceive_packet_pipelinexxwrite_data_wptr_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req,
        read_ack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack,
        read_data => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data,
        write_req => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req,
        write_ack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack,
        write_data => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : simple_obj_ref_3330_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3330_inst_ack_0 then -- 
            assert false report " ReadPipe in_data to wire a_3331 value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3330_inst_req_0;
      simple_obj_ref_3330_inst_ack_0 <= ack(0);
      a_3331 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_read_req(0),
          oack => in_data_pipe_read_ack(0),
          odata => in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_3377_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3377_inst_ack_0 then -- 
            assert false report " ReadPipe free_queue_pipe to wire buf_3378 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3377_inst_req_0;
      simple_obj_ref_3377_inst_ack_0 <= ack(0);
      buf_3378 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => free_queue_pipe_pipe_read_req(0),
          oack => free_queue_pipe_pipe_read_ack(0),
          odata => free_queue_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_3416_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3416_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxbuf8_ptr_pipe to wire buf8_ptr_3417 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3416_inst_req_0;
      simple_obj_ref_3416_inst_ack_0 <= ack(0);
      buf8_ptr_3417 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_3419_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3419_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxbuf64_ptr_pipe to wire buf64_ptr_3420 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3419_inst_req_0;
      simple_obj_ref_3419_inst_ack_0 <= ack(0);
      buf64_ptr_3420 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_3422_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3422_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxpkt8_ptr_pipe to wire pkt8_ptr_3423 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3422_inst_req_0;
      simple_obj_ref_3422_inst_ack_0 <= ack(0);
      pkt8_ptr_3423 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : simple_obj_ref_3425_inst 
    InportGroup5: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3425_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxpkt64_ptr_pipe to wire pkt64_ptr_3426 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3425_inst_req_0;
      simple_obj_ref_3425_inst_ack_0 <= ack(0);
      pkt64_ptr_3426 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : simple_obj_ref_3431_inst simple_obj_ref_3458_inst 
    InportGroup6: Block -- 
      signal data_out: std_logic_vector(127 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3431_inst_ack_0 then -- 
            assert false report " ReadPipe swapped_in_data to wire simple_obj_ref_3431_wire value="  &  convert_slv_to_hex_string(data_out(127 downto 64))  severity note; --
          end if;
          if simple_obj_ref_3458_inst_ack_0 then -- 
            assert false report " ReadPipe swapped_in_data to wire simple_obj_ref_3458_wire value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(1) <= simple_obj_ref_3431_inst_req_0;
      req(0) <= simple_obj_ref_3458_inst_req_0;
      simple_obj_ref_3431_inst_ack_0 <= ack(1);
      simple_obj_ref_3458_inst_ack_0 <= ack(0);
      simple_obj_ref_3431_wire <= data_out(127 downto 64);
      simple_obj_ref_3458_wire <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 2,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => swapped_in_data_pipe_read_req(0),
          oack => swapped_in_data_pipe_read_ack(0),
          odata => swapped_in_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : simple_obj_ref_3440_inst simple_obj_ref_3465_inst 
    InportGroup7: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3440_inst_ack_0 then -- 
            assert false report " ReadPipe in_ctrl to wire hdr_in_ctrl_3441 value="  &  convert_slv_to_hex_string(data_out(15 downto 8))  severity note; --
          end if;
          if simple_obj_ref_3465_inst_ack_0 then -- 
            assert false report " ReadPipe in_ctrl to wire pkt_in_ctrl_3466 value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(1) <= simple_obj_ref_3440_inst_req_0;
      req(0) <= simple_obj_ref_3465_inst_req_0;
      simple_obj_ref_3440_inst_ack_0 <= ack(1);
      simple_obj_ref_3465_inst_ack_0 <= ack(0);
      hdr_in_ctrl_3441 <= data_out(15 downto 8);
      pkt_in_ctrl_3466 <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 2,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_ctrl_pipe_read_req(0),
          oack => in_ctrl_pipe_read_ack(0),
          odata => in_ctrl_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : simple_obj_ref_3491_inst 
    InportGroup8: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3491_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data_wptr to wire simple_obj_ref_3491_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3491_inst_req_0;
      simple_obj_ref_3491_inst_ack_0 <= ack(0);
      simple_obj_ref_3491_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : simple_obj_ref_3493_inst 
    InportGroup9: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3493_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data to wire simple_obj_ref_3493_wire value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3493_inst_req_0;
      simple_obj_ref_3493_inst_ack_0 <= ack(0);
      simple_obj_ref_3493_wire <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : simple_obj_ref_3496_inst 
    InportGroup10: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3496_inst_ack_0 then -- 
            assert false report " ReadPipe xxreceive_packet_pipelinexxwrite_data_last_word_flag to wire simple_obj_ref_3496_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3496_inst_req_0;
      simple_obj_ref_3496_inst_ack_0 <= ack(0);
      simple_obj_ref_3496_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : simple_obj_ref_3500_inst 
    InportGroup11: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3500_inst_ack_0 then -- 
            assert false report " ReadPipe receive_packet_buf_queue to wire simple_obj_ref_3500_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3500_inst_req_0;
      simple_obj_ref_3500_inst_ack_0 <= ack(0);
      simple_obj_ref_3500_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => receive_packet_buf_queue_pipe_read_req(0),
          oack => receive_packet_buf_queue_pipe_read_ack(0),
          odata => receive_packet_buf_queue_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3332_inst_ack_0 then -- 
          assert false report " WritePipe swapped_in_data from wire binary_3369_wire value="  &  convert_slv_to_hex_string(binary_3369_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3332_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3332_inst_req_0;
      simple_obj_ref_3332_inst_ack_0 <= ack(0);
      data_in <= binary_3369_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => swapped_in_data_pipe_write_req(0),
          oack => swapped_in_data_pipe_write_ack(0),
          odata => swapped_in_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3393_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxbuf8_ptr_pipe from wire buf8_ptr_3383 value="  &  convert_slv_to_hex_string(buf8_ptr_3383) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_3393_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3393_inst_req_0;
      simple_obj_ref_3393_inst_ack_0 <= ack(0);
      data_in <= buf8_ptr_3383;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxbuf8_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3396_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxbuf64_ptr_pipe from wire buf64_ptr_3387 value="  &  convert_slv_to_hex_string(buf64_ptr_3387) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_3396_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3396_inst_req_0;
      simple_obj_ref_3396_inst_ack_0 <= ack(0);
      data_in <= buf64_ptr_3387;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxbuf64_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3399_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxpkt8_ptr_pipe from wire pkt8_ptr_3391 value="  &  convert_slv_to_hex_string(pkt8_ptr_3391) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_3399_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3399_inst_req_0;
      simple_obj_ref_3399_inst_ack_0 <= ack(0);
      data_in <= pkt8_ptr_3391;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxpkt8_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3402_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxpkt64_ptr_pipe from wire type_cast_3404_wire value="  &  convert_slv_to_hex_string(type_cast_3404_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (4) : simple_obj_ref_3402_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3402_inst_req_0;
      simple_obj_ref_3402_inst_ack_0 <= ack(0);
      data_in <= type_cast_3404_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxpkt64_ptr_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3406_inst_ack_0 then -- 
          assert false report " WritePipe receive_packet_buf_queue from wire buf_3378 value="  &  convert_slv_to_hex_string(buf_3378) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (5) : simple_obj_ref_3406_inst 
    OutportGroup5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3406_inst_req_0;
      simple_obj_ref_3406_inst_ack_0 <= ack(0);
      data_in <= buf_3378;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => receive_packet_buf_queue_pipe_write_req(0),
          oack => receive_packet_buf_queue_pipe_write_ack(0),
          odata => receive_packet_buf_queue_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3430_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data from wire simple_obj_ref_3431_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3431_wire) severity note; --
        end if;
        if simple_obj_ref_3457_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data from wire simple_obj_ref_3458_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3458_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (6) : simple_obj_ref_3430_inst simple_obj_ref_3457_inst 
    OutportGroup6: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_3430_inst_req_0;
      req(0) <= simple_obj_ref_3457_inst_req_0;
      simple_obj_ref_3430_inst_ack_0 <= ack(1);
      simple_obj_ref_3457_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3431_wire & simple_obj_ref_3458_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3433_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_last_word_flag from wire expr_3434_wire_constant value="  &  convert_slv_to_hex_string(expr_3434_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3473_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_last_word_flag from wire ternary_3479_wire value="  &  convert_slv_to_hex_string(ternary_3479_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (7) : simple_obj_ref_3433_inst simple_obj_ref_3473_inst 
    OutportGroup7: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_3433_inst_req_0;
      req(0) <= simple_obj_ref_3473_inst_req_0;
      simple_obj_ref_3433_inst_ack_0 <= ack(1);
      simple_obj_ref_3473_inst_ack_0 <= ack(0);
      data_in <= expr_3434_wire_constant & ternary_3479_wire;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_last_word_flag_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3436_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_wptr from wire buf64_ptr_3420 value="  &  convert_slv_to_hex_string(buf64_ptr_3420) severity note; --
        end if;
        if simple_obj_ref_3460_inst_ack_0 then -- 
          assert false report " WritePipe xxreceive_packet_pipelinexxwrite_data_wptr from wire array_obj_ref_3462_wire value="  &  convert_slv_to_hex_string(array_obj_ref_3462_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (8) : simple_obj_ref_3436_inst simple_obj_ref_3460_inst 
    OutportGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      req(1) <= simple_obj_ref_3436_inst_req_0;
      req(0) <= simple_obj_ref_3460_inst_req_0;
      simple_obj_ref_3436_inst_ack_0 <= ack(1);
      simple_obj_ref_3460_inst_ack_0 <= ack(0);
      data_in <= buf64_ptr_3420 & array_obj_ref_3462_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 2,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_req(0),
          oack => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_ack(0),
          odata => xxreceive_packet_pipelinexxwrite_data_wptr_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3499_inst_ack_0 then -- 
          assert false report " WritePipe receive_packet_pipe from wire type_cast_3501_wire value="  &  convert_slv_to_hex_string(type_cast_3501_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (9) : simple_obj_ref_3499_inst 
    OutportGroup9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3499_inst_req_0;
      simple_obj_ref_3499_inst_ack_0 <= ack(0);
      data_in <= type_cast_3501_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => receive_packet_pipe_pipe_write_req(0),
          oack => receive_packet_pipe_pipe_write_ack(0),
          odata => receive_packet_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 9
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity send_packet_pipeline is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
    memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
    memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
    memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
    send_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
    send_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
    out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
    send_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
    send_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
    analyze_packet_call_reqs : out  std_logic_vector(0 downto 0);
    analyze_packet_call_acks : in   std_logic_vector(0 downto 0);
    analyze_packet_call_data : out  std_logic_vector(31 downto 0);
    analyze_packet_call_tag  :  out  std_logic_vector(0 downto 0);
    analyze_packet_return_reqs : out  std_logic_vector(0 downto 0);
    analyze_packet_return_acks : in   std_logic_vector(0 downto 0);
    analyze_packet_return_data : in   std_logic_vector(63 downto 0);
    analyze_packet_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity send_packet_pipeline;
architecture Default of send_packet_pipeline is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal send_packet_pipeline_CP_17966_start: Boolean;
  -- links between control-path and data-path
  signal binary_3707_inst_ack_0 : boolean;
  signal binary_3705_inst_req_0 : boolean;
  signal binary_3703_inst_ack_0 : boolean;
  signal binary_3706_inst_ack_0 : boolean;
  signal simple_obj_ref_3725_inst_req_0 : boolean;
  signal binary_3728_inst_req_0 : boolean;
  signal simple_obj_ref_3709_inst_ack_0 : boolean;
  signal type_cast_3704_inst_ack_0 : boolean;
  signal simple_obj_ref_3713_inst_req_0 : boolean;
  signal binary_3728_inst_ack_1 : boolean;
  signal binary_3728_inst_req_1 : boolean;
  signal binary_3705_inst_ack_1 : boolean;
  signal binary_3707_inst_req_0 : boolean;
  signal binary_3703_inst_req_0 : boolean;
  signal simple_obj_ref_3725_inst_ack_0 : boolean;
  signal binary_3705_inst_ack_0 : boolean;
  signal type_cast_3704_inst_req_0 : boolean;
  signal type_cast_3700_inst_ack_0 : boolean;
  signal binary_3705_inst_req_1 : boolean;
  signal simple_obj_ref_3710_inst_ack_0 : boolean;
  signal simple_obj_ref_3670_inst_req_0 : boolean;
  signal simple_obj_ref_3709_inst_req_0 : boolean;
  signal simple_obj_ref_3670_inst_ack_0 : boolean;
  signal binary_3703_inst_ack_1 : boolean;
  signal if_stmt_3720_branch_ack_0 : boolean;
  signal binary_3706_inst_req_0 : boolean;
  signal simple_obj_ref_3712_inst_req_0 : boolean;
  signal binary_3706_inst_req_1 : boolean;
  signal simple_obj_ref_3712_inst_ack_0 : boolean;
  signal simple_obj_ref_3726_inst_ack_0 : boolean;
  signal binary_3706_inst_ack_1 : boolean;
  signal binary_3703_inst_req_1 : boolean;
  signal binary_3707_inst_ack_1 : boolean;
  signal binary_3728_inst_ack_0 : boolean;
  signal simple_obj_ref_3726_inst_req_0 : boolean;
  signal simple_obj_ref_3713_inst_ack_0 : boolean;
  signal type_cast_3700_inst_req_0 : boolean;
  signal binary_3707_inst_req_1 : boolean;
  signal ptr_deref_3653_addr_0_req_0 : boolean;
  signal ptr_deref_3653_addr_0_ack_0 : boolean;
  signal ptr_deref_3653_addr_0_req_1 : boolean;
  signal ptr_deref_3653_root_address_inst_req_0 : boolean;
  signal ptr_deref_3653_base_resize_req_0 : boolean;
  signal ptr_deref_3653_base_resize_ack_0 : boolean;
  signal phi_stmt_3591_req_0 : boolean;
  signal phi_stmt_3591_req_1 : boolean;
  signal simple_obj_ref_3652_inst_req_0 : boolean;
  signal ptr_deref_3653_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3653_addr_1_req_0 : boolean;
  signal ptr_deref_3653_addr_1_ack_0 : boolean;
  signal simple_obj_ref_3652_inst_ack_0 : boolean;
  signal ptr_deref_3653_addr_0_ack_1 : boolean;
  signal phi_stmt_3591_ack_0 : boolean;
  signal simple_obj_ref_3710_inst_req_0 : boolean;
  signal simple_obj_ref_3524_inst_req_0 : boolean;
  signal simple_obj_ref_3524_inst_ack_0 : boolean;
  signal type_cast_3527_inst_req_0 : boolean;
  signal type_cast_3527_inst_ack_0 : boolean;
  signal call_stmt_3531_call_req_0 : boolean;
  signal call_stmt_3531_call_ack_0 : boolean;
  signal call_stmt_3531_call_req_1 : boolean;
  signal call_stmt_3531_call_ack_1 : boolean;
  signal type_cast_3535_inst_req_0 : boolean;
  signal type_cast_3535_inst_ack_0 : boolean;
  signal simple_obj_ref_3533_inst_req_0 : boolean;
  signal simple_obj_ref_3533_inst_ack_0 : boolean;
  signal type_cast_3539_inst_req_0 : boolean;
  signal type_cast_3539_inst_ack_0 : boolean;
  signal simple_obj_ref_3537_inst_req_0 : boolean;
  signal simple_obj_ref_3537_inst_ack_0 : boolean;
  signal simple_obj_ref_3541_inst_req_0 : boolean;
  signal simple_obj_ref_3541_inst_ack_0 : boolean;
  signal simple_obj_ref_3544_inst_req_0 : boolean;
  signal simple_obj_ref_3544_inst_ack_0 : boolean;
  signal type_cast_3549_inst_req_0 : boolean;
  signal type_cast_3549_inst_ack_0 : boolean;
  signal simple_obj_ref_3547_inst_req_0 : boolean;
  signal simple_obj_ref_3547_inst_ack_0 : boolean;
  signal simple_obj_ref_3558_inst_req_0 : boolean;
  signal simple_obj_ref_3558_inst_ack_0 : boolean;
  signal simple_obj_ref_3561_inst_req_0 : boolean;
  signal simple_obj_ref_3561_inst_ack_0 : boolean;
  signal simple_obj_ref_3564_inst_req_0 : boolean;
  signal simple_obj_ref_3564_inst_ack_0 : boolean;
  signal simple_obj_ref_3567_inst_req_0 : boolean;
  signal simple_obj_ref_3567_inst_ack_0 : boolean;
  signal binary_3573_inst_req_0 : boolean;
  signal binary_3573_inst_ack_0 : boolean;
  signal binary_3573_inst_req_1 : boolean;
  signal binary_3573_inst_ack_1 : boolean;
  signal if_stmt_3570_branch_req_0 : boolean;
  signal if_stmt_3570_branch_ack_1 : boolean;
  signal if_stmt_3570_branch_ack_0 : boolean;
  signal simple_obj_ref_3575_inst_req_0 : boolean;
  signal simple_obj_ref_3575_inst_ack_0 : boolean;
  signal simple_obj_ref_3578_inst_req_0 : boolean;
  signal simple_obj_ref_3578_inst_ack_0 : boolean;
  signal simple_obj_ref_3581_inst_req_0 : boolean;
  signal simple_obj_ref_3581_inst_ack_0 : boolean;
  signal binary_3587_inst_req_0 : boolean;
  signal binary_3587_inst_ack_0 : boolean;
  signal binary_3587_inst_req_1 : boolean;
  signal binary_3587_inst_ack_1 : boolean;
  signal simple_obj_ref_3598_inst_req_0 : boolean;
  signal simple_obj_ref_3598_inst_ack_0 : boolean;
  signal array_obj_ref_3603_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3603_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_3603_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3603_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3603_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3603_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_3603_offset_inst_req_0 : boolean;
  signal array_obj_ref_3603_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3603_base_resize_req_0 : boolean;
  signal array_obj_ref_3603_base_resize_ack_0 : boolean;
  signal array_obj_ref_3603_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3603_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3603_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3603_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3603_final_reg_req_0 : boolean;
  signal array_obj_ref_3603_final_reg_ack_0 : boolean;
  signal simple_obj_ref_3601_inst_req_0 : boolean;
  signal simple_obj_ref_3601_inst_ack_0 : boolean;
  signal simple_obj_ref_3605_inst_req_0 : boolean;
  signal simple_obj_ref_3605_inst_ack_0 : boolean;
  signal binary_3611_inst_req_0 : boolean;
  signal binary_3611_inst_ack_0 : boolean;
  signal binary_3611_inst_req_1 : boolean;
  signal binary_3611_inst_ack_1 : boolean;
  signal binary_3617_inst_req_0 : boolean;
  signal binary_3617_inst_ack_0 : boolean;
  signal binary_3617_inst_req_1 : boolean;
  signal binary_3617_inst_ack_1 : boolean;
  signal if_stmt_3614_branch_req_0 : boolean;
  signal if_stmt_3614_branch_ack_1 : boolean;
  signal if_stmt_3614_branch_ack_0 : boolean;
  signal array_obj_ref_3622_index_0_resize_req_0 : boolean;
  signal array_obj_ref_3622_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_3622_index_0_scale_req_0 : boolean;
  signal array_obj_ref_3622_index_0_scale_ack_0 : boolean;
  signal array_obj_ref_3622_index_0_scale_req_1 : boolean;
  signal array_obj_ref_3622_index_0_scale_ack_1 : boolean;
  signal array_obj_ref_3622_offset_inst_req_0 : boolean;
  signal array_obj_ref_3622_offset_inst_ack_0 : boolean;
  signal array_obj_ref_3622_base_resize_req_0 : boolean;
  signal array_obj_ref_3622_base_resize_ack_0 : boolean;
  signal array_obj_ref_3622_root_address_inst_req_0 : boolean;
  signal array_obj_ref_3622_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_3622_root_address_inst_req_1 : boolean;
  signal array_obj_ref_3622_root_address_inst_ack_1 : boolean;
  signal array_obj_ref_3622_final_reg_req_0 : boolean;
  signal array_obj_ref_3622_final_reg_ack_0 : boolean;
  signal binary_3631_inst_req_0 : boolean;
  signal binary_3631_inst_ack_0 : boolean;
  signal binary_3631_inst_req_1 : boolean;
  signal binary_3631_inst_ack_1 : boolean;
  signal binary_3632_inst_req_0 : boolean;
  signal binary_3632_inst_ack_0 : boolean;
  signal binary_3632_inst_req_1 : boolean;
  signal binary_3632_inst_ack_1 : boolean;
  signal binary_3634_inst_req_0 : boolean;
  signal binary_3634_inst_ack_0 : boolean;
  signal binary_3634_inst_req_1 : boolean;
  signal binary_3634_inst_ack_1 : boolean;
  signal type_cast_3635_inst_req_0 : boolean;
  signal type_cast_3635_inst_ack_0 : boolean;
  signal binary_3636_inst_req_0 : boolean;
  signal binary_3636_inst_ack_0 : boolean;
  signal binary_3636_inst_req_1 : boolean;
  signal binary_3636_inst_ack_1 : boolean;
  signal simple_obj_ref_3625_inst_req_0 : boolean;
  signal simple_obj_ref_3625_inst_ack_0 : boolean;
  signal simple_obj_ref_3638_inst_req_0 : boolean;
  signal simple_obj_ref_3638_inst_ack_0 : boolean;
  signal simple_obj_ref_3641_inst_req_0 : boolean;
  signal simple_obj_ref_3641_inst_ack_0 : boolean;
  signal ptr_deref_3653_addr_1_req_1 : boolean;
  signal ptr_deref_3653_addr_1_ack_1 : boolean;
  signal ptr_deref_3653_addr_2_req_0 : boolean;
  signal ptr_deref_3653_addr_2_ack_0 : boolean;
  signal ptr_deref_3653_addr_2_req_1 : boolean;
  signal ptr_deref_3653_addr_2_ack_1 : boolean;
  signal ptr_deref_3653_addr_3_req_0 : boolean;
  signal ptr_deref_3653_addr_3_ack_0 : boolean;
  signal ptr_deref_3653_addr_3_req_1 : boolean;
  signal ptr_deref_3653_addr_3_ack_1 : boolean;
  signal ptr_deref_3653_addr_4_req_0 : boolean;
  signal ptr_deref_3653_addr_4_ack_0 : boolean;
  signal ptr_deref_3653_addr_4_req_1 : boolean;
  signal ptr_deref_3653_addr_4_ack_1 : boolean;
  signal ptr_deref_3653_addr_5_req_0 : boolean;
  signal ptr_deref_3653_addr_5_ack_0 : boolean;
  signal ptr_deref_3653_addr_5_req_1 : boolean;
  signal ptr_deref_3653_addr_5_ack_1 : boolean;
  signal ptr_deref_3653_addr_6_req_0 : boolean;
  signal ptr_deref_3653_addr_6_ack_0 : boolean;
  signal ptr_deref_3653_addr_6_req_1 : boolean;
  signal ptr_deref_3653_addr_6_ack_1 : boolean;
  signal ptr_deref_3653_addr_7_req_0 : boolean;
  signal ptr_deref_3653_addr_7_ack_0 : boolean;
  signal ptr_deref_3653_addr_7_req_1 : boolean;
  signal ptr_deref_3653_addr_7_ack_1 : boolean;
  signal ptr_deref_3653_load_0_req_0 : boolean;
  signal ptr_deref_3653_load_0_ack_0 : boolean;
  signal ptr_deref_3653_load_1_req_0 : boolean;
  signal ptr_deref_3653_load_1_ack_0 : boolean;
  signal ptr_deref_3653_load_2_req_0 : boolean;
  signal ptr_deref_3653_load_2_ack_0 : boolean;
  signal ptr_deref_3653_load_3_req_0 : boolean;
  signal ptr_deref_3653_load_3_ack_0 : boolean;
  signal ptr_deref_3653_load_4_req_0 : boolean;
  signal ptr_deref_3653_load_4_ack_0 : boolean;
  signal ptr_deref_3653_load_5_req_0 : boolean;
  signal ptr_deref_3653_load_5_ack_0 : boolean;
  signal ptr_deref_3653_load_6_req_0 : boolean;
  signal ptr_deref_3653_load_6_ack_0 : boolean;
  signal ptr_deref_3653_load_7_req_0 : boolean;
  signal ptr_deref_3653_load_7_ack_0 : boolean;
  signal ptr_deref_3653_load_0_req_1 : boolean;
  signal ptr_deref_3653_load_0_ack_1 : boolean;
  signal ptr_deref_3653_load_1_req_1 : boolean;
  signal ptr_deref_3653_load_1_ack_1 : boolean;
  signal ptr_deref_3653_load_2_req_1 : boolean;
  signal ptr_deref_3653_load_2_ack_1 : boolean;
  signal ptr_deref_3653_load_3_req_1 : boolean;
  signal ptr_deref_3653_load_3_ack_1 : boolean;
  signal ptr_deref_3653_load_4_req_1 : boolean;
  signal ptr_deref_3653_load_4_ack_1 : boolean;
  signal ptr_deref_3653_load_5_req_1 : boolean;
  signal ptr_deref_3653_load_5_ack_1 : boolean;
  signal ptr_deref_3653_load_6_req_1 : boolean;
  signal ptr_deref_3653_load_6_ack_1 : boolean;
  signal ptr_deref_3653_load_7_req_1 : boolean;
  signal ptr_deref_3653_load_7_ack_1 : boolean;
  signal ptr_deref_3653_gather_scatter_req_0 : boolean;
  signal ptr_deref_3653_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_3651_inst_req_0 : boolean;
  signal simple_obj_ref_3651_inst_ack_0 : boolean;
  signal if_stmt_3720_branch_ack_1 : boolean;
  signal if_stmt_3720_branch_req_0 : boolean;
  signal binary_3723_inst_ack_1 : boolean;
  signal simple_obj_ref_3656_inst_req_0 : boolean;
  signal binary_3723_inst_req_1 : boolean;
  signal simple_obj_ref_3656_inst_ack_0 : boolean;
  signal binary_3723_inst_ack_0 : boolean;
  signal binary_3723_inst_req_0 : boolean;
  signal simple_obj_ref_3655_inst_req_0 : boolean;
  signal simple_obj_ref_3721_inst_ack_0 : boolean;
  signal simple_obj_ref_3655_inst_ack_0 : boolean;
  signal simple_obj_ref_3721_inst_req_0 : boolean;
  signal simple_obj_ref_3659_inst_req_0 : boolean;
  signal simple_obj_ref_3659_inst_ack_0 : boolean;
  signal simple_obj_ref_3658_inst_req_0 : boolean;
  signal simple_obj_ref_3658_inst_ack_0 : boolean;
  signal simple_obj_ref_3667_inst_req_0 : boolean;
  signal simple_obj_ref_3667_inst_ack_0 : boolean;
  signal type_cast_3672_inst_req_0 : boolean;
  signal type_cast_3672_inst_ack_0 : boolean;
  signal binary_3675_inst_req_0 : boolean;
  signal binary_3675_inst_ack_0 : boolean;
  signal binary_3675_inst_req_1 : boolean;
  signal binary_3675_inst_ack_1 : boolean;
  signal type_cast_3676_inst_req_0 : boolean;
  signal type_cast_3676_inst_ack_0 : boolean;
  signal binary_3677_inst_req_0 : boolean;
  signal binary_3677_inst_ack_0 : boolean;
  signal binary_3677_inst_req_1 : boolean;
  signal binary_3677_inst_ack_1 : boolean;
  signal binary_3680_inst_req_0 : boolean;
  signal binary_3680_inst_ack_0 : boolean;
  signal binary_3680_inst_req_1 : boolean;
  signal binary_3680_inst_ack_1 : boolean;
  signal type_cast_3681_inst_req_0 : boolean;
  signal type_cast_3681_inst_ack_0 : boolean;
  signal binary_3684_inst_req_0 : boolean;
  signal binary_3684_inst_ack_0 : boolean;
  signal binary_3684_inst_req_1 : boolean;
  signal binary_3684_inst_ack_1 : boolean;
  signal type_cast_3685_inst_req_0 : boolean;
  signal type_cast_3685_inst_ack_0 : boolean;
  signal binary_3686_inst_req_0 : boolean;
  signal binary_3686_inst_ack_0 : boolean;
  signal binary_3686_inst_req_1 : boolean;
  signal binary_3686_inst_ack_1 : boolean;
  signal binary_3687_inst_req_0 : boolean;
  signal binary_3687_inst_ack_0 : boolean;
  signal binary_3687_inst_req_1 : boolean;
  signal binary_3687_inst_ack_1 : boolean;
  signal binary_3690_inst_req_0 : boolean;
  signal binary_3690_inst_ack_0 : boolean;
  signal binary_3690_inst_req_1 : boolean;
  signal binary_3690_inst_ack_1 : boolean;
  signal type_cast_3691_inst_req_0 : boolean;
  signal type_cast_3691_inst_ack_0 : boolean;
  signal binary_3694_inst_req_0 : boolean;
  signal binary_3694_inst_ack_0 : boolean;
  signal binary_3694_inst_req_1 : boolean;
  signal binary_3694_inst_ack_1 : boolean;
  signal type_cast_3695_inst_req_0 : boolean;
  signal type_cast_3695_inst_ack_0 : boolean;
  signal binary_3696_inst_req_0 : boolean;
  signal binary_3696_inst_ack_0 : boolean;
  signal binary_3696_inst_req_1 : boolean;
  signal binary_3696_inst_ack_1 : boolean;
  signal binary_3699_inst_req_0 : boolean;
  signal binary_3699_inst_ack_0 : boolean;
  signal binary_3699_inst_req_1 : boolean;
  signal binary_3699_inst_ack_1 : boolean;
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  send_packet_pipeline_CP_17966: Block -- control-path 
    signal cp_elements: BooleanArray(402 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(402);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(402), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(0);
    cp_elements(2) <= false; 
    cp_elements(3) <= OrReduce(cp_elements(39) & cp_elements(42));
    req_17995_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => simple_obj_ref_3524_inst_req_0); -- 
    cp_elements(4) <= cp_elements(36);
    ack_17996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3524_inst_ack_0, ack => cp_elements(5)); -- 
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(8) & cp_elements(9));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18006_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => type_cast_3527_inst_req_0); -- 
    cp_elements(8) <= cp_elements(6);
    cp_elements(9) <= cp_elements(6);
    ack_18007_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3527_inst_ack_0, ack => cp_elements(10)); -- 
    crr_18013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => call_stmt_3531_call_req_0); -- 
    cra_18014_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3531_call_ack_0, ack => cp_elements(11)); -- 
    ccr_18018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => call_stmt_3531_call_req_1); -- 
    cca_18019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3531_call_ack_1, ack => cp_elements(12)); -- 
    cp_elements(13) <= cp_elements(12);
    cp_elements(14) <= cp_elements(13);
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(17));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => type_cast_3535_inst_req_0); -- 
    cp_elements(16) <= cp_elements(14);
    cp_elements(17) <= cp_elements(14);
    ack_18037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3535_inst_ack_0, ack => cp_elements(18)); -- 
    pipe_wreq_18042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => simple_obj_ref_3533_inst_req_0); -- 
    pipe_wack_18043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3533_inst_ack_0, ack => cp_elements(19)); -- 
    cp_elements(20) <= cp_elements(13);
    cpelement_group_21 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(22) & cp_elements(23));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(21),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18055_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => type_cast_3539_inst_req_0); -- 
    cp_elements(22) <= cp_elements(20);
    cp_elements(23) <= cp_elements(20);
    ack_18056_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3539_inst_ack_0, ack => cp_elements(24)); -- 
    pipe_wreq_18061_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => simple_obj_ref_3537_inst_req_0); -- 
    pipe_wack_18062_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3537_inst_ack_0, ack => cp_elements(25)); -- 
    cp_elements(26) <= cp_elements(13);
    pipe_wreq_18073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => simple_obj_ref_3541_inst_req_0); -- 
    pipe_wack_18074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3541_inst_ack_0, ack => cp_elements(27)); -- 
    cp_elements(28) <= cp_elements(13);
    pipe_wreq_18085_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => simple_obj_ref_3544_inst_req_0); -- 
    pipe_wack_18086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3544_inst_ack_0, ack => cp_elements(29)); -- 
    cp_elements(30) <= cp_elements(13);
    cpelement_group_31 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(32) & cp_elements(33));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(31),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18098_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => type_cast_3549_inst_req_0); -- 
    cp_elements(32) <= cp_elements(30);
    cp_elements(33) <= cp_elements(30);
    ack_18099_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3549_inst_ack_0, ack => cp_elements(34)); -- 
    pipe_wreq_18104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => simple_obj_ref_3547_inst_req_0); -- 
    pipe_wack_18105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3547_inst_ack_0, ack => cp_elements(35)); -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(25) & cp_elements(27) & cp_elements(29) & cp_elements(35));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(37) <= cp_elements(1);
    cp_elements(38) <= false;
    cp_elements(39) <= cp_elements(38);
    cp_elements(40) <= cp_elements(1);
    cp_elements(41) <= OrReduce(cp_elements(4) & cp_elements(40));
    cp_elements(42) <= cp_elements(41);
    cp_elements(43) <= cp_elements(0);
    cp_elements(44) <= false; 
    cp_elements(45) <= OrReduce(cp_elements(177) & cp_elements(180));
    cp_elements(46) <= cp_elements(57);
    cp_elements(47) <= OrReduce(cp_elements(60) & cp_elements(68) & cp_elements(73));
    cp_elements(48) <= cp_elements(45);
    cp_elements(49) <= cp_elements(48);
    req_18145_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => simple_obj_ref_3558_inst_req_0); -- 
    ack_18146_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3558_inst_ack_0, ack => cp_elements(50)); -- 
    cp_elements(51) <= cp_elements(48);
    req_18156_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => simple_obj_ref_3561_inst_req_0); -- 
    ack_18157_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3561_inst_ack_0, ack => cp_elements(52)); -- 
    cp_elements(53) <= cp_elements(48);
    req_18167_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => simple_obj_ref_3564_inst_req_0); -- 
    ack_18168_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3564_inst_ack_0, ack => cp_elements(54)); -- 
    cp_elements(55) <= cp_elements(48);
    req_18178_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => simple_obj_ref_3567_inst_req_0); -- 
    ack_18179_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3567_inst_ack_0, ack => cp_elements(56)); -- 
    cpelement_group_57 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(50) & cp_elements(52) & cp_elements(54) & cp_elements(56));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(57),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(58) <= cp_elements(46);
    cp_elements(59) <= false;
    cp_elements(60) <= cp_elements(59);
    cp_elements(61) <= cp_elements(46);
    rr_18193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => binary_3573_inst_req_0); -- 
    ra_18194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3573_inst_ack_0, ack => cp_elements(62)); -- 
    cr_18195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => binary_3573_inst_req_1); -- 
    ca_18196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3573_inst_ack_1, ack => cp_elements(63)); -- 
    branch_req_18197_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => if_stmt_3570_branch_req_0); -- 
    cp_elements(64) <= cp_elements(63);
    cp_elements(65) <= cp_elements(64);
    if_choice_transition_18202_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3570_branch_ack_1, ack => cp_elements(66)); -- 
    cp_elements(67) <= cp_elements(64);
    else_choice_transition_18206_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3570_branch_ack_0, ack => cp_elements(68)); -- 
    cp_elements(69) <= cp_elements(87);
    cp_elements(70) <= OrReduce(cp_elements(170) & cp_elements(174));
    cp_elements(71) <= cp_elements(114);
    cp_elements(72) <= OrReduce(cp_elements(117) & cp_elements(125));
    cp_elements(73) <= cp_elements(167);
    cp_elements(74) <= cp_elements(66);
    cp_elements(75) <= cp_elements(74);
    pipe_wreq_18231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => simple_obj_ref_3575_inst_req_0); -- 
    pipe_wack_18232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3575_inst_ack_0, ack => cp_elements(76)); -- 
    cp_elements(77) <= cp_elements(74);
    pipe_wreq_18243_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => simple_obj_ref_3578_inst_req_0); -- 
    pipe_wack_18244_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3578_inst_ack_0, ack => cp_elements(78)); -- 
    cp_elements(79) <= cp_elements(74);
    pipe_wreq_18254_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => simple_obj_ref_3581_inst_req_0); -- 
    pipe_wack_18255_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3581_inst_ack_0, ack => cp_elements(80)); -- 
    cp_elements(81) <= cp_elements(74);
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(83) & cp_elements(84));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18267_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => binary_3587_inst_req_0); -- 
    cp_elements(83) <= cp_elements(81);
    cp_elements(84) <= cp_elements(81);
    ra_18268_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3587_inst_ack_0, ack => cp_elements(85)); -- 
    cr_18269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(85), ack => binary_3587_inst_req_1); -- 
    ca_18270_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3587_inst_ack_1, ack => cp_elements(86)); -- 
    cpelement_group_87 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(78) & cp_elements(80) & cp_elements(86));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(87),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(88) <= cp_elements(70);
    cp_elements(89) <= cp_elements(88);
    pipe_wreq_18283_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => simple_obj_ref_3598_inst_req_0); -- 
    pipe_wack_18284_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3598_inst_ack_0, ack => cp_elements(90)); -- 
    cp_elements(91) <= cp_elements(88);
    cp_elements(92) <= cp_elements(91);
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(92) & cp_elements(103));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_18333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => array_obj_ref_3603_final_reg_req_0); -- 
    cp_elements(94) <= cp_elements(91);
    base_resize_req_18320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => array_obj_ref_3603_base_resize_req_0); -- 
    cp_elements(95) <= cp_elements(91);
    index_resize_req_18302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_3603_index_0_resize_req_0); -- 
    index_resize_ack_18303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_index_0_resize_ack_0, ack => cp_elements(96)); -- 
    scale_rr_18307_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => array_obj_ref_3603_index_0_scale_req_0); -- 
    scale_ra_18308_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_index_0_scale_ack_0, ack => cp_elements(97)); -- 
    scale_cr_18309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => array_obj_ref_3603_index_0_scale_req_1); -- 
    scale_ca_18310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_index_0_scale_ack_1, ack => cp_elements(98)); -- 
    final_index_req_18314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => array_obj_ref_3603_offset_inst_req_0); -- 
    final_index_ack_18315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_offset_inst_ack_0, ack => cp_elements(99)); -- 
    base_resize_ack_18321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_base_resize_ack_0, ack => cp_elements(100)); -- 
    cpelement_group_101 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(99) & cp_elements(100));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(101),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_18326_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(101), ack => array_obj_ref_3603_root_address_inst_req_0); -- 
    plus_base_ra_18327_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_root_address_inst_ack_0, ack => cp_elements(102)); -- 
    plus_base_cr_18328_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => array_obj_ref_3603_root_address_inst_req_1); -- 
    plus_base_ca_18329_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_root_address_inst_ack_1, ack => cp_elements(103)); -- 
    final_reg_ack_18334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3603_final_reg_ack_0, ack => cp_elements(104)); -- 
    pipe_wreq_18339_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(104), ack => simple_obj_ref_3601_inst_req_0); -- 
    pipe_wack_18340_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3601_inst_ack_0, ack => cp_elements(105)); -- 
    cp_elements(106) <= cp_elements(88);
    pipe_wreq_18350_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => simple_obj_ref_3605_inst_req_0); -- 
    pipe_wack_18351_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3605_inst_ack_0, ack => cp_elements(107)); -- 
    cp_elements(108) <= cp_elements(88);
    cpelement_group_109 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(110) & cp_elements(111));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(109),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18363_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => binary_3611_inst_req_0); -- 
    cp_elements(110) <= cp_elements(108);
    cp_elements(111) <= cp_elements(108);
    ra_18364_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3611_inst_ack_0, ack => cp_elements(112)); -- 
    cr_18365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(112), ack => binary_3611_inst_req_1); -- 
    ca_18366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3611_inst_ack_1, ack => cp_elements(113)); -- 
    cpelement_group_114 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(90) & cp_elements(105) & cp_elements(107) & cp_elements(113));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(115) <= cp_elements(71);
    cp_elements(116) <= false;
    cp_elements(117) <= cp_elements(116);
    cp_elements(118) <= cp_elements(71);
    rr_18380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => binary_3617_inst_req_0); -- 
    ra_18381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3617_inst_ack_0, ack => cp_elements(119)); -- 
    cr_18382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => binary_3617_inst_req_1); -- 
    ca_18383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3617_inst_ack_1, ack => cp_elements(120)); -- 
    branch_req_18384_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => if_stmt_3614_branch_req_0); -- 
    cp_elements(121) <= cp_elements(120);
    cp_elements(122) <= cp_elements(121);
    if_choice_transition_18389_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3614_branch_ack_1, ack => cp_elements(123)); -- 
    phi_stmt_3591_req_18549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(123), ack => phi_stmt_3591_req_1); -- 
    cp_elements(124) <= cp_elements(121);
    else_choice_transition_18393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3614_branch_ack_0, ack => cp_elements(125)); -- 
    cp_elements(126) <= cp_elements(72);
    cp_elements(127) <= cp_elements(126);
    cpelement_group_128 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(127) & cp_elements(138));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(128),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_18443_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(128), ack => array_obj_ref_3622_final_reg_req_0); -- 
    cp_elements(129) <= cp_elements(126);
    base_resize_req_18430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => array_obj_ref_3622_base_resize_req_0); -- 
    cp_elements(130) <= cp_elements(126);
    index_resize_req_18412_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(130), ack => array_obj_ref_3622_index_0_resize_req_0); -- 
    index_resize_ack_18413_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_index_0_resize_ack_0, ack => cp_elements(131)); -- 
    scale_rr_18417_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(131), ack => array_obj_ref_3622_index_0_scale_req_0); -- 
    scale_ra_18418_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_index_0_scale_ack_0, ack => cp_elements(132)); -- 
    scale_cr_18419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(132), ack => array_obj_ref_3622_index_0_scale_req_1); -- 
    scale_ca_18420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_index_0_scale_ack_1, ack => cp_elements(133)); -- 
    final_index_req_18424_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(133), ack => array_obj_ref_3622_offset_inst_req_0); -- 
    final_index_ack_18425_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_offset_inst_ack_0, ack => cp_elements(134)); -- 
    base_resize_ack_18431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_base_resize_ack_0, ack => cp_elements(135)); -- 
    cpelement_group_136 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(134) & cp_elements(135));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(136),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    plus_base_rr_18436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => array_obj_ref_3622_root_address_inst_req_0); -- 
    plus_base_ra_18437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_root_address_inst_ack_0, ack => cp_elements(137)); -- 
    plus_base_cr_18438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(137), ack => array_obj_ref_3622_root_address_inst_req_1); -- 
    plus_base_ca_18439_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_root_address_inst_ack_1, ack => cp_elements(138)); -- 
    final_reg_ack_18444_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_3622_final_reg_ack_0, ack => cp_elements(139)); -- 
    cp_elements(140) <= cp_elements(139);
    cp_elements(141) <= cp_elements(140);
    cpelement_group_142 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(143) & cp_elements(159));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(142),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => binary_3636_inst_req_0); -- 
    cp_elements(143) <= cp_elements(141);
    cpelement_group_144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(145) & cp_elements(158));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => type_cast_3635_inst_req_0); -- 
    cp_elements(145) <= cp_elements(141);
    cpelement_group_146 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(147) & cp_elements(156));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(146),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18481_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(146), ack => binary_3634_inst_req_0); -- 
    cp_elements(147) <= cp_elements(141);
    cpelement_group_148 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(149) & cp_elements(154));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(148),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(148), ack => binary_3632_inst_req_0); -- 
    cp_elements(149) <= cp_elements(141);
    cpelement_group_150 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(151) & cp_elements(152));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(150),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(150), ack => binary_3631_inst_req_0); -- 
    cp_elements(151) <= cp_elements(141);
    cp_elements(152) <= cp_elements(141);
    ra_18468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3631_inst_ack_0, ack => cp_elements(153)); -- 
    cr_18469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(153), ack => binary_3631_inst_req_1); -- 
    ca_18470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3631_inst_ack_1, ack => cp_elements(154)); -- 
    ra_18475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3632_inst_ack_0, ack => cp_elements(155)); -- 
    cr_18476_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(155), ack => binary_3632_inst_req_1); -- 
    ca_18477_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3632_inst_ack_1, ack => cp_elements(156)); -- 
    ra_18482_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3634_inst_ack_0, ack => cp_elements(157)); -- 
    cr_18483_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(157), ack => binary_3634_inst_req_1); -- 
    ca_18484_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3634_inst_ack_1, ack => cp_elements(158)); -- 
    ack_18489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3635_inst_ack_0, ack => cp_elements(159)); -- 
    ra_18494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3636_inst_ack_0, ack => cp_elements(160)); -- 
    cr_18495_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => binary_3636_inst_req_1); -- 
    ca_18496_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3636_inst_ack_1, ack => cp_elements(161)); -- 
    pipe_wreq_18501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(161), ack => simple_obj_ref_3625_inst_req_0); -- 
    pipe_wack_18502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3625_inst_ack_0, ack => cp_elements(162)); -- 
    cp_elements(163) <= cp_elements(140);
    pipe_wreq_18513_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(163), ack => simple_obj_ref_3638_inst_req_0); -- 
    pipe_wack_18514_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3638_inst_ack_0, ack => cp_elements(164)); -- 
    cp_elements(165) <= cp_elements(140);
    pipe_wreq_18524_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(165), ack => simple_obj_ref_3641_inst_req_0); -- 
    pipe_wack_18525_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3641_inst_ack_0, ack => cp_elements(166)); -- 
    cpelement_group_167 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(162) & cp_elements(164) & cp_elements(166));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(167),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(168) <= cp_elements(69);
    cp_elements(169) <= false;
    cp_elements(170) <= cp_elements(169);
    cp_elements(171) <= cp_elements(69);
    phi_stmt_3591_req_18539_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => phi_stmt_3591_req_0); -- 
    cp_elements(172) <= OrReduce(cp_elements(123) & cp_elements(171));
    cp_elements(173) <= cp_elements(172);
    phi_stmt_3591_ack_18554_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3591_ack_0, ack => cp_elements(174)); -- 
    cp_elements(175) <= cp_elements(43);
    cp_elements(176) <= false;
    cp_elements(177) <= cp_elements(176);
    cp_elements(178) <= cp_elements(43);
    cp_elements(179) <= OrReduce(cp_elements(47) & cp_elements(178));
    cp_elements(180) <= cp_elements(179);
    cp_elements(181) <= cp_elements(0);
    cp_elements(182) <= false; 
    cp_elements(183) <= OrReduce(cp_elements(260) & cp_elements(263));
    cp_elements(184) <= cp_elements(257);
    cp_elements(185) <= cp_elements(183);
    cp_elements(186) <= cp_elements(185);
    req_18595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(186), ack => simple_obj_ref_3652_inst_req_0); -- 
    ack_18596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3652_inst_ack_0, ack => cp_elements(187)); -- 
    base_resize_req_18603_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => ptr_deref_3653_base_resize_req_0); -- 
    base_resize_ack_18604_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_base_resize_ack_0, ack => cp_elements(188)); -- 
    sum_rename_req_18608_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(188), ack => ptr_deref_3653_root_address_inst_req_0); -- 
    cp_elements(189) <= ptr_deref_3653_root_address_inst_ack_0;
    cp_elements(190) <= cp_elements(189);
    rr_18616_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(190), ack => ptr_deref_3653_addr_0_req_0); -- 
    ra_18617_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_0_ack_0, ack => cp_elements(191)); -- 
    cr_18618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => ptr_deref_3653_addr_0_req_1); -- 
    ca_18619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_0_ack_1, ack => cp_elements(192)); -- 
    cp_elements(193) <= cp_elements(189);
    rr_18623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(193), ack => ptr_deref_3653_addr_1_req_0); -- 
    ra_18624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_1_ack_0, ack => cp_elements(194)); -- 
    cr_18625_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(194), ack => ptr_deref_3653_addr_1_req_1); -- 
    ca_18626_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_1_ack_1, ack => cp_elements(195)); -- 
    cp_elements(196) <= cp_elements(189);
    rr_18630_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(196), ack => ptr_deref_3653_addr_2_req_0); -- 
    ra_18631_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_2_ack_0, ack => cp_elements(197)); -- 
    cr_18632_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(197), ack => ptr_deref_3653_addr_2_req_1); -- 
    ca_18633_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_2_ack_1, ack => cp_elements(198)); -- 
    cp_elements(199) <= cp_elements(189);
    rr_18637_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(199), ack => ptr_deref_3653_addr_3_req_0); -- 
    ra_18638_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_3_ack_0, ack => cp_elements(200)); -- 
    cr_18639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(200), ack => ptr_deref_3653_addr_3_req_1); -- 
    ca_18640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_3_ack_1, ack => cp_elements(201)); -- 
    cp_elements(202) <= cp_elements(189);
    rr_18644_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(202), ack => ptr_deref_3653_addr_4_req_0); -- 
    ra_18645_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_4_ack_0, ack => cp_elements(203)); -- 
    cr_18646_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => ptr_deref_3653_addr_4_req_1); -- 
    ca_18647_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_4_ack_1, ack => cp_elements(204)); -- 
    cp_elements(205) <= cp_elements(189);
    rr_18651_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => ptr_deref_3653_addr_5_req_0); -- 
    ra_18652_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_5_ack_0, ack => cp_elements(206)); -- 
    cr_18653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(206), ack => ptr_deref_3653_addr_5_req_1); -- 
    ca_18654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_5_ack_1, ack => cp_elements(207)); -- 
    cp_elements(208) <= cp_elements(189);
    rr_18658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(208), ack => ptr_deref_3653_addr_6_req_0); -- 
    ra_18659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_6_ack_0, ack => cp_elements(209)); -- 
    cr_18660_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => ptr_deref_3653_addr_6_req_1); -- 
    ca_18661_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_6_ack_1, ack => cp_elements(210)); -- 
    cp_elements(211) <= cp_elements(189);
    rr_18665_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(211), ack => ptr_deref_3653_addr_7_req_0); -- 
    ra_18666_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_7_ack_0, ack => cp_elements(212)); -- 
    cr_18667_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(212), ack => ptr_deref_3653_addr_7_req_1); -- 
    ca_18668_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_addr_7_ack_1, ack => cp_elements(213)); -- 
    cpelement_group_214 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(192) & cp_elements(195) & cp_elements(198) & cp_elements(201) & cp_elements(204) & cp_elements(207) & cp_elements(210) & cp_elements(213));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(214),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(215) <= cp_elements(214);
    rr_18678_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(215), ack => ptr_deref_3653_load_0_req_0); -- 
    ra_18679_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_0_ack_0, ack => cp_elements(216)); -- 
    cp_elements(217) <= cp_elements(214);
    rr_18683_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(217), ack => ptr_deref_3653_load_1_req_0); -- 
    ra_18684_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_1_ack_0, ack => cp_elements(218)); -- 
    cp_elements(219) <= cp_elements(214);
    rr_18688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => ptr_deref_3653_load_2_req_0); -- 
    ra_18689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_2_ack_0, ack => cp_elements(220)); -- 
    cp_elements(221) <= cp_elements(214);
    rr_18693_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => ptr_deref_3653_load_3_req_0); -- 
    ra_18694_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_3_ack_0, ack => cp_elements(222)); -- 
    cp_elements(223) <= cp_elements(214);
    rr_18698_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => ptr_deref_3653_load_4_req_0); -- 
    ra_18699_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_4_ack_0, ack => cp_elements(224)); -- 
    cp_elements(225) <= cp_elements(214);
    rr_18703_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => ptr_deref_3653_load_5_req_0); -- 
    ra_18704_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_5_ack_0, ack => cp_elements(226)); -- 
    cp_elements(227) <= cp_elements(214);
    rr_18708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => ptr_deref_3653_load_6_req_0); -- 
    ra_18709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_6_ack_0, ack => cp_elements(228)); -- 
    cp_elements(229) <= cp_elements(214);
    rr_18713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(229), ack => ptr_deref_3653_load_7_req_0); -- 
    ra_18714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_7_ack_0, ack => cp_elements(230)); -- 
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(216) & cp_elements(218) & cp_elements(220) & cp_elements(222) & cp_elements(224) & cp_elements(226) & cp_elements(228) & cp_elements(230));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(232) <= cp_elements(231);
    cr_18724_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(232), ack => ptr_deref_3653_load_0_req_1); -- 
    ca_18725_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_0_ack_1, ack => cp_elements(233)); -- 
    cp_elements(234) <= cp_elements(231);
    cr_18729_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(234), ack => ptr_deref_3653_load_1_req_1); -- 
    ca_18730_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_1_ack_1, ack => cp_elements(235)); -- 
    cp_elements(236) <= cp_elements(231);
    cr_18734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => ptr_deref_3653_load_2_req_1); -- 
    ca_18735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_2_ack_1, ack => cp_elements(237)); -- 
    cp_elements(238) <= cp_elements(231);
    cr_18739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => ptr_deref_3653_load_3_req_1); -- 
    ca_18740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_3_ack_1, ack => cp_elements(239)); -- 
    cp_elements(240) <= cp_elements(231);
    cr_18744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(240), ack => ptr_deref_3653_load_4_req_1); -- 
    ca_18745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_4_ack_1, ack => cp_elements(241)); -- 
    cp_elements(242) <= cp_elements(231);
    cr_18749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(242), ack => ptr_deref_3653_load_5_req_1); -- 
    ca_18750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_5_ack_1, ack => cp_elements(243)); -- 
    cp_elements(244) <= cp_elements(231);
    cr_18754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(244), ack => ptr_deref_3653_load_6_req_1); -- 
    ca_18755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_6_ack_1, ack => cp_elements(245)); -- 
    cp_elements(246) <= cp_elements(231);
    cr_18759_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(246), ack => ptr_deref_3653_load_7_req_1); -- 
    ca_18760_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_load_7_ack_1, ack => cp_elements(247)); -- 
    cpelement_group_248 : Block -- 
      signal predecessors: BooleanArray(7 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(233) & cp_elements(235) & cp_elements(237) & cp_elements(239) & cp_elements(241) & cp_elements(243) & cp_elements(245) & cp_elements(247));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(248),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    merge_req_18761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => ptr_deref_3653_gather_scatter_req_0); -- 
    merge_ack_18762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3653_gather_scatter_ack_0, ack => cp_elements(249)); -- 
    pipe_wreq_18767_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(249), ack => simple_obj_ref_3651_inst_req_0); -- 
    pipe_wack_18768_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3651_inst_ack_0, ack => cp_elements(250)); -- 
    cp_elements(251) <= cp_elements(185);
    req_18778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(251), ack => simple_obj_ref_3656_inst_req_0); -- 
    ack_18779_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3656_inst_ack_0, ack => cp_elements(252)); -- 
    pipe_wreq_18784_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => simple_obj_ref_3655_inst_req_0); -- 
    pipe_wack_18785_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3655_inst_ack_0, ack => cp_elements(253)); -- 
    cp_elements(254) <= cp_elements(185);
    req_18795_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => simple_obj_ref_3659_inst_req_0); -- 
    ack_18796_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3659_inst_ack_0, ack => cp_elements(255)); -- 
    pipe_wreq_18801_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(255), ack => simple_obj_ref_3658_inst_req_0); -- 
    pipe_wack_18802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3658_inst_ack_0, ack => cp_elements(256)); -- 
    cpelement_group_257 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(250) & cp_elements(253) & cp_elements(256));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(257),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(258) <= cp_elements(181);
    cp_elements(259) <= false;
    cp_elements(260) <= cp_elements(259);
    cp_elements(261) <= cp_elements(181);
    cp_elements(262) <= OrReduce(cp_elements(184) & cp_elements(261));
    cp_elements(263) <= cp_elements(262);
    cp_elements(264) <= cp_elements(0);
    cp_elements(265) <= false; 
    cp_elements(266) <= OrReduce(cp_elements(369) & cp_elements(372));
    req_18839_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => simple_obj_ref_3667_inst_req_0); -- 
    cp_elements(267) <= cp_elements(366);
    ack_18840_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3667_inst_ack_0, ack => cp_elements(268)); -- 
    cp_elements(269) <= cp_elements(268);
    cp_elements(270) <= cp_elements(269);
    cpelement_group_271 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(272) & cp_elements(312) & cp_elements(356));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(271),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19035_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(271), ack => binary_3707_inst_req_0); -- 
    cp_elements(272) <= cp_elements(270);
    cpelement_group_273 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(274) & cp_elements(290) & cp_elements(310));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(273),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(273), ack => binary_3687_inst_req_0); -- 
    cp_elements(274) <= cp_elements(270);
    cpelement_group_275 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(276) & cp_elements(280) & cp_elements(288));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(275),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(275), ack => binary_3677_inst_req_0); -- 
    cp_elements(276) <= cp_elements(270);
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(278) & cp_elements(279));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(277), ack => type_cast_3672_inst_req_0); -- 
    cp_elements(278) <= cp_elements(270);
    cp_elements(279) <= cp_elements(270);
    ack_18862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3672_inst_ack_0, ack => cp_elements(280)); -- 
    cpelement_group_281 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(282) & cp_elements(287));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(281),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18878_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(281), ack => type_cast_3676_inst_req_0); -- 
    cp_elements(282) <= cp_elements(270);
    cpelement_group_283 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(284) & cp_elements(285));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(283),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18871_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(283), ack => binary_3675_inst_req_0); -- 
    cp_elements(284) <= cp_elements(270);
    cp_elements(285) <= cp_elements(270);
    ra_18872_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3675_inst_ack_0, ack => cp_elements(286)); -- 
    cr_18873_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => binary_3675_inst_req_1); -- 
    ca_18874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3675_inst_ack_1, ack => cp_elements(287)); -- 
    ack_18879_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3676_inst_ack_0, ack => cp_elements(288)); -- 
    ra_18884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3677_inst_ack_0, ack => cp_elements(289)); -- 
    cr_18885_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(289), ack => binary_3677_inst_req_1); -- 
    ca_18886_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3677_inst_ack_1, ack => cp_elements(290)); -- 
    cpelement_group_291 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(292) & cp_elements(300) & cp_elements(308));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(291),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(291), ack => binary_3686_inst_req_0); -- 
    cp_elements(292) <= cp_elements(270);
    cpelement_group_293 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(294) & cp_elements(299));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(293),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18904_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(293), ack => type_cast_3681_inst_req_0); -- 
    cp_elements(294) <= cp_elements(270);
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(296) & cp_elements(297));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18897_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(295), ack => binary_3680_inst_req_0); -- 
    cp_elements(296) <= cp_elements(270);
    cp_elements(297) <= cp_elements(270);
    ra_18898_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3680_inst_ack_0, ack => cp_elements(298)); -- 
    cr_18899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(298), ack => binary_3680_inst_req_1); -- 
    ca_18900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3680_inst_ack_1, ack => cp_elements(299)); -- 
    ack_18905_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3681_inst_ack_0, ack => cp_elements(300)); -- 
    cpelement_group_301 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(302) & cp_elements(307));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(301),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => type_cast_3685_inst_req_0); -- 
    cp_elements(302) <= cp_elements(270);
    cpelement_group_303 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(304) & cp_elements(305));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(303),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18914_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(303), ack => binary_3684_inst_req_0); -- 
    cp_elements(304) <= cp_elements(270);
    cp_elements(305) <= cp_elements(270);
    ra_18915_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3684_inst_ack_0, ack => cp_elements(306)); -- 
    cr_18916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(306), ack => binary_3684_inst_req_1); -- 
    ca_18917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3684_inst_ack_1, ack => cp_elements(307)); -- 
    ack_18922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3685_inst_ack_0, ack => cp_elements(308)); -- 
    ra_18927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3686_inst_ack_0, ack => cp_elements(309)); -- 
    cr_18928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(309), ack => binary_3686_inst_req_1); -- 
    ca_18929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3686_inst_ack_1, ack => cp_elements(310)); -- 
    ra_18934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3687_inst_ack_0, ack => cp_elements(311)); -- 
    cr_18935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(311), ack => binary_3687_inst_req_1); -- 
    ca_18936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3687_inst_ack_1, ack => cp_elements(312)); -- 
    cpelement_group_313 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(314) & cp_elements(334) & cp_elements(354));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(313),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19028_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => binary_3706_inst_req_0); -- 
    cp_elements(314) <= cp_elements(270);
    cpelement_group_315 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(316) & cp_elements(324) & cp_elements(332));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(315),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18978_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => binary_3696_inst_req_0); -- 
    cp_elements(316) <= cp_elements(270);
    cpelement_group_317 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(318) & cp_elements(323));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(317),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(317), ack => type_cast_3691_inst_req_0); -- 
    cp_elements(318) <= cp_elements(270);
    cpelement_group_319 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(320) & cp_elements(321));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(319),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18949_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => binary_3690_inst_req_0); -- 
    cp_elements(320) <= cp_elements(270);
    cp_elements(321) <= cp_elements(270);
    ra_18950_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3690_inst_ack_0, ack => cp_elements(322)); -- 
    cr_18951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(322), ack => binary_3690_inst_req_1); -- 
    ca_18952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3690_inst_ack_1, ack => cp_elements(323)); -- 
    ack_18957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3691_inst_ack_0, ack => cp_elements(324)); -- 
    cpelement_group_325 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(326) & cp_elements(331));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(325),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18973_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(325), ack => type_cast_3695_inst_req_0); -- 
    cp_elements(326) <= cp_elements(270);
    cpelement_group_327 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(328) & cp_elements(329));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(327),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18966_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(327), ack => binary_3694_inst_req_0); -- 
    cp_elements(328) <= cp_elements(270);
    cp_elements(329) <= cp_elements(270);
    ra_18967_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3694_inst_ack_0, ack => cp_elements(330)); -- 
    cr_18968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(330), ack => binary_3694_inst_req_1); -- 
    ca_18969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3694_inst_ack_1, ack => cp_elements(331)); -- 
    ack_18974_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3695_inst_ack_0, ack => cp_elements(332)); -- 
    ra_18979_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3696_inst_ack_0, ack => cp_elements(333)); -- 
    cr_18980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => binary_3696_inst_req_1); -- 
    ca_18981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3696_inst_ack_1, ack => cp_elements(334)); -- 
    cpelement_group_335 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(336) & cp_elements(344) & cp_elements(352));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(335),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19021_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => binary_3705_inst_req_0); -- 
    cp_elements(336) <= cp_elements(270);
    cpelement_group_337 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(338) & cp_elements(343));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(337),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_18999_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(337), ack => type_cast_3700_inst_req_0); -- 
    cp_elements(338) <= cp_elements(270);
    cpelement_group_339 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(340) & cp_elements(341));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(339),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_18992_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => binary_3699_inst_req_0); -- 
    cp_elements(340) <= cp_elements(270);
    cp_elements(341) <= cp_elements(270);
    ra_18993_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3699_inst_ack_0, ack => cp_elements(342)); -- 
    cr_18994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(342), ack => binary_3699_inst_req_1); -- 
    ca_18995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3699_inst_ack_1, ack => cp_elements(343)); -- 
    ack_19000_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3700_inst_ack_0, ack => cp_elements(344)); -- 
    cpelement_group_345 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(346) & cp_elements(351));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(345),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19016_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(345), ack => type_cast_3704_inst_req_0); -- 
    cp_elements(346) <= cp_elements(270);
    cpelement_group_347 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(348) & cp_elements(349));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(347),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19009_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(347), ack => binary_3703_inst_req_0); -- 
    cp_elements(348) <= cp_elements(270);
    cp_elements(349) <= cp_elements(270);
    ra_19010_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3703_inst_ack_0, ack => cp_elements(350)); -- 
    cr_19011_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(350), ack => binary_3703_inst_req_1); -- 
    ca_19012_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3703_inst_ack_1, ack => cp_elements(351)); -- 
    ack_19017_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3704_inst_ack_0, ack => cp_elements(352)); -- 
    ra_19022_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3705_inst_ack_0, ack => cp_elements(353)); -- 
    cr_19023_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => binary_3705_inst_req_1); -- 
    ca_19024_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3705_inst_ack_1, ack => cp_elements(354)); -- 
    ra_19029_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3706_inst_ack_0, ack => cp_elements(355)); -- 
    cr_19030_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(355), ack => binary_3706_inst_req_1); -- 
    ca_19031_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3706_inst_ack_1, ack => cp_elements(356)); -- 
    ra_19036_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3707_inst_ack_0, ack => cp_elements(357)); -- 
    cr_19037_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => binary_3707_inst_req_1); -- 
    ca_19038_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3707_inst_ack_1, ack => cp_elements(358)); -- 
    pipe_wreq_19043_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(358), ack => simple_obj_ref_3670_inst_req_0); -- 
    pipe_wack_19044_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3670_inst_ack_0, ack => cp_elements(359)); -- 
    cp_elements(360) <= cp_elements(269);
    req_19054_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(360), ack => simple_obj_ref_3710_inst_req_0); -- 
    ack_19055_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3710_inst_ack_0, ack => cp_elements(361)); -- 
    pipe_wreq_19060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(361), ack => simple_obj_ref_3709_inst_req_0); -- 
    pipe_wack_19061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3709_inst_ack_0, ack => cp_elements(362)); -- 
    cp_elements(363) <= cp_elements(269);
    req_19071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(363), ack => simple_obj_ref_3713_inst_req_0); -- 
    ack_19072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3713_inst_ack_0, ack => cp_elements(364)); -- 
    pipe_wreq_19077_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(364), ack => simple_obj_ref_3712_inst_req_0); -- 
    pipe_wack_19078_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3712_inst_ack_0, ack => cp_elements(365)); -- 
    cpelement_group_366 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(359) & cp_elements(362) & cp_elements(365));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(366),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(367) <= cp_elements(264);
    cp_elements(368) <= false;
    cp_elements(369) <= cp_elements(368);
    cp_elements(370) <= cp_elements(264);
    cp_elements(371) <= OrReduce(cp_elements(267) & cp_elements(370));
    cp_elements(372) <= cp_elements(371);
    cp_elements(373) <= cp_elements(0);
    cp_elements(374) <= false; 
    cp_elements(375) <= OrReduce(cp_elements(398) & cp_elements(401));
    cp_elements(376) <= OrReduce(cp_elements(379) & cp_elements(388) & cp_elements(395));
    cp_elements(377) <= cp_elements(375);
    cp_elements(378) <= false;
    cp_elements(379) <= cp_elements(378);
    cp_elements(380) <= cp_elements(375);
    req_19120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => simple_obj_ref_3721_inst_req_0); -- 
    ack_19121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3721_inst_ack_0, ack => cp_elements(381)); -- 
    rr_19122_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(381), ack => binary_3723_inst_req_0); -- 
    ra_19123_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3723_inst_ack_0, ack => cp_elements(382)); -- 
    cr_19124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(382), ack => binary_3723_inst_req_1); -- 
    ca_19125_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3723_inst_ack_1, ack => cp_elements(383)); -- 
    branch_req_19126_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(383), ack => if_stmt_3720_branch_req_0); -- 
    cp_elements(384) <= cp_elements(383);
    cp_elements(385) <= cp_elements(384);
    cp_elements(386) <= if_stmt_3720_branch_ack_1;
    cp_elements(387) <= cp_elements(384);
    else_choice_transition_19135_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3720_branch_ack_0, ack => cp_elements(388)); -- 
    cpelement_group_389 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(390) & cp_elements(392));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19157_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(389), ack => binary_3728_inst_req_0); -- 
    cp_elements(390) <= cp_elements(386);
    cp_elements(391) <= cp_elements(386);
    req_19152_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(391), ack => simple_obj_ref_3726_inst_req_0); -- 
    ack_19153_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3726_inst_ack_0, ack => cp_elements(392)); -- 
    ra_19158_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3728_inst_ack_0, ack => cp_elements(393)); -- 
    cr_19159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(393), ack => binary_3728_inst_req_1); -- 
    ca_19160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_3728_inst_ack_1, ack => cp_elements(394)); -- 
    pipe_wreq_19165_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(394), ack => simple_obj_ref_3725_inst_req_0); -- 
    pipe_wack_19166_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3725_inst_ack_0, ack => cp_elements(395)); -- 
    cp_elements(396) <= cp_elements(373);
    cp_elements(397) <= false;
    cp_elements(398) <= cp_elements(397);
    cp_elements(399) <= cp_elements(373);
    cp_elements(400) <= OrReduce(cp_elements(376) & cp_elements(399));
    cp_elements(401) <= cp_elements(400);
    cpelement_group_402 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(2) & cp_elements(44) & cp_elements(182) & cp_elements(265) & cp_elements(374));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(402),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal I_3591 : std_logic_vector(15 downto 0);
    signal LI_3588 : std_logic_vector(15 downto 0);
    signal NI_3612 : std_logic_vector(15 downto 0);
    signal a_3668 : std_logic_vector(63 downto 0);
    signal array_obj_ref_3603_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3603_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3603_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3603_root_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3603_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_3622_final_offset : std_logic_vector(15 downto 0);
    signal array_obj_ref_3622_offset_scale_factor_0 : std_logic_vector(15 downto 0);
    signal array_obj_ref_3622_resized_base_address : std_logic_vector(15 downto 0);
    signal array_obj_ref_3622_root_address : std_logic_vector(15 downto 0);
    signal binary_3573_wire : std_logic_vector(0 downto 0);
    signal binary_3617_wire : std_logic_vector(0 downto 0);
    signal binary_3631_wire : std_logic_vector(15 downto 0);
    signal binary_3632_wire : std_logic_vector(15 downto 0);
    signal binary_3634_wire : std_logic_vector(15 downto 0);
    signal binary_3636_wire : std_logic_vector(7 downto 0);
    signal binary_3675_wire : std_logic_vector(63 downto 0);
    signal binary_3677_wire : std_logic_vector(15 downto 0);
    signal binary_3680_wire : std_logic_vector(63 downto 0);
    signal binary_3684_wire : std_logic_vector(63 downto 0);
    signal binary_3686_wire : std_logic_vector(15 downto 0);
    signal binary_3687_wire : std_logic_vector(31 downto 0);
    signal binary_3690_wire : std_logic_vector(63 downto 0);
    signal binary_3694_wire : std_logic_vector(63 downto 0);
    signal binary_3696_wire : std_logic_vector(15 downto 0);
    signal binary_3699_wire : std_logic_vector(63 downto 0);
    signal binary_3703_wire : std_logic_vector(63 downto 0);
    signal binary_3705_wire : std_logic_vector(15 downto 0);
    signal binary_3706_wire : std_logic_vector(31 downto 0);
    signal binary_3707_wire : std_logic_vector(63 downto 0);
    signal binary_3723_wire : std_logic_vector(0 downto 0);
    signal binary_3728_wire : std_logic_vector(31 downto 0);
    signal blen_3531 : std_logic_vector(15 downto 0);
    signal blen_3562 : std_logic_vector(15 downto 0);
    signal buf64_3565 : std_logic_vector(31 downto 0);
    signal buf_3531 : std_logic_vector(31 downto 0);
    signal expr_3572_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3576_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3582_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3586_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3599_wire_constant : std_logic_vector(7 downto 0);
    signal expr_3606_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3610_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3628_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3630_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3633_wire_constant : std_logic_vector(15 downto 0);
    signal expr_3642_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3674_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3679_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3683_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3689_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3693_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3698_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3702_wire_constant : std_logic_vector(63 downto 0);
    signal expr_3722_wire_constant : std_logic_vector(0 downto 0);
    signal expr_3727_wire_constant : std_logic_vector(31 downto 0);
    signal last_word_ptr_3623 : std_logic_vector(31 downto 0);
    signal pkt64_3568 : std_logic_vector(31 downto 0);
    signal pkt_3525 : std_logic_vector(31 downto 0);
    signal ptr_deref_3653_data_0 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_1 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_2 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_3 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_4 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_5 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_6 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_data_7 : std_logic_vector(7 downto 0);
    signal ptr_deref_3653_resized_base_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_root_address : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_wire : std_logic_vector(63 downto 0);
    signal ptr_deref_3653_word_address_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_address_7 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_0 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_1 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_2 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_3 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_4 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_5 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_6 : std_logic_vector(15 downto 0);
    signal ptr_deref_3653_word_offset_7 : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3602_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3602_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3621_resized : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3621_scaled : std_logic_vector(15 downto 0);
    signal simple_obj_ref_3652_wire : std_logic_vector(31 downto 0);
    signal simple_obj_ref_3656_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_3659_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3710_wire : std_logic_vector(7 downto 0);
    signal simple_obj_ref_3713_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3721_wire : std_logic_vector(0 downto 0);
    signal simple_obj_ref_3726_wire : std_logic_vector(31 downto 0);
    signal type_cast_3527_wire : std_logic_vector(31 downto 0);
    signal type_cast_3535_wire : std_logic_vector(31 downto 0);
    signal type_cast_3539_wire : std_logic_vector(31 downto 0);
    signal type_cast_3549_wire : std_logic_vector(31 downto 0);
    signal type_cast_3594_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_3627_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3635_wire : std_logic_vector(7 downto 0);
    signal type_cast_3672_wire : std_logic_vector(7 downto 0);
    signal type_cast_3676_wire : std_logic_vector(7 downto 0);
    signal type_cast_3681_wire : std_logic_vector(7 downto 0);
    signal type_cast_3685_wire : std_logic_vector(7 downto 0);
    signal type_cast_3691_wire : std_logic_vector(7 downto 0);
    signal type_cast_3695_wire : std_logic_vector(7 downto 0);
    signal type_cast_3700_wire : std_logic_vector(7 downto 0);
    signal type_cast_3704_wire : std_logic_vector(7 downto 0);
    signal wlen_3531 : std_logic_vector(15 downto 0);
    signal wlen_3559 : std_logic_vector(15 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxblen_pipe
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxblen_pipe
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxblen_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxbuf64_pipe
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxbuf64_pipe
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxfree_packet_in
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxfree_packet_in
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxfree_packet_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxpkt64_pipe
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxpkt64_pipe
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_ctrl_in
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_ctrl_in
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_last_word_in
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_last_word_in
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxread_pointer
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxread_pointer
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_data: std_logic_vector(31 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxread_pointer_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_ctrl_in
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_ctrl_in
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data: std_logic_vector(7 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_data_in
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_data: std_logic_vector(63 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_data_in
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_data: std_logic_vector(63 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_data_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxswap_last_word_in
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxswap_last_word_in
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for write to pipe xxsend_packet_pipelinexxwlen_pipe
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
    -- aggregate signals for read from pipe xxsend_packet_pipelinexxwlen_pipe
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_data: std_logic_vector(15 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_req: std_logic_vector(0 downto 0);
    signal xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_3603_offset_scale_factor_0 <= "0000000000001000";
    array_obj_ref_3622_offset_scale_factor_0 <= "0000000000001000";
    expr_3572_wire_constant <= "0000000000000000";
    expr_3576_wire_constant <= "11111111";
    expr_3582_wire_constant <= "0";
    expr_3586_wire_constant <= "0000000000000001";
    expr_3599_wire_constant <= "00000000";
    expr_3606_wire_constant <= "0";
    expr_3610_wire_constant <= "0000000000000001";
    expr_3628_wire_constant <= "0000000000001000";
    expr_3630_wire_constant <= "0000000000000111";
    expr_3633_wire_constant <= "0000000000000111";
    expr_3642_wire_constant <= "1";
    expr_3674_wire_constant <= "0000000000000000000000000000000000000000000000000000000000001000";
    expr_3679_wire_constant <= "0000000000000000000000000000000000000000000000000000000000010000";
    expr_3683_wire_constant <= "0000000000000000000000000000000000000000000000000000000000011000";
    expr_3689_wire_constant <= "0000000000000000000000000000000000000000000000000000000000100000";
    expr_3693_wire_constant <= "0000000000000000000000000000000000000000000000000000000000101000";
    expr_3698_wire_constant <= "0000000000000000000000000000000000000000000000000000000000110000";
    expr_3702_wire_constant <= "0000000000000000000000000000000000000000000000000000000000111000";
    expr_3722_wire_constant <= "0";
    expr_3727_wire_constant <= "11111111111111111111100000000000";
    ptr_deref_3653_word_offset_0 <= "0000000000000000";
    ptr_deref_3653_word_offset_1 <= "0000000000000001";
    ptr_deref_3653_word_offset_2 <= "0000000000000010";
    ptr_deref_3653_word_offset_3 <= "0000000000000011";
    ptr_deref_3653_word_offset_4 <= "0000000000000100";
    ptr_deref_3653_word_offset_5 <= "0000000000000101";
    ptr_deref_3653_word_offset_6 <= "0000000000000110";
    ptr_deref_3653_word_offset_7 <= "0000000000000111";
    type_cast_3594_wire_constant <= "0000000000000000";
    type_cast_3627_wire_constant <= "00000001";
    phi_stmt_3591: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3594_wire_constant & NI_3612;
      req <= phi_stmt_3591_req_0 & phi_stmt_3591_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 16) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3591_ack_0,
          idata => idata,
          odata => I_3591,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3591
    array_obj_ref_3603_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_3568, dout => array_obj_ref_3603_resized_base_address, req => array_obj_ref_3603_base_resize_req_0, ack => array_obj_ref_3603_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3603_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3603_root_address, dout => array_obj_ref_3603_wire, req => array_obj_ref_3603_final_reg_req_0, ack => array_obj_ref_3603_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3603_index_0_resize: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => I_3591, dout => simple_obj_ref_3602_resized, req => array_obj_ref_3603_index_0_resize_req_0, ack => array_obj_ref_3603_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3603_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3602_scaled, dout => array_obj_ref_3603_final_offset, req => array_obj_ref_3603_offset_inst_req_0, ack => array_obj_ref_3603_offset_inst_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3622_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => pkt64_3568, dout => array_obj_ref_3622_resized_base_address, req => array_obj_ref_3622_base_resize_req_0, ack => array_obj_ref_3622_base_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3622_final_reg: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 32, flow_through => false ) 
      port map( din => array_obj_ref_3622_root_address, dout => last_word_ptr_3623, req => array_obj_ref_3622_final_reg_req_0, ack => array_obj_ref_3622_final_reg_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3622_index_0_resize: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => LI_3588, dout => simple_obj_ref_3621_resized, req => array_obj_ref_3622_index_0_resize_req_0, ack => array_obj_ref_3622_index_0_resize_ack_0, clk => clk, reset => reset); -- 
    array_obj_ref_3622_offset_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3621_scaled, dout => array_obj_ref_3622_final_offset, req => array_obj_ref_3622_offset_inst_req_0, ack => array_obj_ref_3622_offset_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3653_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 16, flow_through => true ) 
      port map( din => simple_obj_ref_3652_wire, dout => ptr_deref_3653_resized_base_address, req => ptr_deref_3653_base_resize_req_0, ack => ptr_deref_3653_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_3527_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_3525, dout => type_cast_3527_wire, req => type_cast_3527_inst_req_0, ack => type_cast_3527_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3535_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => buf_3531, dout => type_cast_3535_wire, req => type_cast_3535_inst_req_0, ack => type_cast_3535_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3539_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_3525, dout => type_cast_3539_wire, req => type_cast_3539_inst_req_0, ack => type_cast_3539_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3549_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => true ) 
      port map( din => pkt_3525, dout => type_cast_3549_wire, req => type_cast_3549_inst_req_0, ack => type_cast_3549_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3635_inst: RegisterBase --
      generic map(in_data_width => 16,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3634_wire, dout => type_cast_3635_wire, req => type_cast_3635_inst_req_0, ack => type_cast_3635_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3672_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => a_3668, dout => type_cast_3672_wire, req => type_cast_3672_inst_req_0, ack => type_cast_3672_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3676_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3675_wire, dout => type_cast_3676_wire, req => type_cast_3676_inst_req_0, ack => type_cast_3676_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3681_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3680_wire, dout => type_cast_3681_wire, req => type_cast_3681_inst_req_0, ack => type_cast_3681_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3685_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3684_wire, dout => type_cast_3685_wire, req => type_cast_3685_inst_req_0, ack => type_cast_3685_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3691_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3690_wire, dout => type_cast_3691_wire, req => type_cast_3691_inst_req_0, ack => type_cast_3691_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3695_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3694_wire, dout => type_cast_3695_wire, req => type_cast_3695_inst_req_0, ack => type_cast_3695_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3700_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3699_wire, dout => type_cast_3700_wire, req => type_cast_3700_inst_req_0, ack => type_cast_3700_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3704_inst: RegisterBase --
      generic map(in_data_width => 64,out_data_width => 8, flow_through => true ) 
      port map( din => binary_3703_wire, dout => type_cast_3704_wire, req => type_cast_3704_inst_req_0, ack => type_cast_3704_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3653_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(63 downto 0); --
    begin -- 
      ptr_deref_3653_gather_scatter_ack_0 <= ptr_deref_3653_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3653_data_7 & ptr_deref_3653_data_6 & ptr_deref_3653_data_5 & ptr_deref_3653_data_4 & ptr_deref_3653_data_3 & ptr_deref_3653_data_2 & ptr_deref_3653_data_1 & ptr_deref_3653_data_0;
      ptr_deref_3653_wire <= aggregated_sig(63 downto 0);
      --
    end Block;
    ptr_deref_3653_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(15 downto 0); --
    begin -- 
      ptr_deref_3653_root_address_inst_ack_0 <= ptr_deref_3653_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3653_resized_base_address;
      ptr_deref_3653_root_address <= aggregated_sig(15 downto 0);
      --
    end Block;
    if_stmt_3570_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3573_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3570_branch_req_0,
          ack0 => if_stmt_3570_branch_ack_0,
          ack1 => if_stmt_3570_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3614_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3617_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3614_branch_req_0,
          ack0 => if_stmt_3614_branch_ack_0,
          ack1 => if_stmt_3614_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3720_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= binary_3723_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3720_branch_req_0,
          ack0 => if_stmt_3720_branch_ack_0,
          ack1 => if_stmt_3720_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : array_obj_ref_3603_index_0_scale array_obj_ref_3622_index_0_scale 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3602_resized & simple_obj_ref_3621_resized;
      simple_obj_ref_3602_scaled <= data_out(31 downto 16);
      simple_obj_ref_3621_scaled <= data_out(15 downto 0);
      reqL(1) <= array_obj_ref_3603_index_0_scale_req_0;
      reqL(0) <= array_obj_ref_3622_index_0_scale_req_0;
      array_obj_ref_3603_index_0_scale_ack_0 <= ackL(1);
      array_obj_ref_3622_index_0_scale_ack_0 <= ackL(0);
      reqR(1) <= array_obj_ref_3603_index_0_scale_req_1;
      reqR(0) <= array_obj_ref_3622_index_0_scale_req_1;
      array_obj_ref_3603_index_0_scale_ack_1 <= ackR(1);
      array_obj_ref_3622_index_0_scale_ack_1 <= ackR(0);
      SplitOperator: SplitOperatorShared -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000001000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          no_arbitration => false,
          min_clock_period => true,
          num_reqs => 2--
        ) -- 
      port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset);
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : array_obj_ref_3603_root_address_inst 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3603_final_offset & array_obj_ref_3603_resized_base_address;
      array_obj_ref_3603_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3603_root_address_inst_req_0,
          ackL => array_obj_ref_3603_root_address_inst_ack_0,
          reqR => array_obj_ref_3603_root_address_inst_req_1,
          ackR => array_obj_ref_3603_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : array_obj_ref_3622_root_address_inst 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= array_obj_ref_3622_final_offset & array_obj_ref_3622_resized_base_address;
      array_obj_ref_3622_root_address <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => array_obj_ref_3622_root_address_inst_req_0,
          ackL => array_obj_ref_3622_root_address_inst_ack_0,
          reqR => array_obj_ref_3622_root_address_inst_req_1,
          ackR => array_obj_ref_3622_root_address_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : binary_3573_inst 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= wlen_3559;
      binary_3573_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUgt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3573_inst_req_0,
          ackL => binary_3573_inst_ack_0,
          reqR => binary_3573_inst_req_1,
          ackR => binary_3573_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared split operator group (4) : binary_3587_inst 
    SplitOperatorGroup4: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= wlen_3559;
      LI_3588 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3587_inst_req_0,
          ackL => binary_3587_inst_ack_0,
          reqR => binary_3587_inst_req_1,
          ackR => binary_3587_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : binary_3611_inst 
    SplitOperatorGroup5: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= I_3591;
      NI_3612 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3611_inst_req_0,
          ackL => binary_3611_inst_ack_0,
          reqR => binary_3611_inst_req_1,
          ackR => binary_3611_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : binary_3617_inst 
    SplitOperatorGroup6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= NI_3612 & LI_3588;
      binary_3617_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntUlt",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3617_inst_req_0,
          ackL => binary_3617_inst_ack_0,
          reqR => binary_3617_inst_req_1,
          ackR => binary_3617_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : binary_3631_inst 
    SplitOperatorGroup7: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= blen_3562;
      binary_3631_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3631_inst_req_0,
          ackL => binary_3631_inst_ack_0,
          reqR => binary_3631_inst_req_1,
          ackR => binary_3631_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- shared split operator group (8) : binary_3632_inst 
    SplitOperatorGroup8: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= expr_3628_wire_constant & binary_3631_wire;
      binary_3632_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3632_inst_req_0,
          ackL => binary_3632_inst_ack_0,
          reqR => binary_3632_inst_req_1,
          ackR => binary_3632_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- shared split operator group (9) : binary_3634_inst 
    SplitOperatorGroup9: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3632_wire;
      binary_3634_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3634_inst_req_0,
          ackL => binary_3634_inst_ack_0,
          reqR => binary_3634_inst_req_1,
          ackR => binary_3634_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    -- shared split operator group (10) : binary_3636_inst 
    SplitOperatorGroup10: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(7 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3627_wire_constant & type_cast_3635_wire;
      binary_3636_wire <= data_out(7 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntSHL",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 8,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3636_inst_req_0,
          ackL => binary_3636_inst_ack_0,
          reqR => binary_3636_inst_req_1,
          ackR => binary_3636_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- shared split operator group (11) : binary_3675_inst 
    SplitOperatorGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3675_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000001000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3675_inst_req_0,
          ackL => binary_3675_inst_ack_0,
          reqR => binary_3675_inst_req_1,
          ackR => binary_3675_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- shared split operator group (12) : binary_3677_inst 
    SplitOperatorGroup12: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3672_wire & type_cast_3676_wire;
      binary_3677_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3677_inst_req_0,
          ackL => binary_3677_inst_ack_0,
          reqR => binary_3677_inst_req_1,
          ackR => binary_3677_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 12
    -- shared split operator group (13) : binary_3680_inst 
    SplitOperatorGroup13: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3680_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000010000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3680_inst_req_0,
          ackL => binary_3680_inst_ack_0,
          reqR => binary_3680_inst_req_1,
          ackR => binary_3680_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 13
    -- shared split operator group (14) : binary_3684_inst 
    SplitOperatorGroup14: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3684_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000011000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3684_inst_req_0,
          ackL => binary_3684_inst_ack_0,
          reqR => binary_3684_inst_req_1,
          ackR => binary_3684_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 14
    -- shared split operator group (15) : binary_3686_inst 
    SplitOperatorGroup15: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3681_wire & type_cast_3685_wire;
      binary_3686_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3686_inst_req_0,
          ackL => binary_3686_inst_ack_0,
          reqR => binary_3686_inst_req_1,
          ackR => binary_3686_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 15
    -- shared split operator group (16) : binary_3687_inst 
    SplitOperatorGroup16: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3677_wire & binary_3686_wire;
      binary_3687_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3687_inst_req_0,
          ackL => binary_3687_inst_ack_0,
          reqR => binary_3687_inst_req_1,
          ackR => binary_3687_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 16
    -- shared split operator group (17) : binary_3690_inst 
    SplitOperatorGroup17: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3690_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000100000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3690_inst_req_0,
          ackL => binary_3690_inst_ack_0,
          reqR => binary_3690_inst_req_1,
          ackR => binary_3690_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 17
    -- shared split operator group (18) : binary_3694_inst 
    SplitOperatorGroup18: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3694_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000101000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3694_inst_req_0,
          ackL => binary_3694_inst_ack_0,
          reqR => binary_3694_inst_req_1,
          ackR => binary_3694_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 18
    -- shared split operator group (19) : binary_3696_inst 
    SplitOperatorGroup19: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3691_wire & type_cast_3695_wire;
      binary_3696_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3696_inst_req_0,
          ackL => binary_3696_inst_ack_0,
          reqR => binary_3696_inst_req_1,
          ackR => binary_3696_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 19
    -- shared split operator group (20) : binary_3699_inst 
    SplitOperatorGroup20: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3699_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000110000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3699_inst_req_0,
          ackL => binary_3699_inst_ack_0,
          reqR => binary_3699_inst_req_1,
          ackR => binary_3699_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 20
    -- shared split operator group (21) : binary_3703_inst 
    SplitOperatorGroup21: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= a_3668;
      binary_3703_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntLSHR",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 64,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0000000000000000000000000000000000000000000000000000000000111000",
          constant_width => 64,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3703_inst_req_0,
          ackL => binary_3703_inst_ack_0,
          reqR => binary_3703_inst_req_1,
          ackR => binary_3703_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 21
    -- shared split operator group (22) : binary_3705_inst 
    SplitOperatorGroup22: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= type_cast_3700_wire & type_cast_3704_wire;
      binary_3705_wire <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 8,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3705_inst_req_0,
          ackL => binary_3705_inst_ack_0,
          reqR => binary_3705_inst_req_1,
          ackR => binary_3705_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 22
    -- shared split operator group (23) : binary_3706_inst 
    SplitOperatorGroup23: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3696_wire & binary_3705_wire;
      binary_3706_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3706_inst_req_0,
          ackL => binary_3706_inst_ack_0,
          reqR => binary_3706_inst_req_1,
          ackR => binary_3706_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 23
    -- shared split operator group (24) : binary_3707_inst 
    SplitOperatorGroup24: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= binary_3687_wire & binary_3706_wire;
      binary_3707_wire <= data_out(63 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApConcat",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 64,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3707_inst_req_0,
          ackL => binary_3707_inst_ack_0,
          reqR => binary_3707_inst_req_1,
          ackR => binary_3707_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 24
    -- shared split operator group (25) : binary_3723_inst 
    SplitOperatorGroup25: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3721_wire;
      binary_3723_wire <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNe",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => binary_3723_inst_req_0,
          ackL => binary_3723_inst_ack_0,
          reqR => binary_3723_inst_req_1,
          ackR => binary_3723_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 25
    -- shared split operator group (26) : binary_3728_inst 
    SplitOperatorGroup26: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= simple_obj_ref_3726_wire;
      binary_3728_wire <= data_out(31 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "11111111111111111111100000000000",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => true--
        ) 
        port map ( -- 
          reqL => binary_3728_inst_req_0,
          ackL => binary_3728_inst_ack_0,
          reqR => binary_3728_inst_req_1,
          ackR => binary_3728_inst_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 26
    -- shared split operator group (27) : ptr_deref_3653_addr_0 
    SplitOperatorGroup27: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_0 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000000",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_0_req_0,
          ackL => ptr_deref_3653_addr_0_ack_0,
          reqR => ptr_deref_3653_addr_0_req_1,
          ackR => ptr_deref_3653_addr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 27
    -- shared split operator group (28) : ptr_deref_3653_addr_1 
    SplitOperatorGroup28: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_1 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000001",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_1_req_0,
          ackL => ptr_deref_3653_addr_1_ack_0,
          reqR => ptr_deref_3653_addr_1_req_1,
          ackR => ptr_deref_3653_addr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 28
    -- shared split operator group (29) : ptr_deref_3653_addr_2 
    SplitOperatorGroup29: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_2 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000010",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_2_req_0,
          ackL => ptr_deref_3653_addr_2_ack_0,
          reqR => ptr_deref_3653_addr_2_req_1,
          ackR => ptr_deref_3653_addr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 29
    -- shared split operator group (30) : ptr_deref_3653_addr_3 
    SplitOperatorGroup30: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_3 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000011",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_3_req_0,
          ackL => ptr_deref_3653_addr_3_ack_0,
          reqR => ptr_deref_3653_addr_3_req_1,
          ackR => ptr_deref_3653_addr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 30
    -- shared split operator group (31) : ptr_deref_3653_addr_4 
    SplitOperatorGroup31: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_4 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000100",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_4_req_0,
          ackL => ptr_deref_3653_addr_4_ack_0,
          reqR => ptr_deref_3653_addr_4_req_1,
          ackR => ptr_deref_3653_addr_4_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 31
    -- shared split operator group (32) : ptr_deref_3653_addr_5 
    SplitOperatorGroup32: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_5 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000101",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_5_req_0,
          ackL => ptr_deref_3653_addr_5_ack_0,
          reqR => ptr_deref_3653_addr_5_req_1,
          ackR => ptr_deref_3653_addr_5_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 32
    -- shared split operator group (33) : ptr_deref_3653_addr_6 
    SplitOperatorGroup33: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_6 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000110",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_6_req_0,
          ackL => ptr_deref_3653_addr_6_ack_0,
          reqR => ptr_deref_3653_addr_6_req_1,
          ackR => ptr_deref_3653_addr_6_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 33
    -- shared split operator group (34) : ptr_deref_3653_addr_7 
    SplitOperatorGroup34: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(15 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= ptr_deref_3653_root_address;
      ptr_deref_3653_word_address_7 <= data_out(15 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 16,
          constant_operand => "0000000000000111",
          constant_width => 16,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => ptr_deref_3653_addr_7_req_0,
          ackL => ptr_deref_3653_addr_7_ack_0,
          reqR => ptr_deref_3653_addr_7_req_1,
          ackR => ptr_deref_3653_addr_7_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 34
    -- shared load operator group (0) : ptr_deref_3653_load_0 ptr_deref_3653_load_6 ptr_deref_3653_load_2 ptr_deref_3653_load_4 ptr_deref_3653_load_5 ptr_deref_3653_load_1 ptr_deref_3653_load_3 ptr_deref_3653_load_7 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3653_load_0_req_0,
        ptr_deref_3653_load_0_ack_0,
        ptr_deref_3653_load_0_req_1,
        ptr_deref_3653_load_0_ack_1,
        "ptr_deref_3653_load_0",
        "memory_space_5" ,
        ptr_deref_3653_data_0,
        ptr_deref_3653_word_address_0,
        "ptr_deref_3653_data_0",
        "ptr_deref_3653_word_address_0" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_6_req_0,
        ptr_deref_3653_load_6_ack_0,
        ptr_deref_3653_load_6_req_1,
        ptr_deref_3653_load_6_ack_1,
        "ptr_deref_3653_load_6",
        "memory_space_5" ,
        ptr_deref_3653_data_6,
        ptr_deref_3653_word_address_6,
        "ptr_deref_3653_data_6",
        "ptr_deref_3653_word_address_6" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_2_req_0,
        ptr_deref_3653_load_2_ack_0,
        ptr_deref_3653_load_2_req_1,
        ptr_deref_3653_load_2_ack_1,
        "ptr_deref_3653_load_2",
        "memory_space_5" ,
        ptr_deref_3653_data_2,
        ptr_deref_3653_word_address_2,
        "ptr_deref_3653_data_2",
        "ptr_deref_3653_word_address_2" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_4_req_0,
        ptr_deref_3653_load_4_ack_0,
        ptr_deref_3653_load_4_req_1,
        ptr_deref_3653_load_4_ack_1,
        "ptr_deref_3653_load_4",
        "memory_space_5" ,
        ptr_deref_3653_data_4,
        ptr_deref_3653_word_address_4,
        "ptr_deref_3653_data_4",
        "ptr_deref_3653_word_address_4" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_5_req_0,
        ptr_deref_3653_load_5_ack_0,
        ptr_deref_3653_load_5_req_1,
        ptr_deref_3653_load_5_ack_1,
        "ptr_deref_3653_load_5",
        "memory_space_5" ,
        ptr_deref_3653_data_5,
        ptr_deref_3653_word_address_5,
        "ptr_deref_3653_data_5",
        "ptr_deref_3653_word_address_5" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_1_req_0,
        ptr_deref_3653_load_1_ack_0,
        ptr_deref_3653_load_1_req_1,
        ptr_deref_3653_load_1_ack_1,
        "ptr_deref_3653_load_1",
        "memory_space_5" ,
        ptr_deref_3653_data_1,
        ptr_deref_3653_word_address_1,
        "ptr_deref_3653_data_1",
        "ptr_deref_3653_word_address_1" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_3_req_0,
        ptr_deref_3653_load_3_ack_0,
        ptr_deref_3653_load_3_req_1,
        ptr_deref_3653_load_3_ack_1,
        "ptr_deref_3653_load_3",
        "memory_space_5" ,
        ptr_deref_3653_data_3,
        ptr_deref_3653_word_address_3,
        "ptr_deref_3653_data_3",
        "ptr_deref_3653_word_address_3" -- 
      );
      LogMemRead(clk, -- 
        ptr_deref_3653_load_7_req_0,
        ptr_deref_3653_load_7_ack_0,
        ptr_deref_3653_load_7_req_1,
        ptr_deref_3653_load_7_ack_1,
        "ptr_deref_3653_load_7",
        "memory_space_5" ,
        ptr_deref_3653_data_7,
        ptr_deref_3653_word_address_7,
        "ptr_deref_3653_data_7",
        "ptr_deref_3653_word_address_7" -- 
      );
      reqL(7) <= ptr_deref_3653_load_0_req_0;
      reqL(6) <= ptr_deref_3653_load_6_req_0;
      reqL(5) <= ptr_deref_3653_load_2_req_0;
      reqL(4) <= ptr_deref_3653_load_4_req_0;
      reqL(3) <= ptr_deref_3653_load_5_req_0;
      reqL(2) <= ptr_deref_3653_load_1_req_0;
      reqL(1) <= ptr_deref_3653_load_3_req_0;
      reqL(0) <= ptr_deref_3653_load_7_req_0;
      ptr_deref_3653_load_0_ack_0 <= ackL(7);
      ptr_deref_3653_load_6_ack_0 <= ackL(6);
      ptr_deref_3653_load_2_ack_0 <= ackL(5);
      ptr_deref_3653_load_4_ack_0 <= ackL(4);
      ptr_deref_3653_load_5_ack_0 <= ackL(3);
      ptr_deref_3653_load_1_ack_0 <= ackL(2);
      ptr_deref_3653_load_3_ack_0 <= ackL(1);
      ptr_deref_3653_load_7_ack_0 <= ackL(0);
      reqR(7) <= ptr_deref_3653_load_0_req_1;
      reqR(6) <= ptr_deref_3653_load_6_req_1;
      reqR(5) <= ptr_deref_3653_load_2_req_1;
      reqR(4) <= ptr_deref_3653_load_4_req_1;
      reqR(3) <= ptr_deref_3653_load_5_req_1;
      reqR(2) <= ptr_deref_3653_load_1_req_1;
      reqR(1) <= ptr_deref_3653_load_3_req_1;
      reqR(0) <= ptr_deref_3653_load_7_req_1;
      ptr_deref_3653_load_0_ack_1 <= ackR(7);
      ptr_deref_3653_load_6_ack_1 <= ackR(6);
      ptr_deref_3653_load_2_ack_1 <= ackR(5);
      ptr_deref_3653_load_4_ack_1 <= ackR(4);
      ptr_deref_3653_load_5_ack_1 <= ackR(3);
      ptr_deref_3653_load_1_ack_1 <= ackR(2);
      ptr_deref_3653_load_3_ack_1 <= ackR(1);
      ptr_deref_3653_load_7_ack_1 <= ackR(0);
      data_in <= ptr_deref_3653_word_address_0 & ptr_deref_3653_word_address_6 & ptr_deref_3653_word_address_2 & ptr_deref_3653_word_address_4 & ptr_deref_3653_word_address_5 & ptr_deref_3653_word_address_1 & ptr_deref_3653_word_address_3 & ptr_deref_3653_word_address_7;
      ptr_deref_3653_data_0 <= data_out(63 downto 56);
      ptr_deref_3653_data_6 <= data_out(55 downto 48);
      ptr_deref_3653_data_2 <= data_out(47 downto 40);
      ptr_deref_3653_data_4 <= data_out(39 downto 32);
      ptr_deref_3653_data_5 <= data_out(31 downto 24);
      ptr_deref_3653_data_1 <= data_out(23 downto 16);
      ptr_deref_3653_data_3 <= data_out(15 downto 8);
      ptr_deref_3653_data_7 <= data_out(7 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 16,
        num_reqs => 8,
        tag_length => 5,
        time_stamp_width => 6,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_5_lr_req(0),
          mack => memory_space_5_lr_ack(0),
          maddr => memory_space_5_lr_addr(15 downto 0),
          mtag => memory_space_5_lr_tag(10 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 8,  num_reqs => 8,  tag_length => 5,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_5_lc_req(0),
          mack => memory_space_5_lc_ack(0),
          mdata => memory_space_5_lc_data(7 downto 0),
          mtag => memory_space_5_lc_tag(4 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    xxsend_packet_pipelinexxblen_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxblen_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxblen_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxblen_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxblen_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxblen_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxblen_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxbuf64_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxfree_packet_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxfree_packet_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxfree_packet_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxfree_packet_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxfree_packet_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxfree_packet_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxfree_packet_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxpkt64_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_ctrl_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_last_word_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_last_word_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_last_word_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_last_word_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_last_word_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxread_pointer_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 32,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxread_pointer_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxread_pointer_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxread_pointer_pipe_read_data,
        write_req => xxsend_packet_pipelinexxread_pointer_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxread_pointer_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxread_pointer_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_ctrl_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 8,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_data_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 64,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_data_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_data_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_data_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_data_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_data_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_data_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxswap_last_word_in_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 1,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data,
        write_req => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    xxsend_packet_pipelinexxwlen_pipe_Pipe: PipeBase -- 
      generic map( -- 
        num_reads => 1,
        num_writes => 1,
        data_width => 16,
        depth => 2 --
      )
      port map( -- 
        read_req => xxsend_packet_pipelinexxwlen_pipe_pipe_read_req,
        read_ack => xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack,
        read_data => xxsend_packet_pipelinexxwlen_pipe_pipe_read_data,
        write_req => xxsend_packet_pipelinexxwlen_pipe_pipe_write_req,
        write_ack => xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack,
        write_data => xxsend_packet_pipelinexxwlen_pipe_pipe_write_data,
        clk => clk,reset => reset -- 
      ); -- 
    -- shared inport operator group (0) : simple_obj_ref_3524_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3524_inst_ack_0 then -- 
            assert false report " ReadPipe send_packet_pipe to wire pkt_3525 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3524_inst_req_0;
      simple_obj_ref_3524_inst_ack_0 <= ack(0);
      pkt_3525 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => send_packet_pipe_pipe_read_req(0),
          oack => send_packet_pipe_pipe_read_ack(0),
          odata => send_packet_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_3558_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3558_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxwlen_pipe to wire wlen_3559 value="  &  convert_slv_to_hex_string(data_out(15 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3558_inst_req_0;
      simple_obj_ref_3558_inst_ack_0 <= ack(0);
      wlen_3559 <= data_out(15 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxwlen_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxwlen_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxwlen_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_3561_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3561_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxblen_pipe to wire blen_3562 value="  &  convert_slv_to_hex_string(data_out(15 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3561_inst_req_0;
      simple_obj_ref_3561_inst_ack_0 <= ack(0);
      blen_3562 <= data_out(15 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxblen_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxblen_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxblen_pipe_pipe_read_data(15 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_3564_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3564_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxbuf64_pipe to wire buf64_3565 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3564_inst_req_0;
      simple_obj_ref_3564_inst_ack_0 <= ack(0);
      buf64_3565 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxbuf64_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_3567_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3567_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxpkt64_pipe to wire pkt64_3568 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3567_inst_req_0;
      simple_obj_ref_3567_inst_ack_0 <= ack(0);
      pkt64_3568 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxpkt64_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- shared inport operator group (5) : simple_obj_ref_3652_inst 
    InportGroup5: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3652_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_pointer to wire simple_obj_ref_3652_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3652_inst_req_0;
      simple_obj_ref_3652_inst_ack_0 <= ack(0);
      simple_obj_ref_3652_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_pointer_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_pointer_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_pointer_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 5
    -- shared inport operator group (6) : simple_obj_ref_3656_inst 
    InportGroup6: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3656_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_ctrl_in to wire simple_obj_ref_3656_wire value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3656_inst_req_0;
      simple_obj_ref_3656_inst_ack_0 <= ack(0);
      simple_obj_ref_3656_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_ctrl_in_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 6
    -- shared inport operator group (7) : simple_obj_ref_3659_inst 
    InportGroup7: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3659_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxread_last_word_in to wire simple_obj_ref_3659_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3659_inst_req_0;
      simple_obj_ref_3659_inst_ack_0 <= ack(0);
      simple_obj_ref_3659_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxread_last_word_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxread_last_word_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxread_last_word_in_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 7
    -- shared inport operator group (8) : simple_obj_ref_3667_inst 
    InportGroup8: Block -- 
      signal data_out: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3667_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_data_in to wire a_3668 value="  &  convert_slv_to_hex_string(data_out(63 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3667_inst_req_0;
      simple_obj_ref_3667_inst_ack_0 <= ack(0);
      a_3668 <= data_out(63 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_data_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_data_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_data_in_pipe_read_data(63 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 8
    -- shared inport operator group (9) : simple_obj_ref_3710_inst 
    InportGroup9: Block -- 
      signal data_out: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3710_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_ctrl_in to wire simple_obj_ref_3710_wire value="  &  convert_slv_to_hex_string(data_out(7 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3710_inst_req_0;
      simple_obj_ref_3710_inst_ack_0 <= ack(0);
      simple_obj_ref_3710_wire <= data_out(7 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_ctrl_in_pipe_read_data(7 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 9
    -- shared inport operator group (10) : simple_obj_ref_3713_inst 
    InportGroup10: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3713_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxswap_last_word_in to wire simple_obj_ref_3713_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3713_inst_req_0;
      simple_obj_ref_3713_inst_ack_0 <= ack(0);
      simple_obj_ref_3713_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxswap_last_word_in_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 10
    -- shared inport operator group (11) : simple_obj_ref_3721_inst 
    InportGroup11: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3721_inst_ack_0 then -- 
            assert false report " ReadPipe xxsend_packet_pipelinexxfree_packet_in to wire simple_obj_ref_3721_wire value="  &  convert_slv_to_hex_string(data_out(0 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3721_inst_req_0;
      simple_obj_ref_3721_inst_ack_0 <= ack(0);
      simple_obj_ref_3721_wire <= data_out(0 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => xxsend_packet_pipelinexxfree_packet_in_pipe_read_req(0),
          oack => xxsend_packet_pipelinexxfree_packet_in_pipe_read_ack(0),
          odata => xxsend_packet_pipelinexxfree_packet_in_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 11
    -- shared inport operator group (12) : simple_obj_ref_3726_inst 
    InportGroup12: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3726_inst_ack_0 then -- 
            assert false report " ReadPipe send_packet_buf_queue to wire simple_obj_ref_3726_wire value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3726_inst_req_0;
      simple_obj_ref_3726_inst_ack_0 <= ack(0);
      simple_obj_ref_3726_wire <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => send_packet_buf_queue_pipe_read_req(0),
          oack => send_packet_buf_queue_pipe_read_ack(0),
          odata => send_packet_buf_queue_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 12
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3533_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxbuf64_pipe from wire type_cast_3535_wire value="  &  convert_slv_to_hex_string(type_cast_3535_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3533_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3533_inst_req_0;
      simple_obj_ref_3533_inst_ack_0 <= ack(0);
      data_in <= type_cast_3535_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxbuf64_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3537_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxpkt64_pipe from wire type_cast_3539_wire value="  &  convert_slv_to_hex_string(type_cast_3539_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (1) : simple_obj_ref_3537_inst 
    OutportGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3537_inst_req_0;
      simple_obj_ref_3537_inst_ack_0 <= ack(0);
      data_in <= type_cast_3539_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxpkt64_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3541_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxwlen_pipe from wire wlen_3531 value="  &  convert_slv_to_hex_string(wlen_3531) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (2) : simple_obj_ref_3541_inst 
    OutportGroup2: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3541_inst_req_0;
      simple_obj_ref_3541_inst_ack_0 <= ack(0);
      data_in <= wlen_3531;
      outport: OutputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxwlen_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxwlen_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxwlen_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3544_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxblen_pipe from wire blen_3531 value="  &  convert_slv_to_hex_string(blen_3531) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (3) : simple_obj_ref_3544_inst 
    OutportGroup3: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3544_inst_req_0;
      simple_obj_ref_3544_inst_ack_0 <= ack(0);
      data_in <= blen_3531;
      outport: OutputPort -- 
        generic map ( data_width => 16,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxblen_pipe_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxblen_pipe_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxblen_pipe_pipe_write_data(15 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3547_inst_ack_0 then -- 
          assert false report " WritePipe send_packet_buf_queue from wire type_cast_3549_wire value="  &  convert_slv_to_hex_string(type_cast_3549_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (4) : simple_obj_ref_3547_inst 
    OutportGroup4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3547_inst_req_0;
      simple_obj_ref_3547_inst_ack_0 <= ack(0);
      data_in <= type_cast_3549_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => send_packet_buf_queue_pipe_write_req(0),
          oack => send_packet_buf_queue_pipe_write_ack(0),
          odata => send_packet_buf_queue_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3625_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire binary_3636_wire value="  &  convert_slv_to_hex_string(binary_3636_wire) severity note; --
        end if;
        if simple_obj_ref_3598_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire expr_3599_wire_constant value="  &  convert_slv_to_hex_string(expr_3599_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3575_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_ctrl_in from wire expr_3576_wire_constant value="  &  convert_slv_to_hex_string(expr_3576_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (5) : simple_obj_ref_3625_inst simple_obj_ref_3598_inst simple_obj_ref_3575_inst 
    OutportGroup5: Block -- 
      signal data_in: std_logic_vector(23 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_3625_inst_req_0;
      req(1) <= simple_obj_ref_3598_inst_req_0;
      req(0) <= simple_obj_ref_3575_inst_req_0;
      simple_obj_ref_3625_inst_ack_0 <= ack(2);
      simple_obj_ref_3598_inst_ack_0 <= ack(1);
      simple_obj_ref_3575_inst_ack_0 <= ack(0);
      data_in <= binary_3636_wire & expr_3599_wire_constant & expr_3576_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_ctrl_in_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 5
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3638_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire last_word_ptr_3623 value="  &  convert_slv_to_hex_string(last_word_ptr_3623) severity note; --
        end if;
        if simple_obj_ref_3601_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire array_obj_ref_3603_wire value="  &  convert_slv_to_hex_string(array_obj_ref_3603_wire) severity note; --
        end if;
        if simple_obj_ref_3578_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_pointer from wire buf64_3565 value="  &  convert_slv_to_hex_string(buf64_3565) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (6) : simple_obj_ref_3638_inst simple_obj_ref_3601_inst simple_obj_ref_3578_inst 
    OutportGroup6: Block -- 
      signal data_in: std_logic_vector(95 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_3638_inst_req_0;
      req(1) <= simple_obj_ref_3601_inst_req_0;
      req(0) <= simple_obj_ref_3578_inst_req_0;
      simple_obj_ref_3638_inst_ack_0 <= ack(2);
      simple_obj_ref_3601_inst_ack_0 <= ack(1);
      simple_obj_ref_3578_inst_ack_0 <= ack(0);
      data_in <= last_word_ptr_3623 & array_obj_ref_3603_wire & buf64_3565;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_pointer_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_pointer_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_pointer_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 6
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3605_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_3606_wire_constant value="  &  convert_slv_to_hex_string(expr_3606_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3581_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_3582_wire_constant value="  &  convert_slv_to_hex_string(expr_3582_wire_constant) severity note; --
        end if;
        if simple_obj_ref_3641_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxread_last_word_in from wire expr_3642_wire_constant value="  &  convert_slv_to_hex_string(expr_3642_wire_constant) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (7) : simple_obj_ref_3605_inst simple_obj_ref_3581_inst simple_obj_ref_3641_inst 
    OutportGroup7: Block -- 
      signal data_in: std_logic_vector(2 downto 0);
      signal req, ack : BooleanArray( 2 downto 0);
      -- 
    begin -- 
      req(2) <= simple_obj_ref_3605_inst_req_0;
      req(1) <= simple_obj_ref_3581_inst_req_0;
      req(0) <= simple_obj_ref_3641_inst_req_0;
      simple_obj_ref_3605_inst_ack_0 <= ack(2);
      simple_obj_ref_3581_inst_ack_0 <= ack(1);
      simple_obj_ref_3641_inst_ack_0 <= ack(0);
      data_in <= expr_3606_wire_constant & expr_3582_wire_constant & expr_3642_wire_constant;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 3,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxread_last_word_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxread_last_word_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxread_last_word_in_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 7
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3651_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_data_in from wire ptr_deref_3653_wire value="  &  convert_slv_to_hex_string(ptr_deref_3653_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (8) : simple_obj_ref_3651_inst 
    OutportGroup8: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3651_inst_req_0;
      simple_obj_ref_3651_inst_ack_0 <= ack(0);
      data_in <= ptr_deref_3653_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_data_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_data_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_data_in_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 8
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3655_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_ctrl_in from wire simple_obj_ref_3656_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3656_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (9) : simple_obj_ref_3655_inst 
    OutportGroup9: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3655_inst_req_0;
      simple_obj_ref_3655_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3656_wire;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_ctrl_in_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 9
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3658_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxswap_last_word_in from wire simple_obj_ref_3659_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3659_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (10) : simple_obj_ref_3658_inst 
    OutportGroup10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3658_inst_req_0;
      simple_obj_ref_3658_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3659_wire;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxswap_last_word_in_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 10
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3670_inst_ack_0 then -- 
          assert false report " WritePipe out_data from wire binary_3707_wire value="  &  convert_slv_to_hex_string(binary_3707_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (11) : simple_obj_ref_3670_inst 
    OutportGroup11: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3670_inst_req_0;
      simple_obj_ref_3670_inst_ack_0 <= ack(0);
      data_in <= binary_3707_wire;
      outport: OutputPort -- 
        generic map ( data_width => 64,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_write_req(0),
          oack => out_data_pipe_write_ack(0),
          odata => out_data_pipe_write_data(63 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 11
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3709_inst_ack_0 then -- 
          assert false report " WritePipe out_ctrl from wire simple_obj_ref_3710_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3710_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (12) : simple_obj_ref_3709_inst 
    OutportGroup12: Block -- 
      signal data_in: std_logic_vector(7 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3709_inst_req_0;
      simple_obj_ref_3709_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3710_wire;
      outport: OutputPort -- 
        generic map ( data_width => 8,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_ctrl_pipe_write_req(0),
          oack => out_ctrl_pipe_write_ack(0),
          odata => out_ctrl_pipe_write_data(7 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 12
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3712_inst_ack_0 then -- 
          assert false report " WritePipe xxsend_packet_pipelinexxfree_packet_in from wire simple_obj_ref_3713_wire value="  &  convert_slv_to_hex_string(simple_obj_ref_3713_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (13) : simple_obj_ref_3712_inst 
    OutportGroup13: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3712_inst_req_0;
      simple_obj_ref_3712_inst_ack_0 <= ack(0);
      data_in <= simple_obj_ref_3713_wire;
      outport: OutputPort -- 
        generic map ( data_width => 1,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => xxsend_packet_pipelinexxfree_packet_in_pipe_write_req(0),
          oack => xxsend_packet_pipelinexxfree_packet_in_pipe_write_ack(0),
          odata => xxsend_packet_pipelinexxfree_packet_in_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 13
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3725_inst_ack_0 then -- 
          assert false report " WritePipe free_queue_pipe from wire binary_3728_wire value="  &  convert_slv_to_hex_string(binary_3728_wire) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (14) : simple_obj_ref_3725_inst 
    OutportGroup14: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3725_inst_req_0;
      simple_obj_ref_3725_inst_ack_0 <= ack(0);
      data_in <= binary_3728_wire;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => free_queue_pipe_pipe_write_req(0),
          oack => free_queue_pipe_pipe_write_ack(0),
          odata => free_queue_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 14
    -- shared call operator group (0) : call_stmt_3531_call 
    CallGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3531_call_req_0;
      call_stmt_3531_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3531_call_req_1;
      call_stmt_3531_call_ack_1 <= ackR(0);
      data_in <= type_cast_3527_wire;
      buf_3531 <= data_out(63 downto 32);
      wlen_3531 <= data_out(31 downto 16);
      blen_3531 <= data_out(15 downto 0);
      CallReq: InputMuxBase -- 
        generic map (  iwidth => 32,
        owidth => 32,
        twidth => 1,
        nreqs => 1,
        registered_output => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => analyze_packet_call_reqs(0),
          ackR => analyze_packet_call_acks(0),
          dataR => analyze_packet_call_data(31 downto 0),
          tagR => analyze_packet_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBase -- 
        generic map ( 
        iwidth => 64, owidth => 64, twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => analyze_packet_return_acks(0), -- cross-over
          ackL => analyze_packet_return_reqs(0), -- cross-over
          dataL => analyze_packet_return_data(63 downto 0),
          tagL => analyze_packet_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_input is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    receive_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    receive_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    src_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
    src_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
    src_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
    global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
    global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
    free_queue_init_call_reqs : out  std_logic_vector(0 downto 0);
    free_queue_init_call_acks : in   std_logic_vector(0 downto 0);
    free_queue_init_call_tag  :  out  std_logic_vector(0 downto 0);
    free_queue_init_return_reqs : out  std_logic_vector(0 downto 0);
    free_queue_init_return_acks : in   std_logic_vector(0 downto 0);
    free_queue_init_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_input;
architecture Default of wrapper_input is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_input_CP_19182_start: Boolean;
  -- links between control-path and data-path
  signal ptr_deref_3751_base_resize_req_0 : boolean;
  signal ptr_deref_3756_base_resize_ack_0 : boolean;
  signal ptr_deref_3751_addr_0_ack_0 : boolean;
  signal ptr_deref_3751_base_resize_ack_0 : boolean;
  signal simple_obj_ref_3748_inst_req_0 : boolean;
  signal ptr_deref_3756_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3756_root_address_inst_req_0 : boolean;
  signal ptr_deref_3756_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3756_base_resize_req_0 : boolean;
  signal call_stmt_3744_call_req_0 : boolean;
  signal ptr_deref_3751_root_address_inst_ack_0 : boolean;
  signal call_stmt_3744_call_req_1 : boolean;
  signal ptr_deref_3756_addr_0_req_0 : boolean;
  signal ptr_deref_3751_store_0_ack_0 : boolean;
  signal call_stmt_3744_call_ack_0 : boolean;
  signal ptr_deref_3756_addr_0_ack_0 : boolean;
  signal call_stmt_3744_call_ack_1 : boolean;
  signal ptr_deref_3751_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3751_store_0_req_0 : boolean;
  signal simple_obj_ref_3758_inst_req_0 : boolean;
  signal simple_obj_ref_3758_inst_ack_0 : boolean;
  signal ptr_deref_3751_store_0_ack_1 : boolean;
  signal ptr_deref_3751_store_0_req_1 : boolean;
  signal ptr_deref_3751_addr_0_req_0 : boolean;
  signal ptr_deref_3751_gather_scatter_req_0 : boolean;
  signal ptr_deref_3751_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_3748_inst_ack_0 : boolean;
  signal ptr_deref_3756_load_0_req_0 : boolean;
  signal ptr_deref_3756_load_0_ack_0 : boolean;
  signal call_stmt_3743_call_req_0 : boolean;
  signal call_stmt_3743_call_ack_0 : boolean;
  signal ptr_deref_3756_load_0_req_1 : boolean;
  signal ptr_deref_3756_load_0_ack_1 : boolean;
  signal call_stmt_3743_call_req_1 : boolean;
  signal call_stmt_3743_call_ack_1 : boolean;
  signal ptr_deref_3756_gather_scatter_req_0 : boolean;
  signal memory_space_7_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_7_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_7_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_7_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_7_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_7_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_7_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_7_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_input_CP_19182: Block -- control-path 
    signal cp_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(2);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(2), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    crr_19218_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => call_stmt_3743_call_req_0); -- 
    cp_elements(1) <= cp_elements(29);
    pipe_wreq_19365_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => simple_obj_ref_3758_inst_req_0); -- 
    cp_elements(2) <= false; 
    cra_19219_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3743_call_ack_0, ack => cp_elements(3)); -- 
    ccr_19223_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => call_stmt_3743_call_req_1); -- 
    cca_19224_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3743_call_ack_1, ack => cp_elements(4)); -- 
    crr_19235_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(4), ack => call_stmt_3744_call_req_0); -- 
    cra_19236_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3744_call_ack_0, ack => cp_elements(5)); -- 
    ccr_19240_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(5), ack => call_stmt_3744_call_req_1); -- 
    cca_19241_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3744_call_ack_1, ack => cp_elements(6)); -- 
    ack_19254_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3748_inst_ack_0, ack => cp_elements(7)); -- 
    cp_elements(8) <= cp_elements(7);
    cp_elements(9) <= cp_elements(8);
    cpelement_group_10 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(9) & cp_elements(11) & cp_elements(15));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(10),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19286_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_3751_gather_scatter_req_0); -- 
    cp_elements(11) <= cp_elements(8);
    cp_elements(12) <= cp_elements(11);
    base_resize_req_19271_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => ptr_deref_3751_base_resize_req_0); -- 
    base_resize_ack_19272_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3751_base_resize_ack_0, ack => cp_elements(13)); -- 
    sum_rename_req_19276_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_3751_root_address_inst_req_0); -- 
    sum_rename_ack_19277_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3751_root_address_inst_ack_0, ack => cp_elements(14)); -- 
    root_rename_req_19281_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(14), ack => ptr_deref_3751_addr_0_req_0); -- 
    root_rename_ack_19282_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3751_addr_0_ack_0, ack => cp_elements(15)); -- 
    split_ack_19287_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3751_gather_scatter_ack_0, ack => cp_elements(16)); -- 
    rr_19294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => ptr_deref_3751_store_0_req_0); -- 
    cp_elements(17) <= ptr_deref_3751_store_0_ack_0;
    cp_elements(18) <= cp_elements(17);
    cr_19305_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => ptr_deref_3751_store_0_req_1); -- 
    ca_19306_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3751_store_0_ack_1, ack => cp_elements(19)); -- 
    cpelement_group_20 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(17) & cp_elements(21) & cp_elements(25));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(20),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19340_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_3756_load_0_req_0); -- 
    cp_elements(21) <= cp_elements(8);
    cp_elements(22) <= cp_elements(21);
    base_resize_req_19319_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(22), ack => ptr_deref_3756_base_resize_req_0); -- 
    base_resize_ack_19320_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_base_resize_ack_0, ack => cp_elements(23)); -- 
    sum_rename_req_19324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => ptr_deref_3756_root_address_inst_req_0); -- 
    sum_rename_ack_19325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_root_address_inst_ack_0, ack => cp_elements(24)); -- 
    root_rename_req_19329_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => ptr_deref_3756_addr_0_req_0); -- 
    root_rename_ack_19330_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_addr_0_ack_0, ack => cp_elements(25)); -- 
    ra_19341_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_load_0_ack_0, ack => cp_elements(26)); -- 
    cr_19351_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => ptr_deref_3756_load_0_req_1); -- 
    ca_19352_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_load_0_ack_1, ack => cp_elements(27)); -- 
    merge_req_19353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => ptr_deref_3756_gather_scatter_req_0); -- 
    merge_ack_19354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3756_gather_scatter_ack_0, ack => cp_elements(28)); -- 
    cpelement_group_29 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(19) & cp_elements(28));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(29),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    pipe_wack_19366_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3758_inst_ack_0, ack => cp_elements(30)); -- 
    cp_elements(31) <= OrReduce(cp_elements(6) & cp_elements(30));
    cp_elements(32) <= cp_elements(31);
    req_19253_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => simple_obj_ref_3748_inst_req_0); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal buf1_3742 : std_logic_vector(31 downto 0);
    signal iNsTr_4_3749 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3757 : std_logic_vector(31 downto 0);
    signal ptr_deref_3751_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3751_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3751_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3751_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3751_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3751_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3756_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3756_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3756_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3756_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3756_word_offset_0 : std_logic_vector(0 downto 0);
    signal xxwrapper_inputxxbodyxxbuf1_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    buf1_3742 <= "00000000000000000000000000000000";
    ptr_deref_3751_word_offset_0 <= "0";
    ptr_deref_3756_word_offset_0 <= "0";
    xxwrapper_inputxxbodyxxbuf1_alloc_base_address <= "0";
    ptr_deref_3751_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => buf1_3742, dout => ptr_deref_3751_resized_base_address, req => ptr_deref_3751_base_resize_req_0, ack => ptr_deref_3751_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3756_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => buf1_3742, dout => ptr_deref_3756_resized_base_address, req => ptr_deref_3756_base_resize_req_0, ack => ptr_deref_3756_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3751_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3751_addr_0_ack_0 <= ptr_deref_3751_addr_0_req_0;
      aggregated_sig <= ptr_deref_3751_root_address;
      ptr_deref_3751_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3751_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3751_gather_scatter_ack_0 <= ptr_deref_3751_gather_scatter_req_0;
      aggregated_sig <= iNsTr_4_3749;
      ptr_deref_3751_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3751_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3751_root_address_inst_ack_0 <= ptr_deref_3751_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3751_resized_base_address;
      ptr_deref_3751_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3756_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3756_addr_0_ack_0 <= ptr_deref_3756_addr_0_req_0;
      aggregated_sig <= ptr_deref_3756_root_address;
      ptr_deref_3756_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3756_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3756_gather_scatter_ack_0 <= ptr_deref_3756_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3756_data_0;
      iNsTr_6_3757 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3756_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3756_root_address_inst_ack_0 <= ptr_deref_3756_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3756_resized_base_address;
      ptr_deref_3756_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    -- shared load operator group (0) : ptr_deref_3756_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3756_load_0_req_0,
        ptr_deref_3756_load_0_ack_0,
        ptr_deref_3756_load_0_req_1,
        ptr_deref_3756_load_0_ack_1,
        "ptr_deref_3756_load_0",
        "memory_space_7" ,
        ptr_deref_3756_data_0,
        ptr_deref_3756_word_address_0,
        "ptr_deref_3756_data_0",
        "ptr_deref_3756_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3756_load_0_req_0;
      ptr_deref_3756_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3756_load_0_req_1;
      ptr_deref_3756_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3756_word_address_0;
      ptr_deref_3756_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_7_lr_req(0),
          mack => memory_space_7_lr_ack(0),
          maddr => memory_space_7_lr_addr(0 downto 0),
          mtag => memory_space_7_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_7_lc_req(0),
          mack => memory_space_7_lc_ack(0),
          mdata => memory_space_7_lc_data(31 downto 0),
          mtag => memory_space_7_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3751_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_7 address ptr_deref_3751_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3751_word_address_0) &  " data ptr_deref_3751_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3751_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3751_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_3751_store_0_req_0;
      ptr_deref_3751_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3751_store_0_req_1;
      ptr_deref_3751_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3751_word_address_0;
      data_in <= ptr_deref_3751_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_7_sr_req(0),
          mack => memory_space_7_sr_ack(0),
          maddr => memory_space_7_sr_addr(0 downto 0),
          mdata => memory_space_7_sr_data(31 downto 0),
          mtag => memory_space_7_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_7_sc_req(0),
          mack => memory_space_7_sc_ack(0),
          mtag => memory_space_7_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : simple_obj_ref_3748_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3748_inst_ack_0 then -- 
            assert false report " ReadPipe receive_packet_pipe to wire iNsTr_4_3749 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3748_inst_req_0;
      simple_obj_ref_3748_inst_ack_0 <= ack(0);
      iNsTr_4_3749 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => receive_packet_pipe_pipe_read_req(0),
          oack => receive_packet_pipe_pipe_read_ack(0),
          odata => receive_packet_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3758_inst_ack_0 then -- 
          assert false report " WritePipe src_in0 from wire iNsTr_6_3757 value="  &  convert_slv_to_hex_string(iNsTr_6_3757) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3758_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3758_inst_req_0;
      simple_obj_ref_3758_inst_ack_0 <= ack(0);
      data_in <= iNsTr_6_3757;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => src_in0_pipe_write_req(0),
          oack => src_in0_pipe_write_ack(0),
          odata => src_in0_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_3743_call 
    CallGroup0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3743_call_req_0;
      call_stmt_3743_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3743_call_req_1;
      call_stmt_3743_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => global_storage_initializer_x_call_reqs(0),
          ackR => global_storage_initializer_x_call_acks(0),
          tagR => global_storage_initializer_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => global_storage_initializer_x_return_acks(0), -- cross-over
          ackL => global_storage_initializer_x_return_reqs(0), -- cross-over
          tagL => global_storage_initializer_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_3744_call 
    CallGroup1: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= call_stmt_3744_call_req_0;
      call_stmt_3744_call_ack_0 <= ackL(0);
      reqR(0) <= call_stmt_3744_call_req_1;
      call_stmt_3744_call_ack_1 <= ackR(0);
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => free_queue_init_call_reqs(0),
          ackR => free_queue_init_call_acks(0),
          tagR => free_queue_init_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => free_queue_init_return_acks(0), -- cross-over
          ackL => free_queue_init_return_reqs(0), -- cross-over
          tagL => free_queue_init_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_7: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_7_lr_addr,
      lr_req_in => memory_space_7_lr_req,
      lr_ack_out => memory_space_7_lr_ack,
      lr_tag_in => memory_space_7_lr_tag,
      lc_req_in => memory_space_7_lc_req,
      lc_ack_out => memory_space_7_lc_ack,
      lc_data_out => memory_space_7_lc_data,
      lc_tag_out => memory_space_7_lc_tag,
      sr_addr_in => memory_space_7_sr_addr,
      sr_data_in => memory_space_7_sr_data,
      sr_req_in => memory_space_7_sr_req,
      sr_ack_out => memory_space_7_sr_ack,
      sr_tag_in => memory_space_7_sr_tag,
      sc_req_in=> memory_space_7_sc_req,
      sc_ack_out => memory_space_7_sc_ack,
      sc_tag_out => memory_space_7_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity wrapper_output is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    tofpga0_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga0_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga1_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga1_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga2_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga2_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga3_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga3_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
    tofpga_port_number_pipe_read_req : out  std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_read_ack : in   std_logic_vector(0 downto 0);
    tofpga_port_number_pipe_read_data : in   std_logic_vector(31 downto 0);
    send_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    send_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity wrapper_output;
architecture Default of wrapper_output is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal wrapper_output_CP_19386_start: Boolean;
  -- links between control-path and data-path
  signal simple_obj_ref_3848_inst_ack_0 : boolean;
  signal ptr_deref_3842_root_address_inst_req_0 : boolean;
  signal ptr_deref_3855_base_resize_req_0 : boolean;
  signal ptr_deref_3842_base_resize_req_0 : boolean;
  signal ptr_deref_3842_addr_0_req_0 : boolean;
  signal simple_obj_ref_3868_inst_req_0 : boolean;
  signal ptr_deref_3862_root_address_inst_req_0 : boolean;
  signal ptr_deref_3862_load_0_req_1 : boolean;
  signal ptr_deref_3862_root_address_inst_ack_0 : boolean;
  signal type_cast_3839_inst_ack_0 : boolean;
  signal ptr_deref_3842_addr_0_ack_0 : boolean;
  signal ptr_deref_3842_base_resize_ack_0 : boolean;
  signal ptr_deref_3829_store_0_req_1 : boolean;
  signal ptr_deref_3842_store_0_req_0 : boolean;
  signal simple_obj_ref_3868_inst_ack_0 : boolean;
  signal ptr_deref_3829_addr_0_req_0 : boolean;
  signal ptr_deref_3862_base_resize_req_0 : boolean;
  signal ptr_deref_3829_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3829_store_0_ack_1 : boolean;
  signal ptr_deref_3855_store_0_req_1 : boolean;
  signal simple_obj_ref_3848_inst_req_0 : boolean;
  signal ptr_deref_3862_load_0_ack_0 : boolean;
  signal ptr_deref_3842_root_address_inst_ack_0 : boolean;
  signal type_cast_3866_inst_req_0 : boolean;
  signal simple_obj_ref_3835_inst_req_0 : boolean;
  signal ptr_deref_3829_gather_scatter_req_0 : boolean;
  signal ptr_deref_3855_base_resize_ack_0 : boolean;
  signal ptr_deref_3855_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_3835_inst_ack_0 : boolean;
  signal ptr_deref_3829_root_address_inst_req_0 : boolean;
  signal type_cast_3839_inst_req_0 : boolean;
  signal ptr_deref_3842_gather_scatter_req_0 : boolean;
  signal type_cast_3826_inst_req_0 : boolean;
  signal ptr_deref_3829_addr_0_ack_0 : boolean;
  signal ptr_deref_3855_store_0_ack_1 : boolean;
  signal type_cast_3866_inst_ack_0 : boolean;
  signal ptr_deref_3862_gather_scatter_req_0 : boolean;
  signal ptr_deref_3842_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3862_base_resize_ack_0 : boolean;
  signal ptr_deref_3855_store_0_ack_0 : boolean;
  signal type_cast_3852_inst_ack_0 : boolean;
  signal ptr_deref_3862_gather_scatter_ack_0 : boolean;
  signal type_cast_3826_inst_ack_0 : boolean;
  signal type_cast_3852_inst_req_0 : boolean;
  signal ptr_deref_3855_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3842_store_0_ack_0 : boolean;
  signal ptr_deref_3855_addr_0_req_0 : boolean;
  signal ptr_deref_3855_addr_0_ack_0 : boolean;
  signal ptr_deref_3862_load_0_ack_1 : boolean;
  signal ptr_deref_3862_load_0_req_0 : boolean;
  signal ptr_deref_3829_store_0_req_0 : boolean;
  signal ptr_deref_3829_store_0_ack_0 : boolean;
  signal ptr_deref_3829_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3855_gather_scatter_req_0 : boolean;
  signal ptr_deref_3842_store_0_req_1 : boolean;
  signal ptr_deref_3855_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3842_store_0_ack_1 : boolean;
  signal ptr_deref_3855_store_0_req_0 : boolean;
  signal ptr_deref_3862_addr_0_ack_0 : boolean;
  signal ptr_deref_3829_base_resize_ack_0 : boolean;
  signal ptr_deref_3862_addr_0_req_0 : boolean;
  signal ptr_deref_3829_base_resize_req_0 : boolean;
  signal simple_obj_ref_3781_inst_req_0 : boolean;
  signal simple_obj_ref_3781_inst_ack_0 : boolean;
  signal ptr_deref_3784_base_resize_req_0 : boolean;
  signal ptr_deref_3784_base_resize_ack_0 : boolean;
  signal ptr_deref_3784_root_address_inst_req_0 : boolean;
  signal ptr_deref_3784_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3784_addr_0_req_0 : boolean;
  signal ptr_deref_3784_addr_0_ack_0 : boolean;
  signal ptr_deref_3784_gather_scatter_req_0 : boolean;
  signal ptr_deref_3784_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3784_store_0_req_0 : boolean;
  signal ptr_deref_3784_store_0_ack_0 : boolean;
  signal ptr_deref_3784_store_0_req_1 : boolean;
  signal ptr_deref_3784_store_0_ack_1 : boolean;
  signal ptr_deref_3789_base_resize_req_0 : boolean;
  signal ptr_deref_3789_base_resize_ack_0 : boolean;
  signal ptr_deref_3789_root_address_inst_req_0 : boolean;
  signal ptr_deref_3789_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3789_addr_0_req_0 : boolean;
  signal ptr_deref_3789_addr_0_ack_0 : boolean;
  signal ptr_deref_3789_load_0_req_0 : boolean;
  signal ptr_deref_3789_load_0_ack_0 : boolean;
  signal ptr_deref_3789_load_0_req_1 : boolean;
  signal ptr_deref_3789_load_0_ack_1 : boolean;
  signal ptr_deref_3789_gather_scatter_req_0 : boolean;
  signal ptr_deref_3789_gather_scatter_ack_0 : boolean;
  signal switch_stmt_3791_branch_default_req_0 : boolean;
  signal switch_stmt_3791_select_expr_0_req_0 : boolean;
  signal switch_stmt_3791_select_expr_0_ack_0 : boolean;
  signal switch_stmt_3791_select_expr_0_req_1 : boolean;
  signal switch_stmt_3791_select_expr_0_ack_1 : boolean;
  signal switch_stmt_3791_branch_0_req_0 : boolean;
  signal switch_stmt_3791_select_expr_1_req_0 : boolean;
  signal switch_stmt_3791_select_expr_1_ack_0 : boolean;
  signal switch_stmt_3791_select_expr_1_req_1 : boolean;
  signal switch_stmt_3791_select_expr_1_ack_1 : boolean;
  signal switch_stmt_3791_branch_1_req_0 : boolean;
  signal switch_stmt_3791_select_expr_2_req_0 : boolean;
  signal switch_stmt_3791_select_expr_2_ack_0 : boolean;
  signal switch_stmt_3791_select_expr_2_req_1 : boolean;
  signal switch_stmt_3791_select_expr_2_ack_1 : boolean;
  signal switch_stmt_3791_branch_2_req_0 : boolean;
  signal switch_stmt_3791_select_expr_3_req_0 : boolean;
  signal switch_stmt_3791_select_expr_3_ack_0 : boolean;
  signal switch_stmt_3791_select_expr_3_req_1 : boolean;
  signal switch_stmt_3791_select_expr_3_ack_1 : boolean;
  signal switch_stmt_3791_branch_3_req_0 : boolean;
  signal switch_stmt_3791_branch_0_ack_1 : boolean;
  signal switch_stmt_3791_branch_1_ack_1 : boolean;
  signal switch_stmt_3791_branch_2_ack_1 : boolean;
  signal switch_stmt_3791_branch_3_ack_1 : boolean;
  signal switch_stmt_3791_branch_default_ack_0 : boolean;
  signal simple_obj_ref_3809_inst_req_0 : boolean;
  signal simple_obj_ref_3809_inst_ack_0 : boolean;
  signal type_cast_3813_inst_req_0 : boolean;
  signal type_cast_3813_inst_ack_0 : boolean;
  signal ptr_deref_3816_base_resize_req_0 : boolean;
  signal ptr_deref_3816_base_resize_ack_0 : boolean;
  signal ptr_deref_3816_root_address_inst_req_0 : boolean;
  signal ptr_deref_3816_root_address_inst_ack_0 : boolean;
  signal ptr_deref_3816_addr_0_req_0 : boolean;
  signal ptr_deref_3816_addr_0_ack_0 : boolean;
  signal ptr_deref_3816_gather_scatter_req_0 : boolean;
  signal ptr_deref_3816_gather_scatter_ack_0 : boolean;
  signal ptr_deref_3816_store_0_req_0 : boolean;
  signal ptr_deref_3816_store_0_ack_0 : boolean;
  signal ptr_deref_3816_store_0_req_1 : boolean;
  signal ptr_deref_3816_store_0_ack_1 : boolean;
  signal simple_obj_ref_3822_inst_req_0 : boolean;
  signal simple_obj_ref_3822_inst_ack_0 : boolean;
  signal memory_space_8_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_lr_tag : std_logic_vector(5 downto 0);
  signal memory_space_8_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_8_lc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_8_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_8_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_8_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_8_sr_tag : std_logic_vector(5 downto 0);
  signal memory_space_8_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_8_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_8_sc_tag :  std_logic_vector(2 downto 0);
  signal memory_space_9_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_9_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_9_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_9_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_9_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_9_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_9_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_9_sc_tag :  std_logic_vector(0 downto 0);
  -- 
begin --  
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 1, backward_delay => 1) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  tagQueue: QueueBase generic map(data_width => 1, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  wrapper_output_CP_19386: Block -- control-path 
    signal cp_elements: BooleanArray(133 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(3);
    finAckJoin: join2 
    generic map ( bypass => false)
    port map(pred0 => fin_req_symbol, pred1 => cp_elements(3), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    cp_elements(1) <= cp_elements(26);
    cp_elements(2) <= OrReduce(cp_elements(47) & cp_elements(131));
    req_19626_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(2), ack => simple_obj_ref_3809_inst_req_0); -- 
    cp_elements(3) <= false; 
    ack_19450_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3781_inst_ack_0, ack => cp_elements(4)); -- 
    cp_elements(5) <= cp_elements(4);
    cp_elements(6) <= cp_elements(5);
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(6) & cp_elements(8) & cp_elements(12));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => ptr_deref_3784_gather_scatter_req_0); -- 
    cp_elements(8) <= cp_elements(5);
    cp_elements(9) <= cp_elements(8);
    base_resize_req_19467_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => ptr_deref_3784_base_resize_req_0); -- 
    base_resize_ack_19468_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3784_base_resize_ack_0, ack => cp_elements(10)); -- 
    sum_rename_req_19472_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => ptr_deref_3784_root_address_inst_req_0); -- 
    sum_rename_ack_19473_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3784_root_address_inst_ack_0, ack => cp_elements(11)); -- 
    root_rename_req_19477_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => ptr_deref_3784_addr_0_req_0); -- 
    root_rename_ack_19478_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3784_addr_0_ack_0, ack => cp_elements(12)); -- 
    split_ack_19483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3784_gather_scatter_ack_0, ack => cp_elements(13)); -- 
    rr_19490_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(13), ack => ptr_deref_3784_store_0_req_0); -- 
    cp_elements(14) <= ptr_deref_3784_store_0_ack_0;
    cp_elements(15) <= cp_elements(14);
    cr_19501_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => ptr_deref_3784_store_0_req_1); -- 
    ca_19502_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3784_store_0_ack_1, ack => cp_elements(16)); -- 
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(14) & cp_elements(18) & cp_elements(22));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    rr_19536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => ptr_deref_3789_load_0_req_0); -- 
    cp_elements(18) <= cp_elements(5);
    cp_elements(19) <= cp_elements(18);
    base_resize_req_19515_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => ptr_deref_3789_base_resize_req_0); -- 
    base_resize_ack_19516_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_base_resize_ack_0, ack => cp_elements(20)); -- 
    sum_rename_req_19520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => ptr_deref_3789_root_address_inst_req_0); -- 
    sum_rename_ack_19521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_root_address_inst_ack_0, ack => cp_elements(21)); -- 
    root_rename_req_19525_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(21), ack => ptr_deref_3789_addr_0_req_0); -- 
    root_rename_ack_19526_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_addr_0_ack_0, ack => cp_elements(22)); -- 
    ra_19537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_load_0_ack_0, ack => cp_elements(23)); -- 
    cr_19547_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(23), ack => ptr_deref_3789_load_0_req_1); -- 
    ca_19548_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_load_0_ack_1, ack => cp_elements(24)); -- 
    merge_req_19549_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(24), ack => ptr_deref_3789_gather_scatter_req_0); -- 
    merge_ack_19550_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3789_gather_scatter_ack_0, ack => cp_elements(25)); -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(16) & cp_elements(25));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    cp_elements(27) <= cp_elements(1);
    cp_elements(28) <= false;
    cp_elements(29) <= cp_elements(28);
    cp_elements(30) <= cp_elements(1);
    cp_elements(31) <= cp_elements(30);
    cp_elements(32) <= cp_elements(31);
    rr_19562_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => switch_stmt_3791_select_expr_0_req_0); -- 
    ra_19563_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_0_ack_0, ack => cp_elements(33)); -- 
    cr_19564_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(33), ack => switch_stmt_3791_select_expr_0_req_1); -- 
    ca_19565_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_0_ack_1, ack => cp_elements(34)); -- 
    cmp_19566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(34), ack => switch_stmt_3791_branch_0_req_0); -- 
    cp_elements(35) <= cp_elements(31);
    rr_19570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => switch_stmt_3791_select_expr_1_req_0); -- 
    ra_19571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_1_ack_0, ack => cp_elements(36)); -- 
    cr_19572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => switch_stmt_3791_select_expr_1_req_1); -- 
    ca_19573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_1_ack_1, ack => cp_elements(37)); -- 
    cmp_19574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => switch_stmt_3791_branch_1_req_0); -- 
    cp_elements(38) <= cp_elements(31);
    rr_19578_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => switch_stmt_3791_select_expr_2_req_0); -- 
    ra_19579_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_2_ack_0, ack => cp_elements(39)); -- 
    cr_19580_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(39), ack => switch_stmt_3791_select_expr_2_req_1); -- 
    ca_19581_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_2_ack_1, ack => cp_elements(40)); -- 
    cmp_19582_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => switch_stmt_3791_branch_2_req_0); -- 
    cp_elements(41) <= cp_elements(31);
    rr_19586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => switch_stmt_3791_select_expr_3_req_0); -- 
    ra_19587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_3_ack_0, ack => cp_elements(42)); -- 
    cr_19588_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(42), ack => switch_stmt_3791_select_expr_3_req_1); -- 
    ca_19589_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_select_expr_3_ack_1, ack => cp_elements(43)); -- 
    cmp_19590_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => switch_stmt_3791_branch_3_req_0); -- 
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(3 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(34) & cp_elements(37) & cp_elements(40) & cp_elements(43));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    Xexit_19558_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(44), ack => switch_stmt_3791_branch_default_req_0); -- 
    cp_elements(45) <= cp_elements(44);
    cp_elements(46) <= cp_elements(45);
    ack1_19595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_branch_0_ack_1, ack => cp_elements(47)); -- 
    cp_elements(48) <= cp_elements(45);
    ack1_19600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_branch_1_ack_1, ack => cp_elements(49)); -- 
    req_19699_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(49), ack => simple_obj_ref_3822_inst_req_0); -- 
    cp_elements(50) <= cp_elements(45);
    ack1_19605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_branch_2_ack_1, ack => cp_elements(51)); -- 
    req_19772_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(51), ack => simple_obj_ref_3835_inst_req_0); -- 
    cp_elements(52) <= cp_elements(45);
    ack1_19610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_branch_3_ack_1, ack => cp_elements(53)); -- 
    req_19845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => simple_obj_ref_3848_inst_req_0); -- 
    cp_elements(54) <= cp_elements(45);
    ack0_19615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => switch_stmt_3791_branch_default_ack_0, ack => cp_elements(55)); -- 
    ack_19627_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3809_inst_ack_0, ack => cp_elements(56)); -- 
    cp_elements(57) <= cp_elements(56);
    cpelement_group_58 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(59) & cp_elements(60));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(58),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(58), ack => type_cast_3813_inst_req_0); -- 
    cp_elements(59) <= cp_elements(57);
    cp_elements(60) <= cp_elements(57);
    ack_19640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3813_inst_ack_0, ack => cp_elements(61)); -- 
    cpelement_group_62 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(61) & cp_elements(63) & cp_elements(67));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(62),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19669_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(62), ack => ptr_deref_3816_gather_scatter_req_0); -- 
    cp_elements(63) <= cp_elements(57);
    cp_elements(64) <= cp_elements(63);
    base_resize_req_19654_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(64), ack => ptr_deref_3816_base_resize_req_0); -- 
    base_resize_ack_19655_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_base_resize_ack_0, ack => cp_elements(65)); -- 
    sum_rename_req_19659_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => ptr_deref_3816_root_address_inst_req_0); -- 
    sum_rename_ack_19660_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_root_address_inst_ack_0, ack => cp_elements(66)); -- 
    root_rename_req_19664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => ptr_deref_3816_addr_0_req_0); -- 
    root_rename_ack_19665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_addr_0_ack_0, ack => cp_elements(67)); -- 
    split_ack_19670_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_gather_scatter_ack_0, ack => cp_elements(68)); -- 
    rr_19677_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(68), ack => ptr_deref_3816_store_0_req_0); -- 
    ra_19678_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_store_0_ack_0, ack => cp_elements(69)); -- 
    cr_19688_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(69), ack => ptr_deref_3816_store_0_req_1); -- 
    ca_19689_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3816_store_0_ack_1, ack => cp_elements(70)); -- 
    ack_19700_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3822_inst_ack_0, ack => cp_elements(71)); -- 
    cp_elements(72) <= cp_elements(71);
    cpelement_group_73 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(74) & cp_elements(75));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(73),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19712_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => type_cast_3826_inst_req_0); -- 
    cp_elements(74) <= cp_elements(72);
    cp_elements(75) <= cp_elements(72);
    ack_19713_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3826_inst_ack_0, ack => cp_elements(76)); -- 
    cpelement_group_77 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(76) & cp_elements(78) & cp_elements(82));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(77),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_3829_gather_scatter_req_0); -- 
    cp_elements(78) <= cp_elements(72);
    cp_elements(79) <= cp_elements(78);
    base_resize_req_19727_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_3829_base_resize_req_0); -- 
    base_resize_ack_19728_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_base_resize_ack_0, ack => cp_elements(80)); -- 
    sum_rename_req_19732_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_3829_root_address_inst_req_0); -- 
    sum_rename_ack_19733_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_root_address_inst_ack_0, ack => cp_elements(81)); -- 
    root_rename_req_19737_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_3829_addr_0_req_0); -- 
    root_rename_ack_19738_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_addr_0_ack_0, ack => cp_elements(82)); -- 
    split_ack_19743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_gather_scatter_ack_0, ack => cp_elements(83)); -- 
    rr_19750_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(83), ack => ptr_deref_3829_store_0_req_0); -- 
    ra_19751_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_store_0_ack_0, ack => cp_elements(84)); -- 
    cr_19761_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(84), ack => ptr_deref_3829_store_0_req_1); -- 
    ca_19762_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3829_store_0_ack_1, ack => cp_elements(85)); -- 
    ack_19773_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3835_inst_ack_0, ack => cp_elements(86)); -- 
    cp_elements(87) <= cp_elements(86);
    cpelement_group_88 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(89) & cp_elements(90));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(88),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => type_cast_3839_inst_req_0); -- 
    cp_elements(89) <= cp_elements(87);
    cp_elements(90) <= cp_elements(87);
    ack_19786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3839_inst_ack_0, ack => cp_elements(91)); -- 
    cpelement_group_92 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(91) & cp_elements(93) & cp_elements(97));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(92),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19815_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(92), ack => ptr_deref_3842_gather_scatter_req_0); -- 
    cp_elements(93) <= cp_elements(87);
    cp_elements(94) <= cp_elements(93);
    base_resize_req_19800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => ptr_deref_3842_base_resize_req_0); -- 
    base_resize_ack_19801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_base_resize_ack_0, ack => cp_elements(95)); -- 
    sum_rename_req_19805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => ptr_deref_3842_root_address_inst_req_0); -- 
    sum_rename_ack_19806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_root_address_inst_ack_0, ack => cp_elements(96)); -- 
    root_rename_req_19810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(96), ack => ptr_deref_3842_addr_0_req_0); -- 
    root_rename_ack_19811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_addr_0_ack_0, ack => cp_elements(97)); -- 
    split_ack_19816_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_gather_scatter_ack_0, ack => cp_elements(98)); -- 
    rr_19823_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(98), ack => ptr_deref_3842_store_0_req_0); -- 
    ra_19824_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_store_0_ack_0, ack => cp_elements(99)); -- 
    cr_19834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(99), ack => ptr_deref_3842_store_0_req_1); -- 
    ca_19835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3842_store_0_ack_1, ack => cp_elements(100)); -- 
    ack_19846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3848_inst_ack_0, ack => cp_elements(101)); -- 
    cp_elements(102) <= cp_elements(101);
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(104) & cp_elements(105));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19858_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(103), ack => type_cast_3852_inst_req_0); -- 
    cp_elements(104) <= cp_elements(102);
    cp_elements(105) <= cp_elements(102);
    ack_19859_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3852_inst_ack_0, ack => cp_elements(106)); -- 
    cpelement_group_107 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(106) & cp_elements(108) & cp_elements(112));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(107),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_19888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => ptr_deref_3855_gather_scatter_req_0); -- 
    cp_elements(108) <= cp_elements(102);
    cp_elements(109) <= cp_elements(108);
    base_resize_req_19873_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(109), ack => ptr_deref_3855_base_resize_req_0); -- 
    base_resize_ack_19874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_base_resize_ack_0, ack => cp_elements(110)); -- 
    sum_rename_req_19878_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(110), ack => ptr_deref_3855_root_address_inst_req_0); -- 
    sum_rename_ack_19879_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_root_address_inst_ack_0, ack => cp_elements(111)); -- 
    root_rename_req_19883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(111), ack => ptr_deref_3855_addr_0_req_0); -- 
    root_rename_ack_19884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_addr_0_ack_0, ack => cp_elements(112)); -- 
    split_ack_19889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_gather_scatter_ack_0, ack => cp_elements(113)); -- 
    rr_19896_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(113), ack => ptr_deref_3855_store_0_req_0); -- 
    ra_19897_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_store_0_ack_0, ack => cp_elements(114)); -- 
    cr_19907_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => ptr_deref_3855_store_0_req_1); -- 
    ca_19908_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3855_store_0_ack_1, ack => cp_elements(115)); -- 
    cp_elements(116) <= cp_elements(133);
    cp_elements(117) <= cp_elements(116);
    base_resize_req_19924_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(117), ack => ptr_deref_3862_base_resize_req_0); -- 
    base_resize_ack_19925_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_base_resize_ack_0, ack => cp_elements(118)); -- 
    sum_rename_req_19929_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => ptr_deref_3862_root_address_inst_req_0); -- 
    sum_rename_ack_19930_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_root_address_inst_ack_0, ack => cp_elements(119)); -- 
    root_rename_req_19934_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(119), ack => ptr_deref_3862_addr_0_req_0); -- 
    root_rename_ack_19935_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_addr_0_ack_0, ack => cp_elements(120)); -- 
    rr_19945_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => ptr_deref_3862_load_0_req_0); -- 
    ra_19946_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_load_0_ack_0, ack => cp_elements(121)); -- 
    cr_19956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(121), ack => ptr_deref_3862_load_0_req_1); -- 
    ca_19957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_load_0_ack_1, ack => cp_elements(122)); -- 
    merge_req_19958_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => ptr_deref_3862_gather_scatter_req_0); -- 
    merge_ack_19959_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_3862_gather_scatter_ack_0, ack => cp_elements(123)); -- 
    cpelement_group_124 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors <= (cp_elements(123) & cp_elements(125));
      jNoI: join -- 
        generic map ( bypass => false)
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(124),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    req_19968_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => type_cast_3866_inst_req_0); -- 
    cp_elements(125) <= cp_elements(116);
    ack_19969_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_3866_inst_ack_0, ack => cp_elements(126)); -- 
    pipe_wreq_19980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => simple_obj_ref_3868_inst_req_0); -- 
    pipe_wack_19981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_3868_inst_ack_0, ack => cp_elements(127)); -- 
    cp_elements(128) <= OrReduce(cp_elements(0) & cp_elements(127));
    cp_elements(129) <= cp_elements(128);
    req_19449_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(129), ack => simple_obj_ref_3781_inst_req_0); -- 
    cp_elements(130) <= false;
    cp_elements(131) <= cp_elements(130);
    cp_elements(132) <= OrReduce(cp_elements(55) & cp_elements(70) & cp_elements(85) & cp_elements(100) & cp_elements(115));
    cp_elements(133) <= cp_elements(132);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal expr_3793_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3793_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3796_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3796_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3799_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3799_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal expr_3802_wire_constant : std_logic_vector(31 downto 0);
    signal expr_3802_wire_constant_cmp : std_logic_vector(0 downto 0);
    signal iNsTr_12_3810 : std_logic_vector(31 downto 0);
    signal iNsTr_13_3814 : std_logic_vector(31 downto 0);
    signal iNsTr_17_3823 : std_logic_vector(31 downto 0);
    signal iNsTr_18_3827 : std_logic_vector(31 downto 0);
    signal iNsTr_22_3836 : std_logic_vector(31 downto 0);
    signal iNsTr_23_3840 : std_logic_vector(31 downto 0);
    signal iNsTr_27_3849 : std_logic_vector(31 downto 0);
    signal iNsTr_28_3853 : std_logic_vector(31 downto 0);
    signal iNsTr_2_3782 : std_logic_vector(31 downto 0);
    signal iNsTr_4_3790 : std_logic_vector(31 downto 0);
    signal iNsTr_6_3863 : std_logic_vector(31 downto 0);
    signal iNsTr_7_3867 : std_logic_vector(31 downto 0);
    signal pkt_3773 : std_logic_vector(31 downto 0);
    signal port_number_3777 : std_logic_vector(31 downto 0);
    signal ptr_deref_3784_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3784_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3784_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3784_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3784_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3784_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3789_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3789_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3789_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3789_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3789_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3816_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3816_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3816_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3816_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3816_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3816_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3829_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3829_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3829_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3829_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3829_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3829_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3842_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3842_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3842_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3842_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3842_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3842_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3855_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3855_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3855_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3855_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_3855_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3855_word_offset_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3862_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_3862_resized_base_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3862_root_address : std_logic_vector(0 downto 0);
    signal ptr_deref_3862_word_address_0 : std_logic_vector(0 downto 0);
    signal ptr_deref_3862_word_offset_0 : std_logic_vector(0 downto 0);
    signal xxwrapper_outputxxbodyxxpkt_alloc_base_address : std_logic_vector(0 downto 0);
    signal xxwrapper_outputxxbodyxxport_number_alloc_base_address : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    expr_3793_wire_constant <= "00000000000000000000000000000001";
    expr_3796_wire_constant <= "00000000000000000000000000000010";
    expr_3799_wire_constant <= "00000000000000000000000000000011";
    expr_3802_wire_constant <= "00000000000000000000000000000100";
    pkt_3773 <= "00000000000000000000000000000000";
    port_number_3777 <= "00000000000000000000000000000000";
    ptr_deref_3784_word_offset_0 <= "0";
    ptr_deref_3789_word_offset_0 <= "0";
    ptr_deref_3816_word_offset_0 <= "0";
    ptr_deref_3829_word_offset_0 <= "0";
    ptr_deref_3842_word_offset_0 <= "0";
    ptr_deref_3855_word_offset_0 <= "0";
    ptr_deref_3862_word_offset_0 <= "0";
    xxwrapper_outputxxbodyxxpkt_alloc_base_address <= "0";
    xxwrapper_outputxxbodyxxport_number_alloc_base_address <= "0";
    ptr_deref_3784_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => port_number_3777, dout => ptr_deref_3784_resized_base_address, req => ptr_deref_3784_base_resize_req_0, ack => ptr_deref_3784_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3789_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => port_number_3777, dout => ptr_deref_3789_resized_base_address, req => ptr_deref_3789_base_resize_req_0, ack => ptr_deref_3789_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3816_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3773, dout => ptr_deref_3816_resized_base_address, req => ptr_deref_3816_base_resize_req_0, ack => ptr_deref_3816_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3829_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3773, dout => ptr_deref_3829_resized_base_address, req => ptr_deref_3829_base_resize_req_0, ack => ptr_deref_3829_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3842_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3773, dout => ptr_deref_3842_resized_base_address, req => ptr_deref_3842_base_resize_req_0, ack => ptr_deref_3842_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3855_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3773, dout => ptr_deref_3855_resized_base_address, req => ptr_deref_3855_base_resize_req_0, ack => ptr_deref_3855_base_resize_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3862_base_resize: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 1, flow_through => true ) 
      port map( din => pkt_3773, dout => ptr_deref_3862_resized_base_address, req => ptr_deref_3862_base_resize_req_0, ack => ptr_deref_3862_base_resize_ack_0, clk => clk, reset => reset); -- 
    type_cast_3813_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_12_3810, dout => iNsTr_13_3814, req => type_cast_3813_inst_req_0, ack => type_cast_3813_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3826_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_17_3823, dout => iNsTr_18_3827, req => type_cast_3826_inst_req_0, ack => type_cast_3826_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3839_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_22_3836, dout => iNsTr_23_3840, req => type_cast_3839_inst_req_0, ack => type_cast_3839_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3852_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_27_3849, dout => iNsTr_28_3853, req => type_cast_3852_inst_req_0, ack => type_cast_3852_inst_ack_0, clk => clk, reset => reset); -- 
    type_cast_3866_inst: RegisterBase --
      generic map(in_data_width => 32,out_data_width => 32, flow_through => false ) 
      port map( din => iNsTr_6_3863, dout => iNsTr_7_3867, req => type_cast_3866_inst_req_0, ack => type_cast_3866_inst_ack_0, clk => clk, reset => reset); -- 
    ptr_deref_3784_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3784_addr_0_ack_0 <= ptr_deref_3784_addr_0_req_0;
      aggregated_sig <= ptr_deref_3784_root_address;
      ptr_deref_3784_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3784_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3784_gather_scatter_ack_0 <= ptr_deref_3784_gather_scatter_req_0;
      aggregated_sig <= iNsTr_2_3782;
      ptr_deref_3784_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3784_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3784_root_address_inst_ack_0 <= ptr_deref_3784_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3784_resized_base_address;
      ptr_deref_3784_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3789_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3789_addr_0_ack_0 <= ptr_deref_3789_addr_0_req_0;
      aggregated_sig <= ptr_deref_3789_root_address;
      ptr_deref_3789_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3789_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3789_gather_scatter_ack_0 <= ptr_deref_3789_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3789_data_0;
      iNsTr_4_3790 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3789_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3789_root_address_inst_ack_0 <= ptr_deref_3789_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3789_resized_base_address;
      ptr_deref_3789_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3816_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3816_addr_0_ack_0 <= ptr_deref_3816_addr_0_req_0;
      aggregated_sig <= ptr_deref_3816_root_address;
      ptr_deref_3816_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3816_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3816_gather_scatter_ack_0 <= ptr_deref_3816_gather_scatter_req_0;
      aggregated_sig <= iNsTr_13_3814;
      ptr_deref_3816_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3816_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3816_root_address_inst_ack_0 <= ptr_deref_3816_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3816_resized_base_address;
      ptr_deref_3816_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3829_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3829_addr_0_ack_0 <= ptr_deref_3829_addr_0_req_0;
      aggregated_sig <= ptr_deref_3829_root_address;
      ptr_deref_3829_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3829_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3829_gather_scatter_ack_0 <= ptr_deref_3829_gather_scatter_req_0;
      aggregated_sig <= iNsTr_18_3827;
      ptr_deref_3829_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3829_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3829_root_address_inst_ack_0 <= ptr_deref_3829_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3829_resized_base_address;
      ptr_deref_3829_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3842_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3842_addr_0_ack_0 <= ptr_deref_3842_addr_0_req_0;
      aggregated_sig <= ptr_deref_3842_root_address;
      ptr_deref_3842_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3842_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3842_gather_scatter_ack_0 <= ptr_deref_3842_gather_scatter_req_0;
      aggregated_sig <= iNsTr_23_3840;
      ptr_deref_3842_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3842_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3842_root_address_inst_ack_0 <= ptr_deref_3842_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3842_resized_base_address;
      ptr_deref_3842_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3855_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3855_addr_0_ack_0 <= ptr_deref_3855_addr_0_req_0;
      aggregated_sig <= ptr_deref_3855_root_address;
      ptr_deref_3855_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3855_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3855_gather_scatter_ack_0 <= ptr_deref_3855_gather_scatter_req_0;
      aggregated_sig <= iNsTr_28_3853;
      ptr_deref_3855_data_0 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3855_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3855_root_address_inst_ack_0 <= ptr_deref_3855_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3855_resized_base_address;
      ptr_deref_3855_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3862_addr_0: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3862_addr_0_ack_0 <= ptr_deref_3862_addr_0_req_0;
      aggregated_sig <= ptr_deref_3862_root_address;
      ptr_deref_3862_word_address_0 <= aggregated_sig(0 downto 0);
      --
    end Block;
    ptr_deref_3862_gather_scatter: Block -- 
      signal aggregated_sig: std_logic_vector(31 downto 0); --
    begin -- 
      ptr_deref_3862_gather_scatter_ack_0 <= ptr_deref_3862_gather_scatter_req_0;
      aggregated_sig <= ptr_deref_3862_data_0;
      iNsTr_6_3863 <= aggregated_sig(31 downto 0);
      --
    end Block;
    ptr_deref_3862_root_address_inst: Block -- 
      signal aggregated_sig: std_logic_vector(0 downto 0); --
    begin -- 
      ptr_deref_3862_root_address_inst_ack_0 <= ptr_deref_3862_root_address_inst_req_0;
      aggregated_sig <= ptr_deref_3862_resized_base_address;
      ptr_deref_3862_root_address <= aggregated_sig(0 downto 0);
      --
    end Block;
    switch_stmt_3791_branch_0: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3793_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3791_branch_0_req_0,
          ack0 => open,
          ack1 => switch_stmt_3791_branch_0_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3791_branch_1: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3796_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3791_branch_1_req_0,
          ack0 => open,
          ack1 => switch_stmt_3791_branch_1_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3791_branch_2: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3799_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3791_branch_2_req_0,
          ack0 => open,
          ack1 => switch_stmt_3791_branch_2_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3791_branch_3: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= expr_3802_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3791_branch_3_req_0,
          ack0 => open,
          ack1 => switch_stmt_3791_branch_3_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    switch_stmt_3791_branch_default: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(3 downto 0);
      begin 
      condition_sig <= expr_3793_wire_constant_cmp & expr_3796_wire_constant_cmp & expr_3799_wire_constant_cmp & expr_3802_wire_constant_cmp;
      branch_instance: BranchBase -- 
        generic map( condition_width => 4)
        port map( -- 
          condition => condition_sig,
          req => switch_stmt_3791_branch_default_req_0,
          ack0 => switch_stmt_3791_branch_default_ack_0,
          ack1 => open,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : switch_stmt_3791_select_expr_0 
    SplitOperatorGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3790;
      expr_3793_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3791_select_expr_0_req_0,
          ackL => switch_stmt_3791_select_expr_0_ack_0,
          reqR => switch_stmt_3791_select_expr_0_req_1,
          ackR => switch_stmt_3791_select_expr_0_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- shared split operator group (1) : switch_stmt_3791_select_expr_1 
    SplitOperatorGroup1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3790;
      expr_3796_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3791_select_expr_1_req_0,
          ackL => switch_stmt_3791_select_expr_1_ack_0,
          reqR => switch_stmt_3791_select_expr_1_req_1,
          ackR => switch_stmt_3791_select_expr_1_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : switch_stmt_3791_select_expr_2 
    SplitOperatorGroup2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3790;
      expr_3799_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3791_select_expr_2_req_0,
          ackL => switch_stmt_3791_select_expr_2_ack_0,
          reqR => switch_stmt_3791_select_expr_2_req_1,
          ackR => switch_stmt_3791_select_expr_2_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : switch_stmt_3791_select_expr_3 
    SplitOperatorGroup3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_4_3790;
      expr_3802_wire_constant_cmp <= data_out(0 downto 0);
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true,
          zero_delay => false, 
          flow_through => false--
        ) 
        port map ( -- 
          reqL => switch_stmt_3791_select_expr_3_req_0,
          ackL => switch_stmt_3791_select_expr_3_ack_0,
          reqR => switch_stmt_3791_select_expr_3_req_1,
          ackR => switch_stmt_3791_select_expr_3_ack_1,
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- shared load operator group (0) : ptr_deref_3789_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3789_load_0_req_0,
        ptr_deref_3789_load_0_ack_0,
        ptr_deref_3789_load_0_req_1,
        ptr_deref_3789_load_0_ack_1,
        "ptr_deref_3789_load_0",
        "memory_space_9" ,
        ptr_deref_3789_data_0,
        ptr_deref_3789_word_address_0,
        "ptr_deref_3789_data_0",
        "ptr_deref_3789_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3789_load_0_req_0;
      ptr_deref_3789_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3789_load_0_req_1;
      ptr_deref_3789_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3789_word_address_0;
      ptr_deref_3789_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_9_lr_req(0),
          mack => memory_space_9_lr_ack(0),
          maddr => memory_space_9_lr_addr(0 downto 0),
          mtag => memory_space_9_lr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 1,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_9_lc_req(0),
          mack => memory_space_9_lc_ack(0),
          mdata => memory_space_9_lc_data(31 downto 0),
          mtag => memory_space_9_lc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared load operator group (1) : ptr_deref_3862_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, -- 
        ptr_deref_3862_load_0_req_0,
        ptr_deref_3862_load_0_ack_0,
        ptr_deref_3862_load_0_req_1,
        ptr_deref_3862_load_0_ack_1,
        "ptr_deref_3862_load_0",
        "memory_space_8" ,
        ptr_deref_3862_data_0,
        ptr_deref_3862_word_address_0,
        "ptr_deref_3862_data_0",
        "ptr_deref_3862_word_address_0" -- 
      );
      reqL(0) <= ptr_deref_3862_load_0_req_0;
      ptr_deref_3862_load_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3862_load_0_req_1;
      ptr_deref_3862_load_0_ack_1 <= ackR(0);
      data_in <= ptr_deref_3862_word_address_0;
      ptr_deref_3862_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 1,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_8_lr_req(0),
          mack => memory_space_8_lr_ack(0),
          maddr => memory_space_8_lr_addr(0 downto 0),
          mtag => memory_space_8_lr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 3,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_8_lc_req(0),
          mack => memory_space_8_lc_ack(0),
          mdata => memory_space_8_lc_data(31 downto 0),
          mtag => memory_space_8_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3784_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_9 address ptr_deref_3784_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3784_word_address_0) &  " data ptr_deref_3784_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3784_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (0) : ptr_deref_3784_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(0 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      reqL(0) <= ptr_deref_3784_store_0_req_0;
      ptr_deref_3784_store_0_ack_0 <= ackL(0);
      reqR(0) <= ptr_deref_3784_store_0_req_1;
      ptr_deref_3784_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3784_word_address_0;
      data_in <= ptr_deref_3784_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 1,
        tag_length => 1,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_9_sr_req(0),
          mack => memory_space_9_sr_ack(0),
          maddr => memory_space_9_sr_addr(0 downto 0),
          mdata => memory_space_9_sr_data(31 downto 0),
          mtag => memory_space_9_sr_tag(3 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 1 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_9_sc_req(0),
          mack => memory_space_9_sc_ack(0),
          mtag => memory_space_9_sc_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if ptr_deref_3829_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3829_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3829_word_address_0) &  " data ptr_deref_3829_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3829_data_0) severity note; --
        end if;
        if ptr_deref_3816_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3816_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3816_word_address_0) &  " data ptr_deref_3816_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3816_data_0) severity note; --
        end if;
        if ptr_deref_3842_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3842_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3842_word_address_0) &  " data ptr_deref_3842_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3842_data_0) severity note; --
        end if;
        if ptr_deref_3855_store_0_ack_1 then -- 
          assert false report " WriteMem  memory_space_8 address ptr_deref_3855_word_address_0 ="  &  convert_slv_to_hex_string(ptr_deref_3855_word_address_0) &  " data ptr_deref_3855_data_0 ="  &  convert_slv_to_hex_string(ptr_deref_3855_data_0) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared store operator group (1) : ptr_deref_3829_store_0 ptr_deref_3816_store_0 ptr_deref_3842_store_0 ptr_deref_3855_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(3 downto 0);
      signal data_in: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      -- 
    begin -- 
      reqL(3) <= ptr_deref_3829_store_0_req_0;
      reqL(2) <= ptr_deref_3816_store_0_req_0;
      reqL(1) <= ptr_deref_3842_store_0_req_0;
      reqL(0) <= ptr_deref_3855_store_0_req_0;
      ptr_deref_3829_store_0_ack_0 <= ackL(3);
      ptr_deref_3816_store_0_ack_0 <= ackL(2);
      ptr_deref_3842_store_0_ack_0 <= ackL(1);
      ptr_deref_3855_store_0_ack_0 <= ackL(0);
      reqR(3) <= ptr_deref_3829_store_0_req_1;
      reqR(2) <= ptr_deref_3816_store_0_req_1;
      reqR(1) <= ptr_deref_3842_store_0_req_1;
      reqR(0) <= ptr_deref_3855_store_0_req_1;
      ptr_deref_3829_store_0_ack_1 <= ackR(3);
      ptr_deref_3816_store_0_ack_1 <= ackR(2);
      ptr_deref_3842_store_0_ack_1 <= ackR(1);
      ptr_deref_3855_store_0_ack_1 <= ackR(0);
      addr_in <= ptr_deref_3829_word_address_0 & ptr_deref_3816_word_address_0 & ptr_deref_3842_word_address_0 & ptr_deref_3855_word_address_0;
      data_in <= ptr_deref_3829_data_0 & ptr_deref_3816_data_0 & ptr_deref_3842_data_0 & ptr_deref_3855_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 1,
        data_width => 32,
        num_reqs => 4,
        tag_length => 3,
        time_stamp_width => 3,
        min_clock_period => true,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_8_sr_req(0),
          mack => memory_space_8_sr_ack(0),
          maddr => memory_space_8_sr_addr(0 downto 0),
          mdata => memory_space_8_sr_data(31 downto 0),
          mtag => memory_space_8_sr_tag(5 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 4,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_8_sc_req(0),
          mack => memory_space_8_sc_ack(0),
          mtag => memory_space_8_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    -- shared inport operator group (0) : simple_obj_ref_3781_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3781_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga_port_number to wire iNsTr_2_3782 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3781_inst_req_0;
      simple_obj_ref_3781_inst_ack_0 <= ack(0);
      iNsTr_2_3782 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga_port_number_pipe_read_req(0),
          oack => tofpga_port_number_pipe_read_ack(0),
          odata => tofpga_port_number_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : simple_obj_ref_3809_inst 
    InportGroup1: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3809_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga0_out0 to wire iNsTr_12_3810 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3809_inst_req_0;
      simple_obj_ref_3809_inst_ack_0 <= ack(0);
      iNsTr_12_3810 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga0_out0_pipe_read_req(0),
          oack => tofpga0_out0_pipe_read_ack(0),
          odata => tofpga0_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : simple_obj_ref_3822_inst 
    InportGroup2: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3822_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga1_out0 to wire iNsTr_17_3823 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3822_inst_req_0;
      simple_obj_ref_3822_inst_ack_0 <= ack(0);
      iNsTr_17_3823 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga1_out0_pipe_read_req(0),
          oack => tofpga1_out0_pipe_read_ack(0),
          odata => tofpga1_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared inport operator group (3) : simple_obj_ref_3835_inst 
    InportGroup3: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3835_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga2_out0 to wire iNsTr_22_3836 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3835_inst_req_0;
      simple_obj_ref_3835_inst_ack_0 <= ack(0);
      iNsTr_22_3836 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga2_out0_pipe_read_req(0),
          oack => tofpga2_out0_pipe_read_ack(0),
          odata => tofpga2_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 3
    -- shared inport operator group (4) : simple_obj_ref_3848_inst 
    InportGroup4: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_3848_inst_ack_0 then -- 
            assert false report " ReadPipe tofpga3_out0 to wire iNsTr_27_3849 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req(0) <= simple_obj_ref_3848_inst_req_0;
      simple_obj_ref_3848_inst_ack_0 <= ack(0);
      iNsTr_27_3849 <= data_out(31 downto 0);
      Inport: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => tofpga3_out0_pipe_read_req(0),
          oack => tofpga3_out0_pipe_read_ack(0),
          odata => tofpga3_out0_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 4
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_3868_inst_ack_0 then -- 
          assert false report " WritePipe send_packet_pipe from wire iNsTr_7_3867 value="  &  convert_slv_to_hex_string(iNsTr_7_3867) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_3868_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      -- 
    begin -- 
      req(0) <= simple_obj_ref_3868_inst_req_0;
      simple_obj_ref_3868_inst_ack_0 <= ack(0);
      data_in <= iNsTr_7_3867;
      outport: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => send_packet_pipe_pipe_write_req(0),
          oack => send_packet_pipe_pipe_write_ack(0),
          odata => send_packet_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  MemorySpace_memory_space_8: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_8_lr_addr,
      lr_req_in => memory_space_8_lr_req,
      lr_ack_out => memory_space_8_lr_ack,
      lr_tag_in => memory_space_8_lr_tag,
      lc_req_in => memory_space_8_lc_req,
      lc_ack_out => memory_space_8_lc_ack,
      lc_data_out => memory_space_8_lc_data,
      lc_tag_out => memory_space_8_lc_tag,
      sr_addr_in => memory_space_8_sr_addr,
      sr_data_in => memory_space_8_sr_data,
      sr_req_in => memory_space_8_sr_req,
      sr_ack_out => memory_space_8_sr_ack,
      sr_tag_in => memory_space_8_sr_tag,
      sc_req_in=> memory_space_8_sc_req,
      sc_ack_out => memory_space_8_sc_ack,
      sc_tag_out => memory_space_8_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_9: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_9_lr_addr,
      lr_req_in => memory_space_9_lr_req,
      lr_ack_out => memory_space_9_lr_ack,
      lr_tag_in => memory_space_9_lr_tag,
      lc_req_in => memory_space_9_lc_req,
      lc_ack_out => memory_space_9_lc_ack,
      lc_data_out => memory_space_9_lc_data,
      lc_tag_out => memory_space_9_lc_tag,
      sr_addr_in => memory_space_9_sr_addr,
      sr_data_in => memory_space_9_sr_data,
      sr_req_in => memory_space_9_sr_req,
      sr_ack_out => memory_space_9_sr_ack,
      sr_tag_in => memory_space_9_sr_tag,
      sc_req_in=> memory_space_9_sc_req,
      sc_ack_out => memory_space_9_sc_ack,
      sc_tag_out => memory_space_9_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
    in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
    in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
    in_data_pipe_write_data: in std_logic_vector(63 downto 0);
    in_data_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
    out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
    out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_read_data: out std_logic_vector(63 downto 0);
    out_data_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(8 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(4 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(4 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_3
  signal memory_space_3_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_lr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_lr_tag : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_lc_data : std_logic_vector(7 downto 0);
  signal memory_space_3_lc_tag :  std_logic_vector(4 downto 0);
  signal memory_space_3_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_3_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_3_sr_addr : std_logic_vector(13 downto 0);
  signal memory_space_3_sr_data : std_logic_vector(7 downto 0);
  signal memory_space_3_sr_tag : std_logic_vector(7 downto 0);
  signal memory_space_3_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_3_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_3_sc_tag :  std_logic_vector(4 downto 0);
  -- interface signals to connect to memory space memory_space_4
  signal memory_space_4_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_lr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_4_lc_tag :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_4_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_addr : std_logic_vector(0 downto 0);
  signal memory_space_4_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_4_sr_tag : std_logic_vector(3 downto 0);
  signal memory_space_4_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_4_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_4_sc_tag :  std_logic_vector(0 downto 0);
  -- interface signals to connect to memory space memory_space_5
  signal memory_space_5_lr_req :  std_logic_vector(9 downto 0);
  signal memory_space_5_lr_ack : std_logic_vector(9 downto 0);
  signal memory_space_5_lr_addr : std_logic_vector(159 downto 0);
  signal memory_space_5_lr_tag : std_logic_vector(109 downto 0);
  signal memory_space_5_lc_req : std_logic_vector(9 downto 0);
  signal memory_space_5_lc_ack :  std_logic_vector(9 downto 0);
  signal memory_space_5_lc_data : std_logic_vector(79 downto 0);
  signal memory_space_5_lc_tag :  std_logic_vector(49 downto 0);
  signal memory_space_5_sr_req :  std_logic_vector(7 downto 0);
  signal memory_space_5_sr_ack : std_logic_vector(7 downto 0);
  signal memory_space_5_sr_addr : std_logic_vector(127 downto 0);
  signal memory_space_5_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_5_sr_tag : std_logic_vector(87 downto 0);
  signal memory_space_5_sc_req : std_logic_vector(7 downto 0);
  signal memory_space_5_sc_ack :  std_logic_vector(7 downto 0);
  signal memory_space_5_sc_tag :  std_logic_vector(39 downto 0);
  -- declarations related to module GV_15_initializer_in_click_bc
  component GV_15_initializer_in_click_bc is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module GV_15_initializer_in_click_bc
  signal GV_15_initializer_in_click_bc_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal GV_15_initializer_in_click_bc_tag_out   : std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_start_req : std_logic;
  signal GV_15_initializer_in_click_bc_start_ack : std_logic;
  signal GV_15_initializer_in_click_bc_fin_req   : std_logic;
  signal GV_15_initializer_in_click_bc_fin_ack : std_logic;
  -- caller side aggregated signals for module GV_15_initializer_in_click_bc
  signal GV_15_initializer_in_click_bc_call_reqs: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_call_acks: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_reqs: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_acks: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_call_tag: std_logic_vector(0 downto 0);
  signal GV_15_initializer_in_click_bc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module GV_16_initializer_in_click_bc
  component GV_16_initializer_in_click_bc is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(4 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module GV_16_initializer_in_click_bc
  signal GV_16_initializer_in_click_bc_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal GV_16_initializer_in_click_bc_tag_out   : std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_start_req : std_logic;
  signal GV_16_initializer_in_click_bc_start_ack : std_logic;
  signal GV_16_initializer_in_click_bc_fin_req   : std_logic;
  signal GV_16_initializer_in_click_bc_fin_ack : std_logic;
  -- caller side aggregated signals for module GV_16_initializer_in_click_bc
  signal GV_16_initializer_in_click_bc_call_reqs: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_call_acks: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_reqs: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_acks: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_call_tag: std_logic_vector(0 downto 0);
  signal GV_16_initializer_in_click_bc_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module ahir_glue_bswap_i16
  component ahir_glue_bswap_i16 is -- 
    generic (tag_length : integer); 
    port ( -- 
      i : in  std_logic_vector(15 downto 0);
      ret_val_x_x : out  std_logic_vector(15 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_bswap_i16
  signal ahir_glue_bswap_i16_i :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_ret_val_x_x :  std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_in_args    : std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_out_args   : std_logic_vector(15 downto 0);
  signal ahir_glue_bswap_i16_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal ahir_glue_bswap_i16_tag_out   : std_logic_vector(2 downto 0);
  signal ahir_glue_bswap_i16_start_req : std_logic;
  signal ahir_glue_bswap_i16_start_ack : std_logic;
  signal ahir_glue_bswap_i16_fin_req   : std_logic;
  signal ahir_glue_bswap_i16_fin_ack : std_logic;
  -- caller side aggregated signals for module ahir_glue_bswap_i16
  signal ahir_glue_bswap_i16_call_reqs: std_logic_vector(6 downto 0);
  signal ahir_glue_bswap_i16_call_acks: std_logic_vector(6 downto 0);
  signal ahir_glue_bswap_i16_return_reqs: std_logic_vector(6 downto 0);
  signal ahir_glue_bswap_i16_return_acks: std_logic_vector(6 downto 0);
  signal ahir_glue_bswap_i16_call_data: std_logic_vector(111 downto 0);
  signal ahir_glue_bswap_i16_call_tag: std_logic_vector(13 downto 0);
  signal ahir_glue_bswap_i16_return_data: std_logic_vector(111 downto 0);
  signal ahir_glue_bswap_i16_return_tag: std_logic_vector(13 downto 0);
  -- declarations related to module ahir_glue_chk
  component ahir_glue_chk is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_chk
  signal ahir_glue_chk_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_chk_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_chk_start_req : std_logic;
  signal ahir_glue_chk_start_ack : std_logic;
  signal ahir_glue_chk_fin_req   : std_logic;
  signal ahir_glue_chk_fin_ack : std_logic;
  -- declarations related to module ahir_glue_chk_1
  component ahir_glue_chk_1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      chk_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      chk_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      chk_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      rtt_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      rtt_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_chk_1
  signal ahir_glue_chk_1_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_chk_1_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_chk_1_start_req : std_logic;
  signal ahir_glue_chk_1_start_ack : std_logic;
  signal ahir_glue_chk_1_fin_req   : std_logic;
  signal ahir_glue_chk_1_fin_ack : std_logic;
  -- declarations related to module ahir_glue_rtt
  component ahir_glue_rtt is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(8 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(4 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_3_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_lr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_3_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_3_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_lr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_4_lc_tag :  in  std_logic_vector(0 downto 0);
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_3_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sr_addr : out  std_logic_vector(13 downto 0);
      memory_space_3_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_3_sr_tag :  out  std_logic_vector(7 downto 0);
      memory_space_3_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_3_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_3_sc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_4_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sr_addr : out  std_logic_vector(0 downto 0);
      memory_space_4_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_4_sr_tag :  out  std_logic_vector(3 downto 0);
      memory_space_4_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_4_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_4_sc_tag :  in  std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      rtt_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      to0_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to0_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to0_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to1_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to1_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to1_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to2_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to2_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to2_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      to3_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      to3_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      to3_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_rtt
  signal ahir_glue_rtt_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_rtt_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_start_req : std_logic;
  signal ahir_glue_rtt_start_ack : std_logic;
  signal ahir_glue_rtt_fin_req   : std_logic;
  signal ahir_glue_rtt_fin_ack : std_logic;
  -- declarations related to module ahir_glue_src
  component ahir_glue_src is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      src_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      src_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      src_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      chk_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      chk_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      chk_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_src
  signal ahir_glue_src_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_src_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_src_start_req : std_logic;
  signal ahir_glue_src_start_ack : std_logic;
  signal ahir_glue_src_fin_req   : std_logic;
  signal ahir_glue_src_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to0
  component ahir_glue_to0 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to0_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to0_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to0_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga0_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to0
  signal ahir_glue_to0_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to0_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to0_start_req : std_logic;
  signal ahir_glue_to0_start_ack : std_logic;
  signal ahir_glue_to0_fin_req   : std_logic;
  signal ahir_glue_to0_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to1
  component ahir_glue_to1 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to1_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to1_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to1_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga1_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to1
  signal ahir_glue_to1_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to1_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to1_start_req : std_logic;
  signal ahir_glue_to1_start_ack : std_logic;
  signal ahir_glue_to1_fin_req   : std_logic;
  signal ahir_glue_to1_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to2
  component ahir_glue_to2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to2_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to2_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to2_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga2_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to2
  signal ahir_glue_to2_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to2_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to2_start_req : std_logic;
  signal ahir_glue_to2_start_ack : std_logic;
  signal ahir_glue_to2_fin_req   : std_logic;
  signal ahir_glue_to2_fin_ack : std_logic;
  -- declarations related to module ahir_glue_to3
  component ahir_glue_to3 is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      to3_in0_pipe_read_req : out  std_logic_vector(0 downto 0);
      to3_in0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      to3_in0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga3_out0_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_write_data : out  std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_write_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_write_data : out  std_logic_vector(31 downto 0);
      ahir_glue_bswap_i16_call_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_call_data : out  std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_call_tag  :  out  std_logic_vector(1 downto 0);
      ahir_glue_bswap_i16_return_reqs : out  std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_acks : in   std_logic_vector(0 downto 0);
      ahir_glue_bswap_i16_return_data : in   std_logic_vector(15 downto 0);
      ahir_glue_bswap_i16_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module ahir_glue_to3
  signal ahir_glue_to3_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal ahir_glue_to3_tag_out   : std_logic_vector(0 downto 0);
  signal ahir_glue_to3_start_req : std_logic;
  signal ahir_glue_to3_start_ack : std_logic;
  signal ahir_glue_to3_fin_req   : std_logic;
  signal ahir_glue_to3_fin_ack : std_logic;
  -- declarations related to module analyze_packet
  component analyze_packet is -- 
    generic (tag_length : integer); 
    port ( -- 
      pkt : in  std_logic_vector(31 downto 0);
      buf : out  std_logic_vector(31 downto 0);
      wlen : out  std_logic_vector(15 downto 0);
      blen : out  std_logic_vector(15 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module analyze_packet
  signal analyze_packet_pkt :  std_logic_vector(31 downto 0);
  signal analyze_packet_buf :  std_logic_vector(31 downto 0);
  signal analyze_packet_wlen :  std_logic_vector(15 downto 0);
  signal analyze_packet_blen :  std_logic_vector(15 downto 0);
  signal analyze_packet_in_args    : std_logic_vector(31 downto 0);
  signal analyze_packet_out_args   : std_logic_vector(63 downto 0);
  signal analyze_packet_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal analyze_packet_tag_out   : std_logic_vector(0 downto 0);
  signal analyze_packet_start_req : std_logic;
  signal analyze_packet_start_ack : std_logic;
  signal analyze_packet_fin_req   : std_logic;
  signal analyze_packet_fin_ack : std_logic;
  -- caller side aggregated signals for module analyze_packet
  signal analyze_packet_call_reqs: std_logic_vector(0 downto 0);
  signal analyze_packet_call_acks: std_logic_vector(0 downto 0);
  signal analyze_packet_return_reqs: std_logic_vector(0 downto 0);
  signal analyze_packet_return_acks: std_logic_vector(0 downto 0);
  signal analyze_packet_call_data: std_logic_vector(31 downto 0);
  signal analyze_packet_call_tag: std_logic_vector(0 downto 0);
  signal analyze_packet_return_data: std_logic_vector(63 downto 0);
  signal analyze_packet_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module click_bc_storage_initializer_x
  component click_bc_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      GV_15_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
      GV_15_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_reqs : out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_acks : in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_call_tag  :  out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_reqs : out  std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_acks : in   std_logic_vector(0 downto 0);
      GV_16_initializer_in_click_bc_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module click_bc_storage_initializer_x
  signal click_bc_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal click_bc_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_start_req : std_logic;
  signal click_bc_storage_initializer_x_start_ack : std_logic;
  signal click_bc_storage_initializer_x_fin_req   : std_logic;
  signal click_bc_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module click_bc_storage_initializer_x
  signal click_bc_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal click_bc_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module free_queue_init
  component free_queue_init is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module free_queue_init
  signal free_queue_init_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal free_queue_init_tag_out   : std_logic_vector(0 downto 0);
  signal free_queue_init_start_req : std_logic;
  signal free_queue_init_start_ack : std_logic;
  signal free_queue_init_fin_req   : std_logic;
  signal free_queue_init_fin_ack : std_logic;
  -- caller side aggregated signals for module free_queue_init
  signal free_queue_init_call_reqs: std_logic_vector(0 downto 0);
  signal free_queue_init_call_acks: std_logic_vector(0 downto 0);
  signal free_queue_init_return_reqs: std_logic_vector(0 downto 0);
  signal free_queue_init_return_acks: std_logic_vector(0 downto 0);
  signal free_queue_init_call_tag: std_logic_vector(0 downto 0);
  signal free_queue_init_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module global_storage_initializer_x
  component global_storage_initializer_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      click_bc_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      click_bc_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module global_storage_initializer_x
  signal global_storage_initializer_x_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal global_storage_initializer_x_tag_out   : std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_start_req : std_logic;
  signal global_storage_initializer_x_start_ack : std_logic;
  signal global_storage_initializer_x_fin_req   : std_logic;
  signal global_storage_initializer_x_fin_ack : std_logic;
  -- caller side aggregated signals for module global_storage_initializer_x
  signal global_storage_initializer_x_call_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_reqs: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_acks: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_call_tag: std_logic_vector(0 downto 0);
  signal global_storage_initializer_x_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module receive_packet_pipeline
  component receive_packet_pipeline is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_sr_data : out  std_logic_vector(7 downto 0);
      memory_space_5_sr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_sc_tag :  in  std_logic_vector(4 downto 0);
      free_queue_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      in_ctrl_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_ctrl_pipe_read_data : in   std_logic_vector(7 downto 0);
      in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      receive_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
      swapped_in_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      swapped_in_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      swapped_in_data_pipe_read_data : in   std_logic_vector(63 downto 0);
      receive_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
      receive_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
      swapped_in_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      swapped_in_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      swapped_in_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      receive_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module receive_packet_pipeline
  signal receive_packet_pipeline_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal receive_packet_pipeline_tag_out   : std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_start_req : std_logic;
  signal receive_packet_pipeline_start_ack : std_logic;
  signal receive_packet_pipeline_fin_req   : std_logic;
  signal receive_packet_pipeline_fin_ack : std_logic;
  -- declarations related to module send_packet_pipeline
  component send_packet_pipeline is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_5_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lr_addr : out  std_logic_vector(15 downto 0);
      memory_space_5_lr_tag :  out  std_logic_vector(10 downto 0);
      memory_space_5_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_5_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_5_lc_data : in   std_logic_vector(7 downto 0);
      memory_space_5_lc_tag :  in  std_logic_vector(4 downto 0);
      send_packet_buf_queue_pipe_read_req : out  std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_read_ack : in   std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_read_data : in   std_logic_vector(31 downto 0);
      send_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      free_queue_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      free_queue_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      out_ctrl_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_ctrl_pipe_write_data : out  std_logic_vector(7 downto 0);
      out_data_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_write_data : out  std_logic_vector(63 downto 0);
      send_packet_buf_queue_pipe_write_req : out  std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_write_ack : in   std_logic_vector(0 downto 0);
      send_packet_buf_queue_pipe_write_data : out  std_logic_vector(31 downto 0);
      analyze_packet_call_reqs : out  std_logic_vector(0 downto 0);
      analyze_packet_call_acks : in   std_logic_vector(0 downto 0);
      analyze_packet_call_data : out  std_logic_vector(31 downto 0);
      analyze_packet_call_tag  :  out  std_logic_vector(0 downto 0);
      analyze_packet_return_reqs : out  std_logic_vector(0 downto 0);
      analyze_packet_return_acks : in   std_logic_vector(0 downto 0);
      analyze_packet_return_data : in   std_logic_vector(63 downto 0);
      analyze_packet_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module send_packet_pipeline
  signal send_packet_pipeline_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal send_packet_pipeline_tag_out   : std_logic_vector(0 downto 0);
  signal send_packet_pipeline_start_req : std_logic;
  signal send_packet_pipeline_start_ack : std_logic;
  signal send_packet_pipeline_fin_req   : std_logic;
  signal send_packet_pipeline_fin_ack : std_logic;
  -- declarations related to module wrapper_input
  component wrapper_input is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      receive_packet_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      receive_packet_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      src_in0_pipe_write_req : out  std_logic_vector(0 downto 0);
      src_in0_pipe_write_ack : in   std_logic_vector(0 downto 0);
      src_in0_pipe_write_data : out  std_logic_vector(31 downto 0);
      global_storage_initializer_x_call_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_call_tag  :  out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_reqs : out  std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_acks : in   std_logic_vector(0 downto 0);
      global_storage_initializer_x_return_tag :  in   std_logic_vector(0 downto 0);
      free_queue_init_call_reqs : out  std_logic_vector(0 downto 0);
      free_queue_init_call_acks : in   std_logic_vector(0 downto 0);
      free_queue_init_call_tag  :  out  std_logic_vector(0 downto 0);
      free_queue_init_return_reqs : out  std_logic_vector(0 downto 0);
      free_queue_init_return_acks : in   std_logic_vector(0 downto 0);
      free_queue_init_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_input
  signal wrapper_input_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_input_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic;
  signal wrapper_input_start_ack : std_logic;
  signal wrapper_input_fin_req   : std_logic;
  signal wrapper_input_fin_ack : std_logic;
  -- declarations related to module wrapper_output
  component wrapper_output is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tofpga0_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga0_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga1_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga1_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga2_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga2_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga3_out0_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga3_out0_pipe_read_data : in   std_logic_vector(31 downto 0);
      tofpga_port_number_pipe_read_req : out  std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_read_ack : in   std_logic_vector(0 downto 0);
      tofpga_port_number_pipe_read_data : in   std_logic_vector(31 downto 0);
      send_packet_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      send_packet_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module wrapper_output
  signal wrapper_output_tag_in    : std_logic_vector(0 downto 0) := (others => '0');
  signal wrapper_output_tag_out   : std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic;
  signal wrapper_output_start_ack : std_logic;
  signal wrapper_output_fin_req   : std_logic;
  signal wrapper_output_fin_ack : std_logic;
  -- aggregate signals for write to pipe chk_in0
  signal chk_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal chk_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal chk_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe chk_in0
  signal chk_in0_pipe_read_data: std_logic_vector(63 downto 0);
  signal chk_in0_pipe_read_req: std_logic_vector(1 downto 0);
  signal chk_in0_pipe_read_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for write to pipe free_queue_pipe
  signal free_queue_pipe_pipe_write_data: std_logic_vector(159 downto 0);
  signal free_queue_pipe_pipe_write_req: std_logic_vector(4 downto 0);
  signal free_queue_pipe_pipe_write_ack: std_logic_vector(4 downto 0);
  -- aggregate signals for read from pipe free_queue_pipe
  signal free_queue_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal free_queue_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal free_queue_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_ctrl
  signal in_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_ctrl_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data
  signal in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_ctrl
  signal out_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_ctrl_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data
  signal out_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe receive_packet_buf_queue
  signal receive_packet_buf_queue_pipe_write_data: std_logic_vector(31 downto 0);
  signal receive_packet_buf_queue_pipe_write_req: std_logic_vector(0 downto 0);
  signal receive_packet_buf_queue_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe receive_packet_buf_queue
  signal receive_packet_buf_queue_pipe_read_data: std_logic_vector(31 downto 0);
  signal receive_packet_buf_queue_pipe_read_req: std_logic_vector(0 downto 0);
  signal receive_packet_buf_queue_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe receive_packet_pipe
  signal receive_packet_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal receive_packet_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal receive_packet_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe receive_packet_pipe
  signal receive_packet_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal receive_packet_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal receive_packet_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe rtt_in0
  signal rtt_in0_pipe_write_data: std_logic_vector(63 downto 0);
  signal rtt_in0_pipe_write_req: std_logic_vector(1 downto 0);
  signal rtt_in0_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe rtt_in0
  signal rtt_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal rtt_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal rtt_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe send_packet_buf_queue
  signal send_packet_buf_queue_pipe_write_data: std_logic_vector(31 downto 0);
  signal send_packet_buf_queue_pipe_write_req: std_logic_vector(0 downto 0);
  signal send_packet_buf_queue_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe send_packet_buf_queue
  signal send_packet_buf_queue_pipe_read_data: std_logic_vector(31 downto 0);
  signal send_packet_buf_queue_pipe_read_req: std_logic_vector(0 downto 0);
  signal send_packet_buf_queue_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe send_packet_pipe
  signal send_packet_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal send_packet_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal send_packet_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe send_packet_pipe
  signal send_packet_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal send_packet_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal send_packet_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe src_in0
  signal src_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal src_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal src_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe src_in0
  signal src_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal src_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal src_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe swapped_in_data
  signal swapped_in_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal swapped_in_data_pipe_write_req: std_logic_vector(0 downto 0);
  signal swapped_in_data_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe swapped_in_data
  signal swapped_in_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal swapped_in_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal swapped_in_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to0_in0
  signal to0_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to0_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to0_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to0_in0
  signal to0_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to0_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to0_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to1_in0
  signal to1_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to1_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to1_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to1_in0
  signal to1_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to1_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to1_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to2_in0
  signal to2_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to2_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to2_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to2_in0
  signal to2_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to2_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to2_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe to3_in0
  signal to3_in0_pipe_write_data: std_logic_vector(31 downto 0);
  signal to3_in0_pipe_write_req: std_logic_vector(0 downto 0);
  signal to3_in0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe to3_in0
  signal to3_in0_pipe_read_data: std_logic_vector(31 downto 0);
  signal to3_in0_pipe_read_req: std_logic_vector(0 downto 0);
  signal to3_in0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga0_out0
  signal tofpga0_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga0_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga0_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga0_out0
  signal tofpga0_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga0_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga0_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga1_out0
  signal tofpga1_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga1_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga1_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga1_out0
  signal tofpga1_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga1_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga1_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga2_out0
  signal tofpga2_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga2_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga2_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga2_out0
  signal tofpga2_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga2_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga2_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga3_out0
  signal tofpga3_out0_pipe_write_data: std_logic_vector(31 downto 0);
  signal tofpga3_out0_pipe_write_req: std_logic_vector(0 downto 0);
  signal tofpga3_out0_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe tofpga3_out0
  signal tofpga3_out0_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga3_out0_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga3_out0_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe tofpga_port_number
  signal tofpga_port_number_pipe_write_data: std_logic_vector(127 downto 0);
  signal tofpga_port_number_pipe_write_req: std_logic_vector(3 downto 0);
  signal tofpga_port_number_pipe_write_ack: std_logic_vector(3 downto 0);
  -- aggregate signals for read from pipe tofpga_port_number
  signal tofpga_port_number_pipe_read_data: std_logic_vector(31 downto 0);
  signal tofpga_port_number_pipe_read_req: std_logic_vector(0 downto 0);
  signal tofpga_port_number_pipe_read_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module GV_15_initializer_in_click_bc
  -- call arbiter for module GV_15_initializer_in_click_bc
  GV_15_initializer_in_click_bc_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => GV_15_initializer_in_click_bc_call_reqs,
      call_acks => GV_15_initializer_in_click_bc_call_acks,
      return_reqs => GV_15_initializer_in_click_bc_return_reqs,
      return_acks => GV_15_initializer_in_click_bc_return_acks,
      call_tag  => GV_15_initializer_in_click_bc_call_tag,
      return_tag  => GV_15_initializer_in_click_bc_return_tag,
      call_mtag => GV_15_initializer_in_click_bc_tag_in,
      return_mtag => GV_15_initializer_in_click_bc_tag_out,
      call_mreq => GV_15_initializer_in_click_bc_start_req,
      call_mack => GV_15_initializer_in_click_bc_start_ack,
      return_mreq => GV_15_initializer_in_click_bc_fin_req,
      return_mack => GV_15_initializer_in_click_bc_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  GV_15_initializer_in_click_bc_instance:GV_15_initializer_in_click_bc-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => GV_15_initializer_in_click_bc_start_req,
      start_ack => GV_15_initializer_in_click_bc_start_ack,
      fin_req => GV_15_initializer_in_click_bc_fin_req,
      fin_ack => GV_15_initializer_in_click_bc_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(8 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(7 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(7 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(4 downto 0),
      tag_in => GV_15_initializer_in_click_bc_tag_in,
      tag_out => GV_15_initializer_in_click_bc_tag_out-- 
    ); -- 
  -- module GV_16_initializer_in_click_bc
  -- call arbiter for module GV_16_initializer_in_click_bc
  GV_16_initializer_in_click_bc_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => GV_16_initializer_in_click_bc_call_reqs,
      call_acks => GV_16_initializer_in_click_bc_call_acks,
      return_reqs => GV_16_initializer_in_click_bc_return_reqs,
      return_acks => GV_16_initializer_in_click_bc_return_acks,
      call_tag  => GV_16_initializer_in_click_bc_call_tag,
      return_tag  => GV_16_initializer_in_click_bc_return_tag,
      call_mtag => GV_16_initializer_in_click_bc_tag_in,
      return_mtag => GV_16_initializer_in_click_bc_tag_out,
      call_mreq => GV_16_initializer_in_click_bc_start_req,
      call_mack => GV_16_initializer_in_click_bc_start_ack,
      return_mreq => GV_16_initializer_in_click_bc_fin_req,
      return_mack => GV_16_initializer_in_click_bc_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  GV_16_initializer_in_click_bc_instance:GV_16_initializer_in_click_bc-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => GV_16_initializer_in_click_bc_start_req,
      start_ack => GV_16_initializer_in_click_bc_start_ack,
      fin_req => GV_16_initializer_in_click_bc_fin_req,
      fin_ack => GV_16_initializer_in_click_bc_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(4 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(6 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      tag_in => GV_16_initializer_in_click_bc_tag_in,
      tag_out => GV_16_initializer_in_click_bc_tag_out-- 
    ); -- 
  -- module ahir_glue_bswap_i16
  ahir_glue_bswap_i16_i <= ahir_glue_bswap_i16_in_args(15 downto 0);
  ahir_glue_bswap_i16_out_args <= ahir_glue_bswap_i16_ret_val_x_x ;
  -- call arbiter for module ahir_glue_bswap_i16
  ahir_glue_bswap_i16_arbiter: SplitCallArbiter -- 
    generic map( --
      num_reqs => 7,
      call_data_width => 16,
      return_data_width => 16,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => ahir_glue_bswap_i16_call_reqs,
      call_acks => ahir_glue_bswap_i16_call_acks,
      return_reqs => ahir_glue_bswap_i16_return_reqs,
      return_acks => ahir_glue_bswap_i16_return_acks,
      call_data  => ahir_glue_bswap_i16_call_data,
      call_tag  => ahir_glue_bswap_i16_call_tag,
      return_tag  => ahir_glue_bswap_i16_return_tag,
      call_mtag => ahir_glue_bswap_i16_tag_in,
      return_mtag => ahir_glue_bswap_i16_tag_out,
      return_data =>ahir_glue_bswap_i16_return_data,
      call_mreq => ahir_glue_bswap_i16_start_req,
      call_mack => ahir_glue_bswap_i16_start_ack,
      return_mreq => ahir_glue_bswap_i16_fin_req,
      return_mack => ahir_glue_bswap_i16_fin_ack,
      call_mdata => ahir_glue_bswap_i16_in_args,
      return_mdata => ahir_glue_bswap_i16_out_args,
      clk => clk, 
      reset => reset --
    ); --
  ahir_glue_bswap_i16_instance:ahir_glue_bswap_i16-- 
    generic map(tag_length => 3)
    port map(-- 
      i => ahir_glue_bswap_i16_i,
      ret_val_x_x => ahir_glue_bswap_i16_ret_val_x_x,
      start_req => ahir_glue_bswap_i16_start_req,
      start_ack => ahir_glue_bswap_i16_start_ack,
      fin_req => ahir_glue_bswap_i16_fin_req,
      fin_ack => ahir_glue_bswap_i16_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => ahir_glue_bswap_i16_tag_in,
      tag_out => ahir_glue_bswap_i16_tag_out-- 
    ); -- 
  -- module ahir_glue_chk
  ahir_glue_chk_instance:ahir_glue_chk-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_chk_start_req,
      start_ack => ahir_glue_chk_start_ack,
      fin_req => ahir_glue_chk_fin_req,
      fin_ack => ahir_glue_chk_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(9 downto 9),
      memory_space_5_lr_ack => memory_space_5_lr_ack(9 downto 9),
      memory_space_5_lr_addr => memory_space_5_lr_addr(159 downto 144),
      memory_space_5_lr_tag => memory_space_5_lr_tag(109 downto 99),
      memory_space_5_lc_req => memory_space_5_lc_req(9 downto 9),
      memory_space_5_lc_ack => memory_space_5_lc_ack(9 downto 9),
      memory_space_5_lc_data => memory_space_5_lc_data(79 downto 72),
      memory_space_5_lc_tag => memory_space_5_lc_tag(49 downto 45),
      memory_space_5_sr_req => memory_space_5_sr_req(7 downto 7),
      memory_space_5_sr_ack => memory_space_5_sr_ack(7 downto 7),
      memory_space_5_sr_addr => memory_space_5_sr_addr(127 downto 112),
      memory_space_5_sr_data => memory_space_5_sr_data(63 downto 56),
      memory_space_5_sr_tag => memory_space_5_sr_tag(87 downto 77),
      memory_space_5_sc_req => memory_space_5_sc_req(7 downto 7),
      memory_space_5_sc_ack => memory_space_5_sc_ack(7 downto 7),
      memory_space_5_sc_tag => memory_space_5_sc_tag(39 downto 35),
      chk_in0_pipe_read_req => chk_in0_pipe_read_req(1 downto 1),
      chk_in0_pipe_read_ack => chk_in0_pipe_read_ack(1 downto 1),
      chk_in0_pipe_read_data => chk_in0_pipe_read_data(63 downto 32),
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(4 downto 4),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(4 downto 4),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(159 downto 128),
      rtt_in0_pipe_write_req => rtt_in0_pipe_write_req(1 downto 1),
      rtt_in0_pipe_write_ack => rtt_in0_pipe_write_ack(1 downto 1),
      rtt_in0_pipe_write_data => rtt_in0_pipe_write_data(63 downto 32),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(6 downto 6),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(6 downto 6),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(111 downto 96),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(13 downto 12),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(6 downto 6),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(6 downto 6),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(111 downto 96),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(13 downto 12),
      tag_in => ahir_glue_chk_tag_in,
      tag_out => ahir_glue_chk_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_chk_tag_in <= (others => '0');
  ahir_glue_chk_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_chk_start_req, start_ack => ahir_glue_chk_start_ack,  fin_req => ahir_glue_chk_fin_req,  fin_ack => ahir_glue_chk_fin_ack);
  -- module ahir_glue_chk_1
  ahir_glue_chk_1_instance:ahir_glue_chk_1-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_chk_1_start_req,
      start_ack => ahir_glue_chk_1_start_ack,
      fin_req => ahir_glue_chk_1_fin_req,
      fin_ack => ahir_glue_chk_1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(8 downto 8),
      memory_space_5_lr_ack => memory_space_5_lr_ack(8 downto 8),
      memory_space_5_lr_addr => memory_space_5_lr_addr(143 downto 128),
      memory_space_5_lr_tag => memory_space_5_lr_tag(98 downto 88),
      memory_space_5_lc_req => memory_space_5_lc_req(8 downto 8),
      memory_space_5_lc_ack => memory_space_5_lc_ack(8 downto 8),
      memory_space_5_lc_data => memory_space_5_lc_data(71 downto 64),
      memory_space_5_lc_tag => memory_space_5_lc_tag(44 downto 40),
      memory_space_5_sr_req => memory_space_5_sr_req(6 downto 6),
      memory_space_5_sr_ack => memory_space_5_sr_ack(6 downto 6),
      memory_space_5_sr_addr => memory_space_5_sr_addr(111 downto 96),
      memory_space_5_sr_data => memory_space_5_sr_data(55 downto 48),
      memory_space_5_sr_tag => memory_space_5_sr_tag(76 downto 66),
      memory_space_5_sc_req => memory_space_5_sc_req(6 downto 6),
      memory_space_5_sc_ack => memory_space_5_sc_ack(6 downto 6),
      memory_space_5_sc_tag => memory_space_5_sc_tag(34 downto 30),
      chk_in0_pipe_read_req => chk_in0_pipe_read_req(0 downto 0),
      chk_in0_pipe_read_ack => chk_in0_pipe_read_ack(0 downto 0),
      chk_in0_pipe_read_data => chk_in0_pipe_read_data(31 downto 0),
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(3 downto 3),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(3 downto 3),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(127 downto 96),
      rtt_in0_pipe_write_req => rtt_in0_pipe_write_req(0 downto 0),
      rtt_in0_pipe_write_ack => rtt_in0_pipe_write_ack(0 downto 0),
      rtt_in0_pipe_write_data => rtt_in0_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(5 downto 5),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(5 downto 5),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(95 downto 80),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(11 downto 10),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(5 downto 5),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(5 downto 5),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(95 downto 80),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(11 downto 10),
      tag_in => ahir_glue_chk_1_tag_in,
      tag_out => ahir_glue_chk_1_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_chk_1_tag_in <= (others => '0');
  ahir_glue_chk_1_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_chk_1_start_req, start_ack => ahir_glue_chk_1_start_ack,  fin_req => ahir_glue_chk_1_fin_req,  fin_ack => ahir_glue_chk_1_fin_ack);
  -- module ahir_glue_rtt
  ahir_glue_rtt_instance:ahir_glue_rtt-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_rtt_start_req,
      start_ack => ahir_glue_rtt_start_ack,
      fin_req => ahir_glue_rtt_fin_req,
      fin_ack => ahir_glue_rtt_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(8 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(7 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(7 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(4 downto 0),
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(4 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(6 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      memory_space_3_lr_req => memory_space_3_lr_req(0 downto 0),
      memory_space_3_lr_ack => memory_space_3_lr_ack(0 downto 0),
      memory_space_3_lr_addr => memory_space_3_lr_addr(13 downto 0),
      memory_space_3_lr_tag => memory_space_3_lr_tag(7 downto 0),
      memory_space_3_lc_req => memory_space_3_lc_req(0 downto 0),
      memory_space_3_lc_ack => memory_space_3_lc_ack(0 downto 0),
      memory_space_3_lc_data => memory_space_3_lc_data(7 downto 0),
      memory_space_3_lc_tag => memory_space_3_lc_tag(4 downto 0),
      memory_space_4_lr_req => memory_space_4_lr_req(0 downto 0),
      memory_space_4_lr_ack => memory_space_4_lr_ack(0 downto 0),
      memory_space_4_lr_addr => memory_space_4_lr_addr(0 downto 0),
      memory_space_4_lr_tag => memory_space_4_lr_tag(3 downto 0),
      memory_space_4_lc_req => memory_space_4_lc_req(0 downto 0),
      memory_space_4_lc_ack => memory_space_4_lc_ack(0 downto 0),
      memory_space_4_lc_data => memory_space_4_lc_data(31 downto 0),
      memory_space_4_lc_tag => memory_space_4_lc_tag(0 downto 0),
      memory_space_5_lr_req => memory_space_5_lr_req(7 downto 7),
      memory_space_5_lr_ack => memory_space_5_lr_ack(7 downto 7),
      memory_space_5_lr_addr => memory_space_5_lr_addr(127 downto 112),
      memory_space_5_lr_tag => memory_space_5_lr_tag(87 downto 77),
      memory_space_5_lc_req => memory_space_5_lc_req(7 downto 7),
      memory_space_5_lc_ack => memory_space_5_lc_ack(7 downto 7),
      memory_space_5_lc_data => memory_space_5_lc_data(63 downto 56),
      memory_space_5_lc_tag => memory_space_5_lc_tag(39 downto 35),
      memory_space_3_sr_req => memory_space_3_sr_req(0 downto 0),
      memory_space_3_sr_ack => memory_space_3_sr_ack(0 downto 0),
      memory_space_3_sr_addr => memory_space_3_sr_addr(13 downto 0),
      memory_space_3_sr_data => memory_space_3_sr_data(7 downto 0),
      memory_space_3_sr_tag => memory_space_3_sr_tag(7 downto 0),
      memory_space_3_sc_req => memory_space_3_sc_req(0 downto 0),
      memory_space_3_sc_ack => memory_space_3_sc_ack(0 downto 0),
      memory_space_3_sc_tag => memory_space_3_sc_tag(4 downto 0),
      memory_space_4_sr_req => memory_space_4_sr_req(0 downto 0),
      memory_space_4_sr_ack => memory_space_4_sr_ack(0 downto 0),
      memory_space_4_sr_addr => memory_space_4_sr_addr(0 downto 0),
      memory_space_4_sr_data => memory_space_4_sr_data(31 downto 0),
      memory_space_4_sr_tag => memory_space_4_sr_tag(3 downto 0),
      memory_space_4_sc_req => memory_space_4_sc_req(0 downto 0),
      memory_space_4_sc_ack => memory_space_4_sc_ack(0 downto 0),
      memory_space_4_sc_tag => memory_space_4_sc_tag(0 downto 0),
      rtt_in0_pipe_read_req => rtt_in0_pipe_read_req(0 downto 0),
      rtt_in0_pipe_read_ack => rtt_in0_pipe_read_ack(0 downto 0),
      rtt_in0_pipe_read_data => rtt_in0_pipe_read_data(31 downto 0),
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(2 downto 2),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(2 downto 2),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(95 downto 64),
      to0_in0_pipe_write_req => to0_in0_pipe_write_req(0 downto 0),
      to0_in0_pipe_write_ack => to0_in0_pipe_write_ack(0 downto 0),
      to0_in0_pipe_write_data => to0_in0_pipe_write_data(31 downto 0),
      to1_in0_pipe_write_req => to1_in0_pipe_write_req(0 downto 0),
      to1_in0_pipe_write_ack => to1_in0_pipe_write_ack(0 downto 0),
      to1_in0_pipe_write_data => to1_in0_pipe_write_data(31 downto 0),
      to2_in0_pipe_write_req => to2_in0_pipe_write_req(0 downto 0),
      to2_in0_pipe_write_ack => to2_in0_pipe_write_ack(0 downto 0),
      to2_in0_pipe_write_data => to2_in0_pipe_write_data(31 downto 0),
      to3_in0_pipe_write_req => to3_in0_pipe_write_req(0 downto 0),
      to3_in0_pipe_write_ack => to3_in0_pipe_write_ack(0 downto 0),
      to3_in0_pipe_write_data => to3_in0_pipe_write_data(31 downto 0),
      tag_in => ahir_glue_rtt_tag_in,
      tag_out => ahir_glue_rtt_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_rtt_tag_in <= (others => '0');
  ahir_glue_rtt_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_rtt_start_req, start_ack => ahir_glue_rtt_start_ack,  fin_req => ahir_glue_rtt_fin_req,  fin_ack => ahir_glue_rtt_fin_ack);
  -- module ahir_glue_src
  ahir_glue_src_instance:ahir_glue_src-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_src_start_req,
      start_ack => ahir_glue_src_start_ack,
      fin_req => ahir_glue_src_fin_req,
      fin_ack => ahir_glue_src_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(6 downto 6),
      memory_space_5_lr_ack => memory_space_5_lr_ack(6 downto 6),
      memory_space_5_lr_addr => memory_space_5_lr_addr(111 downto 96),
      memory_space_5_lr_tag => memory_space_5_lr_tag(76 downto 66),
      memory_space_5_lc_req => memory_space_5_lc_req(6 downto 6),
      memory_space_5_lc_ack => memory_space_5_lc_ack(6 downto 6),
      memory_space_5_lc_data => memory_space_5_lc_data(55 downto 48),
      memory_space_5_lc_tag => memory_space_5_lc_tag(34 downto 30),
      memory_space_5_sr_req => memory_space_5_sr_req(5 downto 5),
      memory_space_5_sr_ack => memory_space_5_sr_ack(5 downto 5),
      memory_space_5_sr_addr => memory_space_5_sr_addr(95 downto 80),
      memory_space_5_sr_data => memory_space_5_sr_data(47 downto 40),
      memory_space_5_sr_tag => memory_space_5_sr_tag(65 downto 55),
      memory_space_5_sc_req => memory_space_5_sc_req(5 downto 5),
      memory_space_5_sc_ack => memory_space_5_sc_ack(5 downto 5),
      memory_space_5_sc_tag => memory_space_5_sc_tag(29 downto 25),
      src_in0_pipe_read_req => src_in0_pipe_read_req(0 downto 0),
      src_in0_pipe_read_ack => src_in0_pipe_read_ack(0 downto 0),
      src_in0_pipe_read_data => src_in0_pipe_read_data(31 downto 0),
      chk_in0_pipe_write_req => chk_in0_pipe_write_req(0 downto 0),
      chk_in0_pipe_write_ack => chk_in0_pipe_write_ack(0 downto 0),
      chk_in0_pipe_write_data => chk_in0_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(4 downto 4),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(4 downto 4),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(79 downto 64),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(9 downto 8),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(4 downto 4),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(4 downto 4),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(79 downto 64),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(9 downto 8),
      tag_in => ahir_glue_src_tag_in,
      tag_out => ahir_glue_src_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_src_tag_in <= (others => '0');
  ahir_glue_src_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_src_start_req, start_ack => ahir_glue_src_start_ack,  fin_req => ahir_glue_src_fin_req,  fin_ack => ahir_glue_src_fin_ack);
  -- module ahir_glue_to0
  ahir_glue_to0_instance:ahir_glue_to0-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to0_start_req,
      start_ack => ahir_glue_to0_start_ack,
      fin_req => ahir_glue_to0_fin_req,
      fin_ack => ahir_glue_to0_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(5 downto 5),
      memory_space_5_lr_ack => memory_space_5_lr_ack(5 downto 5),
      memory_space_5_lr_addr => memory_space_5_lr_addr(95 downto 80),
      memory_space_5_lr_tag => memory_space_5_lr_tag(65 downto 55),
      memory_space_5_lc_req => memory_space_5_lc_req(5 downto 5),
      memory_space_5_lc_ack => memory_space_5_lc_ack(5 downto 5),
      memory_space_5_lc_data => memory_space_5_lc_data(47 downto 40),
      memory_space_5_lc_tag => memory_space_5_lc_tag(29 downto 25),
      memory_space_5_sr_req => memory_space_5_sr_req(4 downto 4),
      memory_space_5_sr_ack => memory_space_5_sr_ack(4 downto 4),
      memory_space_5_sr_addr => memory_space_5_sr_addr(79 downto 64),
      memory_space_5_sr_data => memory_space_5_sr_data(39 downto 32),
      memory_space_5_sr_tag => memory_space_5_sr_tag(54 downto 44),
      memory_space_5_sc_req => memory_space_5_sc_req(4 downto 4),
      memory_space_5_sc_ack => memory_space_5_sc_ack(4 downto 4),
      memory_space_5_sc_tag => memory_space_5_sc_tag(24 downto 20),
      to0_in0_pipe_read_req => to0_in0_pipe_read_req(0 downto 0),
      to0_in0_pipe_read_ack => to0_in0_pipe_read_ack(0 downto 0),
      to0_in0_pipe_read_data => to0_in0_pipe_read_data(31 downto 0),
      tofpga0_out0_pipe_write_req => tofpga0_out0_pipe_write_req(0 downto 0),
      tofpga0_out0_pipe_write_ack => tofpga0_out0_pipe_write_ack(0 downto 0),
      tofpga0_out0_pipe_write_data => tofpga0_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(3 downto 3),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(3 downto 3),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(127 downto 96),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(3 downto 3),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(3 downto 3),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(63 downto 48),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(7 downto 6),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(3 downto 3),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(3 downto 3),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(63 downto 48),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(7 downto 6),
      tag_in => ahir_glue_to0_tag_in,
      tag_out => ahir_glue_to0_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to0_tag_in <= (others => '0');
  ahir_glue_to0_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to0_start_req, start_ack => ahir_glue_to0_start_ack,  fin_req => ahir_glue_to0_fin_req,  fin_ack => ahir_glue_to0_fin_ack);
  -- module ahir_glue_to1
  ahir_glue_to1_instance:ahir_glue_to1-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to1_start_req,
      start_ack => ahir_glue_to1_start_ack,
      fin_req => ahir_glue_to1_fin_req,
      fin_ack => ahir_glue_to1_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(4 downto 4),
      memory_space_5_lr_ack => memory_space_5_lr_ack(4 downto 4),
      memory_space_5_lr_addr => memory_space_5_lr_addr(79 downto 64),
      memory_space_5_lr_tag => memory_space_5_lr_tag(54 downto 44),
      memory_space_5_lc_req => memory_space_5_lc_req(4 downto 4),
      memory_space_5_lc_ack => memory_space_5_lc_ack(4 downto 4),
      memory_space_5_lc_data => memory_space_5_lc_data(39 downto 32),
      memory_space_5_lc_tag => memory_space_5_lc_tag(24 downto 20),
      memory_space_5_sr_req => memory_space_5_sr_req(3 downto 3),
      memory_space_5_sr_ack => memory_space_5_sr_ack(3 downto 3),
      memory_space_5_sr_addr => memory_space_5_sr_addr(63 downto 48),
      memory_space_5_sr_data => memory_space_5_sr_data(31 downto 24),
      memory_space_5_sr_tag => memory_space_5_sr_tag(43 downto 33),
      memory_space_5_sc_req => memory_space_5_sc_req(3 downto 3),
      memory_space_5_sc_ack => memory_space_5_sc_ack(3 downto 3),
      memory_space_5_sc_tag => memory_space_5_sc_tag(19 downto 15),
      to1_in0_pipe_read_req => to1_in0_pipe_read_req(0 downto 0),
      to1_in0_pipe_read_ack => to1_in0_pipe_read_ack(0 downto 0),
      to1_in0_pipe_read_data => to1_in0_pipe_read_data(31 downto 0),
      tofpga1_out0_pipe_write_req => tofpga1_out0_pipe_write_req(0 downto 0),
      tofpga1_out0_pipe_write_ack => tofpga1_out0_pipe_write_ack(0 downto 0),
      tofpga1_out0_pipe_write_data => tofpga1_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(2 downto 2),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(2 downto 2),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(95 downto 64),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(2 downto 2),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(2 downto 2),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(47 downto 32),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(5 downto 4),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(2 downto 2),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(2 downto 2),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(47 downto 32),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(5 downto 4),
      tag_in => ahir_glue_to1_tag_in,
      tag_out => ahir_glue_to1_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to1_tag_in <= (others => '0');
  ahir_glue_to1_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to1_start_req, start_ack => ahir_glue_to1_start_ack,  fin_req => ahir_glue_to1_fin_req,  fin_ack => ahir_glue_to1_fin_ack);
  -- module ahir_glue_to2
  ahir_glue_to2_instance:ahir_glue_to2-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to2_start_req,
      start_ack => ahir_glue_to2_start_ack,
      fin_req => ahir_glue_to2_fin_req,
      fin_ack => ahir_glue_to2_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(3 downto 3),
      memory_space_5_lr_ack => memory_space_5_lr_ack(3 downto 3),
      memory_space_5_lr_addr => memory_space_5_lr_addr(63 downto 48),
      memory_space_5_lr_tag => memory_space_5_lr_tag(43 downto 33),
      memory_space_5_lc_req => memory_space_5_lc_req(3 downto 3),
      memory_space_5_lc_ack => memory_space_5_lc_ack(3 downto 3),
      memory_space_5_lc_data => memory_space_5_lc_data(31 downto 24),
      memory_space_5_lc_tag => memory_space_5_lc_tag(19 downto 15),
      memory_space_5_sr_req => memory_space_5_sr_req(2 downto 2),
      memory_space_5_sr_ack => memory_space_5_sr_ack(2 downto 2),
      memory_space_5_sr_addr => memory_space_5_sr_addr(47 downto 32),
      memory_space_5_sr_data => memory_space_5_sr_data(23 downto 16),
      memory_space_5_sr_tag => memory_space_5_sr_tag(32 downto 22),
      memory_space_5_sc_req => memory_space_5_sc_req(2 downto 2),
      memory_space_5_sc_ack => memory_space_5_sc_ack(2 downto 2),
      memory_space_5_sc_tag => memory_space_5_sc_tag(14 downto 10),
      to2_in0_pipe_read_req => to2_in0_pipe_read_req(0 downto 0),
      to2_in0_pipe_read_ack => to2_in0_pipe_read_ack(0 downto 0),
      to2_in0_pipe_read_data => to2_in0_pipe_read_data(31 downto 0),
      tofpga2_out0_pipe_write_req => tofpga2_out0_pipe_write_req(0 downto 0),
      tofpga2_out0_pipe_write_ack => tofpga2_out0_pipe_write_ack(0 downto 0),
      tofpga2_out0_pipe_write_data => tofpga2_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(1 downto 1),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(1 downto 1),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(63 downto 32),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(1 downto 1),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(1 downto 1),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(31 downto 16),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(3 downto 2),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(1 downto 1),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(1 downto 1),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(31 downto 16),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(3 downto 2),
      tag_in => ahir_glue_to2_tag_in,
      tag_out => ahir_glue_to2_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to2_tag_in <= (others => '0');
  ahir_glue_to2_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to2_start_req, start_ack => ahir_glue_to2_start_ack,  fin_req => ahir_glue_to2_fin_req,  fin_ack => ahir_glue_to2_fin_ack);
  -- module ahir_glue_to3
  ahir_glue_to3_instance:ahir_glue_to3-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => ahir_glue_to3_start_req,
      start_ack => ahir_glue_to3_start_ack,
      fin_req => ahir_glue_to3_fin_req,
      fin_ack => ahir_glue_to3_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(2 downto 2),
      memory_space_5_lr_ack => memory_space_5_lr_ack(2 downto 2),
      memory_space_5_lr_addr => memory_space_5_lr_addr(47 downto 32),
      memory_space_5_lr_tag => memory_space_5_lr_tag(32 downto 22),
      memory_space_5_lc_req => memory_space_5_lc_req(2 downto 2),
      memory_space_5_lc_ack => memory_space_5_lc_ack(2 downto 2),
      memory_space_5_lc_data => memory_space_5_lc_data(23 downto 16),
      memory_space_5_lc_tag => memory_space_5_lc_tag(14 downto 10),
      memory_space_5_sr_req => memory_space_5_sr_req(1 downto 1),
      memory_space_5_sr_ack => memory_space_5_sr_ack(1 downto 1),
      memory_space_5_sr_addr => memory_space_5_sr_addr(31 downto 16),
      memory_space_5_sr_data => memory_space_5_sr_data(15 downto 8),
      memory_space_5_sr_tag => memory_space_5_sr_tag(21 downto 11),
      memory_space_5_sc_req => memory_space_5_sc_req(1 downto 1),
      memory_space_5_sc_ack => memory_space_5_sc_ack(1 downto 1),
      memory_space_5_sc_tag => memory_space_5_sc_tag(9 downto 5),
      to3_in0_pipe_read_req => to3_in0_pipe_read_req(0 downto 0),
      to3_in0_pipe_read_ack => to3_in0_pipe_read_ack(0 downto 0),
      to3_in0_pipe_read_data => to3_in0_pipe_read_data(31 downto 0),
      tofpga3_out0_pipe_write_req => tofpga3_out0_pipe_write_req(0 downto 0),
      tofpga3_out0_pipe_write_ack => tofpga3_out0_pipe_write_ack(0 downto 0),
      tofpga3_out0_pipe_write_data => tofpga3_out0_pipe_write_data(31 downto 0),
      tofpga_port_number_pipe_write_req => tofpga_port_number_pipe_write_req(0 downto 0),
      tofpga_port_number_pipe_write_ack => tofpga_port_number_pipe_write_ack(0 downto 0),
      tofpga_port_number_pipe_write_data => tofpga_port_number_pipe_write_data(31 downto 0),
      ahir_glue_bswap_i16_call_reqs => ahir_glue_bswap_i16_call_reqs(0 downto 0),
      ahir_glue_bswap_i16_call_acks => ahir_glue_bswap_i16_call_acks(0 downto 0),
      ahir_glue_bswap_i16_call_data => ahir_glue_bswap_i16_call_data(15 downto 0),
      ahir_glue_bswap_i16_call_tag => ahir_glue_bswap_i16_call_tag(1 downto 0),
      ahir_glue_bswap_i16_return_reqs => ahir_glue_bswap_i16_return_reqs(0 downto 0),
      ahir_glue_bswap_i16_return_acks => ahir_glue_bswap_i16_return_acks(0 downto 0),
      ahir_glue_bswap_i16_return_data => ahir_glue_bswap_i16_return_data(15 downto 0),
      ahir_glue_bswap_i16_return_tag => ahir_glue_bswap_i16_return_tag(1 downto 0),
      tag_in => ahir_glue_to3_tag_in,
      tag_out => ahir_glue_to3_tag_out-- 
    ); -- 
  -- module will be run forever 
  ahir_glue_to3_tag_in <= (others => '0');
  ahir_glue_to3_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ahir_glue_to3_start_req, start_ack => ahir_glue_to3_start_ack,  fin_req => ahir_glue_to3_fin_req,  fin_ack => ahir_glue_to3_fin_ack);
  -- module analyze_packet
  analyze_packet_pkt <= analyze_packet_in_args(31 downto 0);
  analyze_packet_out_args <= analyze_packet_buf & analyze_packet_wlen & analyze_packet_blen ;
  -- call arbiter for module analyze_packet
  analyze_packet_arbiter: SplitCallArbiter -- 
    generic map( --
      num_reqs => 1,
      call_data_width => 32,
      return_data_width => 64,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => analyze_packet_call_reqs,
      call_acks => analyze_packet_call_acks,
      return_reqs => analyze_packet_return_reqs,
      return_acks => analyze_packet_return_acks,
      call_data  => analyze_packet_call_data,
      call_tag  => analyze_packet_call_tag,
      return_tag  => analyze_packet_return_tag,
      call_mtag => analyze_packet_tag_in,
      return_mtag => analyze_packet_tag_out,
      return_data =>analyze_packet_return_data,
      call_mreq => analyze_packet_start_req,
      call_mack => analyze_packet_start_ack,
      return_mreq => analyze_packet_fin_req,
      return_mack => analyze_packet_fin_ack,
      call_mdata => analyze_packet_in_args,
      return_mdata => analyze_packet_out_args,
      clk => clk, 
      reset => reset --
    ); --
  analyze_packet_instance:analyze_packet-- 
    generic map(tag_length => 1)
    port map(-- 
      pkt => analyze_packet_pkt,
      buf => analyze_packet_buf,
      wlen => analyze_packet_wlen,
      blen => analyze_packet_blen,
      start_req => analyze_packet_start_req,
      start_ack => analyze_packet_start_ack,
      fin_req => analyze_packet_fin_req,
      fin_ack => analyze_packet_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(1 downto 1),
      memory_space_5_lr_ack => memory_space_5_lr_ack(1 downto 1),
      memory_space_5_lr_addr => memory_space_5_lr_addr(31 downto 16),
      memory_space_5_lr_tag => memory_space_5_lr_tag(21 downto 11),
      memory_space_5_lc_req => memory_space_5_lc_req(1 downto 1),
      memory_space_5_lc_ack => memory_space_5_lc_ack(1 downto 1),
      memory_space_5_lc_data => memory_space_5_lc_data(15 downto 8),
      memory_space_5_lc_tag => memory_space_5_lc_tag(9 downto 5),
      tag_in => analyze_packet_tag_in,
      tag_out => analyze_packet_tag_out-- 
    ); -- 
  -- module click_bc_storage_initializer_x
  -- call arbiter for module click_bc_storage_initializer_x
  click_bc_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => click_bc_storage_initializer_x_call_reqs,
      call_acks => click_bc_storage_initializer_x_call_acks,
      return_reqs => click_bc_storage_initializer_x_return_reqs,
      return_acks => click_bc_storage_initializer_x_return_acks,
      call_tag  => click_bc_storage_initializer_x_call_tag,
      return_tag  => click_bc_storage_initializer_x_return_tag,
      call_mtag => click_bc_storage_initializer_x_tag_in,
      return_mtag => click_bc_storage_initializer_x_tag_out,
      call_mreq => click_bc_storage_initializer_x_start_req,
      call_mack => click_bc_storage_initializer_x_start_ack,
      return_mreq => click_bc_storage_initializer_x_fin_req,
      return_mack => click_bc_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  click_bc_storage_initializer_x_instance:click_bc_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => click_bc_storage_initializer_x_start_req,
      start_ack => click_bc_storage_initializer_x_start_ack,
      fin_req => click_bc_storage_initializer_x_fin_req,
      fin_ack => click_bc_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      GV_15_initializer_in_click_bc_call_reqs => GV_15_initializer_in_click_bc_call_reqs(0 downto 0),
      GV_15_initializer_in_click_bc_call_acks => GV_15_initializer_in_click_bc_call_acks(0 downto 0),
      GV_15_initializer_in_click_bc_call_tag => GV_15_initializer_in_click_bc_call_tag(0 downto 0),
      GV_15_initializer_in_click_bc_return_reqs => GV_15_initializer_in_click_bc_return_reqs(0 downto 0),
      GV_15_initializer_in_click_bc_return_acks => GV_15_initializer_in_click_bc_return_acks(0 downto 0),
      GV_15_initializer_in_click_bc_return_tag => GV_15_initializer_in_click_bc_return_tag(0 downto 0),
      GV_16_initializer_in_click_bc_call_reqs => GV_16_initializer_in_click_bc_call_reqs(0 downto 0),
      GV_16_initializer_in_click_bc_call_acks => GV_16_initializer_in_click_bc_call_acks(0 downto 0),
      GV_16_initializer_in_click_bc_call_tag => GV_16_initializer_in_click_bc_call_tag(0 downto 0),
      GV_16_initializer_in_click_bc_return_reqs => GV_16_initializer_in_click_bc_return_reqs(0 downto 0),
      GV_16_initializer_in_click_bc_return_acks => GV_16_initializer_in_click_bc_return_acks(0 downto 0),
      GV_16_initializer_in_click_bc_return_tag => GV_16_initializer_in_click_bc_return_tag(0 downto 0),
      tag_in => click_bc_storage_initializer_x_tag_in,
      tag_out => click_bc_storage_initializer_x_tag_out-- 
    ); -- 
  -- module free_queue_init
  -- call arbiter for module free_queue_init
  free_queue_init_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => free_queue_init_call_reqs,
      call_acks => free_queue_init_call_acks,
      return_reqs => free_queue_init_return_reqs,
      return_acks => free_queue_init_return_acks,
      call_tag  => free_queue_init_call_tag,
      return_tag  => free_queue_init_return_tag,
      call_mtag => free_queue_init_tag_in,
      return_mtag => free_queue_init_tag_out,
      call_mreq => free_queue_init_start_req,
      call_mack => free_queue_init_start_ack,
      return_mreq => free_queue_init_fin_req,
      return_mack => free_queue_init_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  free_queue_init_instance:free_queue_init-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => free_queue_init_start_req,
      start_ack => free_queue_init_start_ack,
      fin_req => free_queue_init_fin_req,
      fin_ack => free_queue_init_fin_ack,
      clk => clk,
      reset => reset,
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(1 downto 1),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(1 downto 1),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(63 downto 32),
      tag_in => free_queue_init_tag_in,
      tag_out => free_queue_init_tag_out-- 
    ); -- 
  -- module global_storage_initializer_x
  -- call arbiter for module global_storage_initializer_x
  global_storage_initializer_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => global_storage_initializer_x_call_reqs,
      call_acks => global_storage_initializer_x_call_acks,
      return_reqs => global_storage_initializer_x_return_reqs,
      return_acks => global_storage_initializer_x_return_acks,
      call_tag  => global_storage_initializer_x_call_tag,
      return_tag  => global_storage_initializer_x_return_tag,
      call_mtag => global_storage_initializer_x_tag_in,
      return_mtag => global_storage_initializer_x_tag_out,
      call_mreq => global_storage_initializer_x_start_req,
      call_mack => global_storage_initializer_x_start_ack,
      return_mreq => global_storage_initializer_x_fin_req,
      return_mack => global_storage_initializer_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  global_storage_initializer_x_instance:global_storage_initializer_x-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => global_storage_initializer_x_start_req,
      start_ack => global_storage_initializer_x_start_ack,
      fin_req => global_storage_initializer_x_fin_req,
      fin_ack => global_storage_initializer_x_fin_ack,
      clk => clk,
      reset => reset,
      click_bc_storage_initializer_x_call_reqs => click_bc_storage_initializer_x_call_reqs(0 downto 0),
      click_bc_storage_initializer_x_call_acks => click_bc_storage_initializer_x_call_acks(0 downto 0),
      click_bc_storage_initializer_x_call_tag => click_bc_storage_initializer_x_call_tag(0 downto 0),
      click_bc_storage_initializer_x_return_reqs => click_bc_storage_initializer_x_return_reqs(0 downto 0),
      click_bc_storage_initializer_x_return_acks => click_bc_storage_initializer_x_return_acks(0 downto 0),
      click_bc_storage_initializer_x_return_tag => click_bc_storage_initializer_x_return_tag(0 downto 0),
      tag_in => global_storage_initializer_x_tag_in,
      tag_out => global_storage_initializer_x_tag_out-- 
    ); -- 
  -- module receive_packet_pipeline
  receive_packet_pipeline_instance:receive_packet_pipeline-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => receive_packet_pipeline_start_req,
      start_ack => receive_packet_pipeline_start_ack,
      fin_req => receive_packet_pipeline_fin_req,
      fin_ack => receive_packet_pipeline_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_sr_req => memory_space_5_sr_req(0 downto 0),
      memory_space_5_sr_ack => memory_space_5_sr_ack(0 downto 0),
      memory_space_5_sr_addr => memory_space_5_sr_addr(15 downto 0),
      memory_space_5_sr_data => memory_space_5_sr_data(7 downto 0),
      memory_space_5_sr_tag => memory_space_5_sr_tag(10 downto 0),
      memory_space_5_sc_req => memory_space_5_sc_req(0 downto 0),
      memory_space_5_sc_ack => memory_space_5_sc_ack(0 downto 0),
      memory_space_5_sc_tag => memory_space_5_sc_tag(4 downto 0),
      free_queue_pipe_pipe_read_req => free_queue_pipe_pipe_read_req(0 downto 0),
      free_queue_pipe_pipe_read_ack => free_queue_pipe_pipe_read_ack(0 downto 0),
      free_queue_pipe_pipe_read_data => free_queue_pipe_pipe_read_data(31 downto 0),
      in_ctrl_pipe_read_req => in_ctrl_pipe_read_req(0 downto 0),
      in_ctrl_pipe_read_ack => in_ctrl_pipe_read_ack(0 downto 0),
      in_ctrl_pipe_read_data => in_ctrl_pipe_read_data(7 downto 0),
      in_data_pipe_read_req => in_data_pipe_read_req(0 downto 0),
      in_data_pipe_read_ack => in_data_pipe_read_ack(0 downto 0),
      in_data_pipe_read_data => in_data_pipe_read_data(63 downto 0),
      receive_packet_buf_queue_pipe_read_req => receive_packet_buf_queue_pipe_read_req(0 downto 0),
      receive_packet_buf_queue_pipe_read_ack => receive_packet_buf_queue_pipe_read_ack(0 downto 0),
      receive_packet_buf_queue_pipe_read_data => receive_packet_buf_queue_pipe_read_data(31 downto 0),
      swapped_in_data_pipe_read_req => swapped_in_data_pipe_read_req(0 downto 0),
      swapped_in_data_pipe_read_ack => swapped_in_data_pipe_read_ack(0 downto 0),
      swapped_in_data_pipe_read_data => swapped_in_data_pipe_read_data(63 downto 0),
      receive_packet_buf_queue_pipe_write_req => receive_packet_buf_queue_pipe_write_req(0 downto 0),
      receive_packet_buf_queue_pipe_write_ack => receive_packet_buf_queue_pipe_write_ack(0 downto 0),
      receive_packet_buf_queue_pipe_write_data => receive_packet_buf_queue_pipe_write_data(31 downto 0),
      swapped_in_data_pipe_write_req => swapped_in_data_pipe_write_req(0 downto 0),
      swapped_in_data_pipe_write_ack => swapped_in_data_pipe_write_ack(0 downto 0),
      swapped_in_data_pipe_write_data => swapped_in_data_pipe_write_data(63 downto 0),
      receive_packet_pipe_pipe_write_req => receive_packet_pipe_pipe_write_req(0 downto 0),
      receive_packet_pipe_pipe_write_ack => receive_packet_pipe_pipe_write_ack(0 downto 0),
      receive_packet_pipe_pipe_write_data => receive_packet_pipe_pipe_write_data(31 downto 0),
      tag_in => receive_packet_pipeline_tag_in,
      tag_out => receive_packet_pipeline_tag_out-- 
    ); -- 
  -- module will be run forever 
  receive_packet_pipeline_tag_in <= (others => '0');
  receive_packet_pipeline_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => receive_packet_pipeline_start_req, start_ack => receive_packet_pipeline_start_ack,  fin_req => receive_packet_pipeline_fin_req,  fin_ack => receive_packet_pipeline_fin_ack);
  -- module send_packet_pipeline
  send_packet_pipeline_instance:send_packet_pipeline-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => send_packet_pipeline_start_req,
      start_ack => send_packet_pipeline_start_ack,
      fin_req => send_packet_pipeline_fin_req,
      fin_ack => send_packet_pipeline_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_5_lr_req => memory_space_5_lr_req(0 downto 0),
      memory_space_5_lr_ack => memory_space_5_lr_ack(0 downto 0),
      memory_space_5_lr_addr => memory_space_5_lr_addr(15 downto 0),
      memory_space_5_lr_tag => memory_space_5_lr_tag(10 downto 0),
      memory_space_5_lc_req => memory_space_5_lc_req(0 downto 0),
      memory_space_5_lc_ack => memory_space_5_lc_ack(0 downto 0),
      memory_space_5_lc_data => memory_space_5_lc_data(7 downto 0),
      memory_space_5_lc_tag => memory_space_5_lc_tag(4 downto 0),
      send_packet_buf_queue_pipe_read_req => send_packet_buf_queue_pipe_read_req(0 downto 0),
      send_packet_buf_queue_pipe_read_ack => send_packet_buf_queue_pipe_read_ack(0 downto 0),
      send_packet_buf_queue_pipe_read_data => send_packet_buf_queue_pipe_read_data(31 downto 0),
      send_packet_pipe_pipe_read_req => send_packet_pipe_pipe_read_req(0 downto 0),
      send_packet_pipe_pipe_read_ack => send_packet_pipe_pipe_read_ack(0 downto 0),
      send_packet_pipe_pipe_read_data => send_packet_pipe_pipe_read_data(31 downto 0),
      free_queue_pipe_pipe_write_req => free_queue_pipe_pipe_write_req(0 downto 0),
      free_queue_pipe_pipe_write_ack => free_queue_pipe_pipe_write_ack(0 downto 0),
      free_queue_pipe_pipe_write_data => free_queue_pipe_pipe_write_data(31 downto 0),
      out_ctrl_pipe_write_req => out_ctrl_pipe_write_req(0 downto 0),
      out_ctrl_pipe_write_ack => out_ctrl_pipe_write_ack(0 downto 0),
      out_ctrl_pipe_write_data => out_ctrl_pipe_write_data(7 downto 0),
      out_data_pipe_write_req => out_data_pipe_write_req(0 downto 0),
      out_data_pipe_write_ack => out_data_pipe_write_ack(0 downto 0),
      out_data_pipe_write_data => out_data_pipe_write_data(63 downto 0),
      send_packet_buf_queue_pipe_write_req => send_packet_buf_queue_pipe_write_req(0 downto 0),
      send_packet_buf_queue_pipe_write_ack => send_packet_buf_queue_pipe_write_ack(0 downto 0),
      send_packet_buf_queue_pipe_write_data => send_packet_buf_queue_pipe_write_data(31 downto 0),
      analyze_packet_call_reqs => analyze_packet_call_reqs(0 downto 0),
      analyze_packet_call_acks => analyze_packet_call_acks(0 downto 0),
      analyze_packet_call_data => analyze_packet_call_data(31 downto 0),
      analyze_packet_call_tag => analyze_packet_call_tag(0 downto 0),
      analyze_packet_return_reqs => analyze_packet_return_reqs(0 downto 0),
      analyze_packet_return_acks => analyze_packet_return_acks(0 downto 0),
      analyze_packet_return_data => analyze_packet_return_data(63 downto 0),
      analyze_packet_return_tag => analyze_packet_return_tag(0 downto 0),
      tag_in => send_packet_pipeline_tag_in,
      tag_out => send_packet_pipeline_tag_out-- 
    ); -- 
  -- module will be run forever 
  send_packet_pipeline_tag_in <= (others => '0');
  send_packet_pipeline_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => send_packet_pipeline_start_req, start_ack => send_packet_pipeline_start_ack,  fin_req => send_packet_pipeline_fin_req,  fin_ack => send_packet_pipeline_fin_ack);
  -- module wrapper_input
  wrapper_input_instance:wrapper_input-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_input_start_req,
      start_ack => wrapper_input_start_ack,
      fin_req => wrapper_input_fin_req,
      fin_ack => wrapper_input_fin_ack,
      clk => clk,
      reset => reset,
      receive_packet_pipe_pipe_read_req => receive_packet_pipe_pipe_read_req(0 downto 0),
      receive_packet_pipe_pipe_read_ack => receive_packet_pipe_pipe_read_ack(0 downto 0),
      receive_packet_pipe_pipe_read_data => receive_packet_pipe_pipe_read_data(31 downto 0),
      src_in0_pipe_write_req => src_in0_pipe_write_req(0 downto 0),
      src_in0_pipe_write_ack => src_in0_pipe_write_ack(0 downto 0),
      src_in0_pipe_write_data => src_in0_pipe_write_data(31 downto 0),
      free_queue_init_call_reqs => free_queue_init_call_reqs(0 downto 0),
      free_queue_init_call_acks => free_queue_init_call_acks(0 downto 0),
      free_queue_init_call_tag => free_queue_init_call_tag(0 downto 0),
      free_queue_init_return_reqs => free_queue_init_return_reqs(0 downto 0),
      free_queue_init_return_acks => free_queue_init_return_acks(0 downto 0),
      free_queue_init_return_tag => free_queue_init_return_tag(0 downto 0),
      global_storage_initializer_x_call_reqs => global_storage_initializer_x_call_reqs(0 downto 0),
      global_storage_initializer_x_call_acks => global_storage_initializer_x_call_acks(0 downto 0),
      global_storage_initializer_x_call_tag => global_storage_initializer_x_call_tag(0 downto 0),
      global_storage_initializer_x_return_reqs => global_storage_initializer_x_return_reqs(0 downto 0),
      global_storage_initializer_x_return_acks => global_storage_initializer_x_return_acks(0 downto 0),
      global_storage_initializer_x_return_tag => global_storage_initializer_x_return_tag(0 downto 0),
      tag_in => wrapper_input_tag_in,
      tag_out => wrapper_input_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_input_tag_in <= (others => '0');
  wrapper_input_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_input_start_req, start_ack => wrapper_input_start_ack,  fin_req => wrapper_input_fin_req,  fin_ack => wrapper_input_fin_ack);
  -- module wrapper_output
  wrapper_output_instance:wrapper_output-- 
    generic map(tag_length => 1)
    port map(-- 
      start_req => wrapper_output_start_req,
      start_ack => wrapper_output_start_ack,
      fin_req => wrapper_output_fin_req,
      fin_ack => wrapper_output_fin_ack,
      clk => clk,
      reset => reset,
      tofpga0_out0_pipe_read_req => tofpga0_out0_pipe_read_req(0 downto 0),
      tofpga0_out0_pipe_read_ack => tofpga0_out0_pipe_read_ack(0 downto 0),
      tofpga0_out0_pipe_read_data => tofpga0_out0_pipe_read_data(31 downto 0),
      tofpga1_out0_pipe_read_req => tofpga1_out0_pipe_read_req(0 downto 0),
      tofpga1_out0_pipe_read_ack => tofpga1_out0_pipe_read_ack(0 downto 0),
      tofpga1_out0_pipe_read_data => tofpga1_out0_pipe_read_data(31 downto 0),
      tofpga2_out0_pipe_read_req => tofpga2_out0_pipe_read_req(0 downto 0),
      tofpga2_out0_pipe_read_ack => tofpga2_out0_pipe_read_ack(0 downto 0),
      tofpga2_out0_pipe_read_data => tofpga2_out0_pipe_read_data(31 downto 0),
      tofpga3_out0_pipe_read_req => tofpga3_out0_pipe_read_req(0 downto 0),
      tofpga3_out0_pipe_read_ack => tofpga3_out0_pipe_read_ack(0 downto 0),
      tofpga3_out0_pipe_read_data => tofpga3_out0_pipe_read_data(31 downto 0),
      tofpga_port_number_pipe_read_req => tofpga_port_number_pipe_read_req(0 downto 0),
      tofpga_port_number_pipe_read_ack => tofpga_port_number_pipe_read_ack(0 downto 0),
      tofpga_port_number_pipe_read_data => tofpga_port_number_pipe_read_data(31 downto 0),
      send_packet_pipe_pipe_write_req => send_packet_pipe_pipe_write_req(0 downto 0),
      send_packet_pipe_pipe_write_ack => send_packet_pipe_pipe_write_ack(0 downto 0),
      send_packet_pipe_pipe_write_data => send_packet_pipe_pipe_write_data(31 downto 0),
      tag_in => wrapper_output_tag_in,
      tag_out => wrapper_output_tag_out-- 
    ); -- 
  -- module will be run forever 
  wrapper_output_tag_in <= (others => '0');
  wrapper_output_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => wrapper_output_start_req, start_ack => wrapper_output_start_ack,  fin_req => wrapper_output_fin_req,  fin_ack => wrapper_output_fin_ack);
  chk_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 2,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => chk_in0_pipe_read_req,
      read_ack => chk_in0_pipe_read_ack,
      read_data => chk_in0_pipe_read_data,
      write_req => chk_in0_pipe_write_req,
      write_ack => chk_in0_pipe_write_ack,
      write_data => chk_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  free_queue_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 5,
      data_width => 32,
      depth => 16 --
    )
    port map( -- 
      read_req => free_queue_pipe_pipe_read_req,
      read_ack => free_queue_pipe_pipe_read_ack,
      read_data => free_queue_pipe_pipe_read_data,
      write_req => free_queue_pipe_pipe_write_req,
      write_ack => free_queue_pipe_pipe_write_ack,
      write_data => free_queue_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => in_ctrl_pipe_read_req,
      read_ack => in_ctrl_pipe_read_ack,
      read_data => in_ctrl_pipe_read_data,
      write_req => in_ctrl_pipe_write_req,
      write_ack => in_ctrl_pipe_write_ack,
      write_data => in_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_read_req,
      read_ack => in_data_pipe_read_ack,
      read_data => in_data_pipe_read_data,
      write_req => in_data_pipe_write_req,
      write_ack => in_data_pipe_write_ack,
      write_data => in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_ctrl_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 8,
      depth => 1 --
    )
    port map( -- 
      read_req => out_ctrl_pipe_read_req,
      read_ack => out_ctrl_pipe_read_ack,
      read_data => out_ctrl_pipe_read_data,
      write_req => out_ctrl_pipe_write_req,
      write_ack => out_ctrl_pipe_write_ack,
      write_data => out_ctrl_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_read_req,
      read_ack => out_data_pipe_read_ack,
      read_data => out_data_pipe_read_data,
      write_req => out_data_pipe_write_req,
      write_ack => out_data_pipe_write_ack,
      write_data => out_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  receive_packet_buf_queue_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 8 --
    )
    port map( -- 
      read_req => receive_packet_buf_queue_pipe_read_req,
      read_ack => receive_packet_buf_queue_pipe_read_ack,
      read_data => receive_packet_buf_queue_pipe_read_data,
      write_req => receive_packet_buf_queue_pipe_write_req,
      write_ack => receive_packet_buf_queue_pipe_write_ack,
      write_data => receive_packet_buf_queue_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  receive_packet_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => receive_packet_pipe_pipe_read_req,
      read_ack => receive_packet_pipe_pipe_read_ack,
      read_data => receive_packet_pipe_pipe_read_data,
      write_req => receive_packet_pipe_pipe_write_req,
      write_ack => receive_packet_pipe_pipe_write_ack,
      write_data => receive_packet_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  rtt_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 2,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => rtt_in0_pipe_read_req,
      read_ack => rtt_in0_pipe_read_ack,
      read_data => rtt_in0_pipe_read_data,
      write_req => rtt_in0_pipe_write_req,
      write_ack => rtt_in0_pipe_write_ack,
      write_data => rtt_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  send_packet_buf_queue_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 8 --
    )
    port map( -- 
      read_req => send_packet_buf_queue_pipe_read_req,
      read_ack => send_packet_buf_queue_pipe_read_ack,
      read_data => send_packet_buf_queue_pipe_read_data,
      write_req => send_packet_buf_queue_pipe_write_req,
      write_ack => send_packet_buf_queue_pipe_write_ack,
      write_data => send_packet_buf_queue_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  send_packet_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => send_packet_pipe_pipe_read_req,
      read_ack => send_packet_pipe_pipe_read_ack,
      read_data => send_packet_pipe_pipe_read_data,
      write_req => send_packet_pipe_pipe_write_req,
      write_ack => send_packet_pipe_pipe_write_ack,
      write_data => send_packet_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  src_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => src_in0_pipe_read_req,
      read_ack => src_in0_pipe_read_ack,
      read_data => src_in0_pipe_read_data,
      write_req => src_in0_pipe_write_req,
      write_ack => src_in0_pipe_write_ack,
      write_data => src_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  swapped_in_data_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 64,
      depth => 2 --
    )
    port map( -- 
      read_req => swapped_in_data_pipe_read_req,
      read_ack => swapped_in_data_pipe_read_ack,
      read_data => swapped_in_data_pipe_read_data,
      write_req => swapped_in_data_pipe_write_req,
      write_ack => swapped_in_data_pipe_write_ack,
      write_data => swapped_in_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to0_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to0_in0_pipe_read_req,
      read_ack => to0_in0_pipe_read_ack,
      read_data => to0_in0_pipe_read_data,
      write_req => to0_in0_pipe_write_req,
      write_ack => to0_in0_pipe_write_ack,
      write_data => to0_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to1_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to1_in0_pipe_read_req,
      read_ack => to1_in0_pipe_read_ack,
      read_data => to1_in0_pipe_read_data,
      write_req => to1_in0_pipe_write_req,
      write_ack => to1_in0_pipe_write_ack,
      write_data => to1_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to2_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to2_in0_pipe_read_req,
      read_ack => to2_in0_pipe_read_ack,
      read_data => to2_in0_pipe_read_data,
      write_req => to2_in0_pipe_write_req,
      write_ack => to2_in0_pipe_write_ack,
      write_data => to2_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  to3_in0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => to3_in0_pipe_read_req,
      read_ack => to3_in0_pipe_read_ack,
      read_data => to3_in0_pipe_read_data,
      write_req => to3_in0_pipe_write_req,
      write_ack => to3_in0_pipe_write_ack,
      write_data => to3_in0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga0_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga0_out0_pipe_read_req,
      read_ack => tofpga0_out0_pipe_read_ack,
      read_data => tofpga0_out0_pipe_read_data,
      write_req => tofpga0_out0_pipe_write_req,
      write_ack => tofpga0_out0_pipe_write_ack,
      write_data => tofpga0_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga1_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga1_out0_pipe_read_req,
      read_ack => tofpga1_out0_pipe_read_ack,
      read_data => tofpga1_out0_pipe_read_data,
      write_req => tofpga1_out0_pipe_write_req,
      write_ack => tofpga1_out0_pipe_write_ack,
      write_data => tofpga1_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga2_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga2_out0_pipe_read_req,
      read_ack => tofpga2_out0_pipe_read_ack,
      read_data => tofpga2_out0_pipe_read_data,
      write_req => tofpga2_out0_pipe_write_req,
      write_ack => tofpga2_out0_pipe_write_ack,
      write_data => tofpga2_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga3_out0_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga3_out0_pipe_read_req,
      read_ack => tofpga3_out0_pipe_read_ack,
      read_data => tofpga3_out0_pipe_read_data,
      write_req => tofpga3_out0_pipe_write_req,
      write_ack => tofpga3_out0_pipe_write_ack,
      write_data => tofpga3_out0_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  tofpga_port_number_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 4,
      data_width => 32,
      depth => 1 --
    )
    port map( -- 
      read_req => tofpga_port_number_pipe_read_req,
      read_ack => tofpga_port_number_pipe_read_ack,
      read_data => tofpga_port_number_pipe_read_data,
      write_req => tofpga_port_number_pipe_write_req,
      write_ack => tofpga_port_number_pipe_write_ack,
      write_data => tofpga_port_number_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 9,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 9,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 5,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 5,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_3: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 14,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 14,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_3_lr_addr,
      lr_req_in => memory_space_3_lr_req,
      lr_ack_out => memory_space_3_lr_ack,
      lr_tag_in => memory_space_3_lr_tag,
      lc_req_in => memory_space_3_lc_req,
      lc_ack_out => memory_space_3_lc_ack,
      lc_data_out => memory_space_3_lc_data,
      lc_tag_out => memory_space_3_lc_tag,
      sr_addr_in => memory_space_3_sr_addr,
      sr_data_in => memory_space_3_sr_data,
      sr_req_in => memory_space_3_sr_req,
      sr_ack_out => memory_space_3_sr_ack,
      sr_tag_in => memory_space_3_sr_tag,
      sc_req_in=> memory_space_3_sc_req,
      sc_ack_out => memory_space_3_sc_ack,
      sc_tag_out => memory_space_3_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_4: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 1,
      data_width => 32,
      tag_width => 1,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 1,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_4_lr_addr,
      lr_req_in => memory_space_4_lr_req,
      lr_ack_out => memory_space_4_lr_ack,
      lr_tag_in => memory_space_4_lr_tag,
      lc_req_in => memory_space_4_lc_req,
      lc_ack_out => memory_space_4_lc_ack,
      lc_data_out => memory_space_4_lc_data,
      lc_tag_out => memory_space_4_lc_tag,
      sr_addr_in => memory_space_4_sr_addr,
      sr_data_in => memory_space_4_sr_data,
      sr_req_in => memory_space_4_sr_req,
      sr_ack_out => memory_space_4_sr_ack,
      sr_tag_in => memory_space_4_sr_tag,
      sc_req_in=> memory_space_4_sc_req,
      sc_ack_out => memory_space_4_sc_ack,
      sc_tag_out => memory_space_4_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_5: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 10,
      num_stores => 8,
      addr_width => 16,
      data_width => 8,
      tag_width => 5,
      time_stamp_width => 6,
      number_of_banks => 2,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 15,
      base_bank_data_width => 8
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_5_lr_addr,
      lr_req_in => memory_space_5_lr_req,
      lr_ack_out => memory_space_5_lr_ack,
      lr_tag_in => memory_space_5_lr_tag,
      lc_req_in => memory_space_5_lc_req,
      lc_ack_out => memory_space_5_lc_ack,
      lc_data_out => memory_space_5_lc_data,
      lc_tag_out => memory_space_5_lc_tag,
      sr_addr_in => memory_space_5_sr_addr,
      sr_data_in => memory_space_5_sr_data,
      sr_req_in => memory_space_5_sr_req,
      sr_ack_out => memory_space_5_sr_ack,
      sr_tag_in => memory_space_5_sr_tag,
      sc_req_in=> memory_space_5_sc_req,
      sc_ack_out => memory_space_5_sc_ack,
      sc_tag_out => memory_space_5_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
library work;
use work.vc_system_package.all;
entity ahir_system_Test_Bench is -- 
  -- 
end entity;
architecture Default of ahir_system_Test_Bench is -- 
  component ahir_system is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      in_ctrl_pipe_write_data: in std_logic_vector(7 downto 0);
      in_ctrl_pipe_write_req : in std_logic_vector(0 downto 0);
      in_ctrl_pipe_write_ack : out std_logic_vector(0 downto 0);
      in_data_pipe_write_data: in std_logic_vector(63 downto 0);
      in_data_pipe_write_req : in std_logic_vector(0 downto 0);
      in_data_pipe_write_ack : out std_logic_vector(0 downto 0);
      out_ctrl_pipe_read_data: out std_logic_vector(7 downto 0);
      out_ctrl_pipe_read_req : in std_logic_vector(0 downto 0);
      out_ctrl_pipe_read_ack : out std_logic_vector(0 downto 0);
      out_data_pipe_read_data: out std_logic_vector(63 downto 0);
      out_data_pipe_read_req : in std_logic_vector(0 downto 0);
      out_data_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  signal clk: std_logic := '0';
  signal reset: std_logic := '1';
  signal ahir_glue_chk_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_start_req : std_logic := '0';
  signal ahir_glue_chk_start_ack : std_logic := '0';
  signal ahir_glue_chk_fin_req   : std_logic := '0';
  signal ahir_glue_chk_fin_ack   : std_logic := '0';
  signal ahir_glue_chk_1_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_1_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_chk_1_start_req : std_logic := '0';
  signal ahir_glue_chk_1_start_ack : std_logic := '0';
  signal ahir_glue_chk_1_fin_req   : std_logic := '0';
  signal ahir_glue_chk_1_fin_ack   : std_logic := '0';
  signal ahir_glue_rtt_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_rtt_start_req : std_logic := '0';
  signal ahir_glue_rtt_start_ack : std_logic := '0';
  signal ahir_glue_rtt_fin_req   : std_logic := '0';
  signal ahir_glue_rtt_fin_ack   : std_logic := '0';
  signal ahir_glue_src_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_src_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_src_start_req : std_logic := '0';
  signal ahir_glue_src_start_ack : std_logic := '0';
  signal ahir_glue_src_fin_req   : std_logic := '0';
  signal ahir_glue_src_fin_ack   : std_logic := '0';
  signal ahir_glue_to0_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to0_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to0_start_req : std_logic := '0';
  signal ahir_glue_to0_start_ack : std_logic := '0';
  signal ahir_glue_to0_fin_req   : std_logic := '0';
  signal ahir_glue_to0_fin_ack   : std_logic := '0';
  signal ahir_glue_to1_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to1_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to1_start_req : std_logic := '0';
  signal ahir_glue_to1_start_ack : std_logic := '0';
  signal ahir_glue_to1_fin_req   : std_logic := '0';
  signal ahir_glue_to1_fin_ack   : std_logic := '0';
  signal ahir_glue_to2_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to2_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to2_start_req : std_logic := '0';
  signal ahir_glue_to2_start_ack : std_logic := '0';
  signal ahir_glue_to2_fin_req   : std_logic := '0';
  signal ahir_glue_to2_fin_ack   : std_logic := '0';
  signal ahir_glue_to3_tag_in: std_logic_vector(0 downto 0);
  signal ahir_glue_to3_tag_out: std_logic_vector(0 downto 0);
  signal ahir_glue_to3_start_req : std_logic := '0';
  signal ahir_glue_to3_start_ack : std_logic := '0';
  signal ahir_glue_to3_fin_req   : std_logic := '0';
  signal ahir_glue_to3_fin_ack   : std_logic := '0';
  signal receive_packet_pipeline_tag_in: std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_tag_out: std_logic_vector(0 downto 0);
  signal receive_packet_pipeline_start_req : std_logic := '0';
  signal receive_packet_pipeline_start_ack : std_logic := '0';
  signal receive_packet_pipeline_fin_req   : std_logic := '0';
  signal receive_packet_pipeline_fin_ack   : std_logic := '0';
  signal send_packet_pipeline_tag_in: std_logic_vector(0 downto 0);
  signal send_packet_pipeline_tag_out: std_logic_vector(0 downto 0);
  signal send_packet_pipeline_start_req : std_logic := '0';
  signal send_packet_pipeline_start_ack : std_logic := '0';
  signal send_packet_pipeline_fin_req   : std_logic := '0';
  signal send_packet_pipeline_fin_ack   : std_logic := '0';
  signal wrapper_input_tag_in: std_logic_vector(0 downto 0);
  signal wrapper_input_tag_out: std_logic_vector(0 downto 0);
  signal wrapper_input_start_req : std_logic := '0';
  signal wrapper_input_start_ack : std_logic := '0';
  signal wrapper_input_fin_req   : std_logic := '0';
  signal wrapper_input_fin_ack   : std_logic := '0';
  signal wrapper_output_tag_in: std_logic_vector(0 downto 0);
  signal wrapper_output_tag_out: std_logic_vector(0 downto 0);
  signal wrapper_output_start_req : std_logic := '0';
  signal wrapper_output_start_ack : std_logic := '0';
  signal wrapper_output_fin_req   : std_logic := '0';
  signal wrapper_output_fin_ack   : std_logic := '0';
  -- write to pipe in_ctrl
  signal in_ctrl_pipe_write_data: std_logic_vector(7 downto 0);
  signal in_ctrl_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal in_ctrl_pipe_write_ack : std_logic_vector(0 downto 0);
  -- write to pipe in_data
  signal in_data_pipe_write_data: std_logic_vector(63 downto 0);
  signal in_data_pipe_write_req : std_logic_vector(0 downto 0) := (others => '0');
  signal in_data_pipe_write_ack : std_logic_vector(0 downto 0);
  -- read from pipe out_ctrl
  signal out_ctrl_pipe_read_data: std_logic_vector(7 downto 0);
  signal out_ctrl_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal out_ctrl_pipe_read_ack : std_logic_vector(0 downto 0);
  -- read from pipe out_data
  signal out_data_pipe_read_data: std_logic_vector(63 downto 0);
  signal out_data_pipe_read_req : std_logic_vector(0 downto 0) := (others => '0');
  signal out_data_pipe_read_ack : std_logic_vector(0 downto 0);
  -- 
begin --
  -- clock/reset generation 
  clk <= not clk after 5 ns;
  process
  begin --
    wait until clk = '1';
    reset <= '0';
    wait;
    --
  end process;
  -- a rudimentary tb.. will start all the top-level modules ..
  ahir_system_instance: ahir_system -- 
    port map ( -- 
      clk => clk,
      reset => reset,
      in_ctrl_pipe_write_data  => in_ctrl_pipe_write_data, 
      in_ctrl_pipe_write_req  => in_ctrl_pipe_write_req, 
      in_ctrl_pipe_write_ack  => in_ctrl_pipe_write_ack,
      in_data_pipe_write_data  => in_data_pipe_write_data, 
      in_data_pipe_write_req  => in_data_pipe_write_req, 
      in_data_pipe_write_ack  => in_data_pipe_write_ack,
      out_ctrl_pipe_read_data  => out_ctrl_pipe_read_data, 
      out_ctrl_pipe_read_req  => out_ctrl_pipe_read_req, 
      out_ctrl_pipe_read_ack  => out_ctrl_pipe_read_ack ,
      out_data_pipe_read_data  => out_data_pipe_read_data, 
      out_data_pipe_read_req  => out_data_pipe_read_req, 
      out_data_pipe_read_ack  => out_data_pipe_read_ack ); -- 
  -- 
end Default;
