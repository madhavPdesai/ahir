-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity vectorSum is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_1_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_0_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_sc_tag :  in  std_logic_vector(3 downto 0);
    in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
    out_data_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    out_data_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    out_data_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
    x_vectorSum_x_call_reqs : out  std_logic_vector(0 downto 0);
    x_vectorSum_x_call_acks : in   std_logic_vector(0 downto 0);
    x_vectorSum_x_call_tag  :  out  std_logic_vector(0 downto 0);
    x_vectorSum_x_return_reqs : out  std_logic_vector(0 downto 0);
    x_vectorSum_x_return_acks : in   std_logic_vector(0 downto 0);
    x_vectorSum_x_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity vectorSum;
architecture Default of vectorSum is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal vectorSum_CP_4500_start: Boolean;
  -- links between control-path and data-path
  signal binary_326_inst_req_1 : boolean;
  signal binary_326_inst_ack_1 : boolean;
  signal call_stmt_345_call_req_1 : boolean;
  signal call_stmt_345_call_req_0 : boolean;
  signal call_stmt_345_call_ack_0 : boolean;
  signal array_obj_ref_358_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_358_index_0_resize_req_0 : boolean;
  signal array_obj_ref_358_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_358_root_address_inst_req_0 : boolean;
  signal binary_326_inst_ack_0 : boolean;
  signal binary_326_inst_req_0 : boolean;
  signal array_obj_ref_358_index_0_rename_req_0 : boolean;
  signal array_obj_ref_358_index_0_rename_ack_0 : boolean;
  signal if_stmt_328_branch_req_0 : boolean;
  signal if_stmt_328_branch_ack_1 : boolean;
  signal array_obj_ref_358_offset_inst_req_0 : boolean;
  signal call_stmt_345_call_ack_1 : boolean;
  signal ptr_deref_363_base_resize_req_0 : boolean;
  signal if_stmt_328_branch_ack_0 : boolean;
  signal binary_372_inst_ack_1 : boolean;
  signal binary_372_inst_req_0 : boolean;
  signal ptr_deref_363_root_address_inst_req_0 : boolean;
  signal ptr_deref_363_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_358_offset_inst_ack_0 : boolean;
  signal ptr_deref_363_base_resize_ack_0 : boolean;
  signal ptr_deref_363_addr_0_req_0 : boolean;
  signal ptr_deref_363_load_0_ack_0 : boolean;
  signal simple_obj_ref_365_inst_req_0 : boolean;
  signal simple_obj_ref_365_inst_ack_0 : boolean;
  signal binary_372_inst_ack_0 : boolean;
  signal binary_372_inst_req_1 : boolean;
  signal ptr_deref_363_load_0_ack_1 : boolean;
  signal ptr_deref_363_root_address_inst_ack_0 : boolean;
  signal ptr_deref_363_addr_0_ack_0 : boolean;
  signal ptr_deref_363_load_0_req_1 : boolean;
  signal ptr_deref_363_gather_scatter_req_0 : boolean;
  signal ptr_deref_363_load_0_req_0 : boolean;
  signal addr_of_359_final_reg_ack_0 : boolean;
  signal array_obj_ref_297_index_0_resize_req_0 : boolean;
  signal array_obj_ref_297_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_297_index_0_rename_req_0 : boolean;
  signal array_obj_ref_297_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_297_offset_inst_req_0 : boolean;
  signal array_obj_ref_297_offset_inst_ack_0 : boolean;
  signal array_obj_ref_297_root_address_inst_req_0 : boolean;
  signal array_obj_ref_297_root_address_inst_ack_0 : boolean;
  signal addr_of_298_final_reg_req_0 : boolean;
  signal addr_of_298_final_reg_ack_0 : boolean;
  signal array_obj_ref_302_index_0_resize_req_0 : boolean;
  signal array_obj_ref_302_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_302_index_0_rename_req_0 : boolean;
  signal array_obj_ref_302_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_302_offset_inst_req_0 : boolean;
  signal array_obj_ref_302_offset_inst_ack_0 : boolean;
  signal array_obj_ref_302_root_address_inst_req_0 : boolean;
  signal array_obj_ref_302_root_address_inst_ack_0 : boolean;
  signal addr_of_303_final_reg_req_0 : boolean;
  signal addr_of_303_final_reg_ack_0 : boolean;
  signal simple_obj_ref_306_inst_req_0 : boolean;
  signal simple_obj_ref_306_inst_ack_0 : boolean;
  signal ptr_deref_309_base_resize_req_0 : boolean;
  signal ptr_deref_309_base_resize_ack_0 : boolean;
  signal ptr_deref_309_root_address_inst_req_0 : boolean;
  signal ptr_deref_309_root_address_inst_ack_0 : boolean;
  signal ptr_deref_309_addr_0_req_0 : boolean;
  signal ptr_deref_309_addr_0_ack_0 : boolean;
  signal ptr_deref_309_gather_scatter_req_0 : boolean;
  signal ptr_deref_309_gather_scatter_ack_0 : boolean;
  signal ptr_deref_309_store_0_req_0 : boolean;
  signal ptr_deref_309_store_0_ack_0 : boolean;
  signal ptr_deref_309_store_0_req_1 : boolean;
  signal ptr_deref_309_store_0_ack_1 : boolean;
  signal addr_of_359_final_reg_req_0 : boolean;
  signal ptr_deref_313_base_resize_req_0 : boolean;
  signal ptr_deref_313_base_resize_ack_0 : boolean;
  signal ptr_deref_313_root_address_inst_req_0 : boolean;
  signal ptr_deref_313_root_address_inst_ack_0 : boolean;
  signal ptr_deref_313_addr_0_req_0 : boolean;
  signal ptr_deref_313_addr_0_ack_0 : boolean;
  signal ptr_deref_313_gather_scatter_req_0 : boolean;
  signal ptr_deref_313_gather_scatter_ack_0 : boolean;
  signal ptr_deref_313_store_0_req_0 : boolean;
  signal ptr_deref_313_store_0_ack_0 : boolean;
  signal ptr_deref_313_store_0_req_1 : boolean;
  signal ptr_deref_313_store_0_ack_1 : boolean;
  signal binary_320_inst_req_0 : boolean;
  signal binary_320_inst_ack_0 : boolean;
  signal binary_320_inst_req_1 : boolean;
  signal binary_320_inst_ack_1 : boolean;
  signal binary_378_inst_req_0 : boolean;
  signal binary_378_inst_ack_0 : boolean;
  signal binary_378_inst_req_1 : boolean;
  signal binary_378_inst_ack_1 : boolean;
  signal if_stmt_380_branch_req_0 : boolean;
  signal if_stmt_380_branch_ack_1 : boolean;
  signal if_stmt_380_branch_ack_0 : boolean;
  signal phi_stmt_287_req_0 : boolean;
  signal type_cast_293_inst_req_0 : boolean;
  signal type_cast_293_inst_ack_0 : boolean;
  signal phi_stmt_287_req_1 : boolean;
  signal phi_stmt_287_ack_0 : boolean;
  signal type_cast_338_inst_req_0 : boolean;
  signal type_cast_338_inst_ack_0 : boolean;
  signal phi_stmt_335_req_0 : boolean;
  signal phi_stmt_335_req_1 : boolean;
  signal phi_stmt_335_ack_0 : boolean;
  signal type_cast_354_inst_req_0 : boolean;
  signal type_cast_354_inst_ack_0 : boolean;
  signal phi_stmt_348_req_1 : boolean;
  signal phi_stmt_348_req_0 : boolean;
  signal phi_stmt_348_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 0, backward_delay => 0) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 0, backward_delay => 0) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"vectorSum start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"vectorSum start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"vectorSum fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"vectorSum fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  vectorSum_CP_4500: Block -- control-path 
    signal cp_elements: BooleanArray(121 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(101);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(101), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  output  bypass 
    -- predecessors 
    -- successors 109 
    -- members (15) 
      -- 	$entry
      -- 	branch_block_stmt_282/$entry
      -- 	branch_block_stmt_282/branch_block_stmt_282__entry__
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/$entry
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/$exit
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/$entry
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/$exit
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/$entry
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/$exit
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/req
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/ack
      -- 	branch_block_stmt_282/bb_0_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_req
      -- 
    phi_stmt_287_req_5027_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => phi_stmt_287_req_0); -- 
    -- CP-element group 1 transition  place  output  bypass 
    -- predecessors 22 
    -- successors 23 
    -- members (7) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304__exit__
      -- 	branch_block_stmt_282/assign_stmt_307__entry__
      -- 	branch_block_stmt_282/assign_stmt_307/$entry
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_trigger_
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_active_
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_complete/req
      -- 
    cp_elements(1) <= cp_elements(22);
    req_4629_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1), ack => simple_obj_ref_306_inst_req_0); -- 
    -- CP-element group 2 branch  place  bypass 
    -- predecessors 56 
    -- successors 57 60 
    -- members (2) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327__exit__
      -- 	branch_block_stmt_282/if_stmt_328__entry__
      -- 
    cp_elements(2) <= cp_elements(56);
    -- CP-element group 3 merge  transition  place  output  bypass 
    -- predecessors 113 117 
    -- successors 108 
    -- members (7) 
      -- 	branch_block_stmt_282/merge_stmt_334__exit__
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/req
      -- 
    cp_elements(3) <= OrReduce(cp_elements(113) & cp_elements(117));
    req_5040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(3), ack => type_cast_293_inst_req_0); -- 
    -- CP-element group 4 branch  place  bypass 
    -- predecessors 98 
    -- successors 99 102 
    -- members (2) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379__exit__
      -- 	branch_block_stmt_282/if_stmt_380__entry__
      -- 
    cp_elements(4) <= cp_elements(98);
    -- CP-element group 5 fork  transition  bypass 
    -- predecessors 111 
    -- successors 16 6 14 8 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/$entry
      -- 
    cp_elements(5) <= cp_elements(111);
    -- CP-element group 6 transition  bypass 
    -- predecessors 5 
    -- successors 7 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_trigger_
      -- 
    cp_elements(6) <= cp_elements(5);
    -- CP-element group 7 join  transition  output  bypass 
    -- predecessors 6 12 
    -- successors 13 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_complete/final_reg_req
      -- 
    cpelement_group_7 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(6);
      predecessors(1) <= cp_elements(12);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(7)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(7),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4576_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(7), ack => addr_of_298_final_reg_req_0); -- 
    -- CP-element group 8 transition  output  bypass 
    -- predecessors 5 
    -- successors 9 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_computed_0
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_296_trigger_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_296_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_296_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_resize_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_resize_0/index_resize_req
      -- 
    cp_elements(8) <= cp_elements(5);
    index_resize_req_4556_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(8), ack => array_obj_ref_297_index_0_resize_req_0); -- 
    -- CP-element group 9 transition  input  output  bypass 
    -- predecessors 8 
    -- successors 10 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_resized_0
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_resize_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_scale_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4557_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_index_0_resize_ack_0, ack => cp_elements(9)); -- 
    scale_rename_req_4561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => array_obj_ref_297_index_0_rename_req_0); -- 
    -- CP-element group 10 transition  input  output  bypass 
    -- predecessors 9 
    -- successors 11 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_indices_scaled
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_scale_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_add_indices/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_add_indices/final_index_req
      -- 
    scale_rename_ack_4562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_index_0_rename_ack_0, ack => cp_elements(10)); -- 
    final_index_req_4566_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(10), ack => array_obj_ref_297_offset_inst_req_0); -- 
    -- CP-element group 11 transition  input  output  bypass 
    -- predecessors 10 
    -- successors 12 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_offset_calculated
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_add_indices/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_add_indices/final_index_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_base_plus_offset/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4567_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_offset_inst_ack_0, ack => cp_elements(11)); -- 
    sum_rename_req_4571_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(11), ack => array_obj_ref_297_root_address_inst_req_0); -- 
    -- CP-element group 12 transition  input  bypass 
    -- predecessors 11 
    -- successors 7 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_root_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_297_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4572_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_297_root_address_inst_ack_0, ack => cp_elements(12)); -- 
    -- CP-element group 13 transition  input  bypass 
    -- predecessors 7 
    -- successors 22 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_299_trigger_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_299_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_299_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_298_complete/final_reg_ack
      -- 
    final_reg_ack_4577_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_298_final_reg_ack_0, ack => cp_elements(13)); -- 
    -- CP-element group 14 transition  bypass 
    -- predecessors 5 
    -- successors 15 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_trigger_
      -- 
    cp_elements(14) <= cp_elements(5);
    -- CP-element group 15 join  transition  output  bypass 
    -- predecessors 14 20 
    -- successors 21 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_complete/final_reg_req
      -- 
    cpelement_group_15 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(14);
      predecessors(1) <= cp_elements(20);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(15)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(15),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4615_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(15), ack => addr_of_303_final_reg_req_0); -- 
    -- CP-element group 16 transition  output  bypass 
    -- predecessors 5 
    -- successors 17 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_computed_0
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_301_trigger_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_301_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/simple_obj_ref_301_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_resize_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_resize_0/index_resize_req
      -- 
    cp_elements(16) <= cp_elements(5);
    index_resize_req_4595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(16), ack => array_obj_ref_302_index_0_resize_req_0); -- 
    -- CP-element group 17 transition  input  output  bypass 
    -- predecessors 16 
    -- successors 18 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_resized_0
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_resize_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_scale_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_scale_0/scale_rename_req
      -- 
    index_resize_ack_4596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_302_index_0_resize_ack_0, ack => cp_elements(17)); -- 
    scale_rename_req_4600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(17), ack => array_obj_ref_302_index_0_rename_req_0); -- 
    -- CP-element group 18 transition  input  output  bypass 
    -- predecessors 17 
    -- successors 19 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_indices_scaled
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_scale_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_add_indices/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_add_indices/final_index_req
      -- 
    scale_rename_ack_4601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_302_index_0_rename_ack_0, ack => cp_elements(18)); -- 
    final_index_req_4605_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(18), ack => array_obj_ref_302_offset_inst_req_0); -- 
    -- CP-element group 19 transition  input  output  bypass 
    -- predecessors 18 
    -- successors 20 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_offset_calculated
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_add_indices/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_add_indices/final_index_ack
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_base_plus_offset/$entry
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_base_plus_offset/sum_rename_req
      -- 
    final_index_ack_4606_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_302_offset_inst_ack_0, ack => cp_elements(19)); -- 
    sum_rename_req_4610_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(19), ack => array_obj_ref_302_root_address_inst_req_0); -- 
    -- CP-element group 20 transition  input  bypass 
    -- predecessors 19 
    -- successors 15 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_root_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/array_obj_ref_302_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4611_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_302_root_address_inst_ack_0, ack => cp_elements(20)); -- 
    -- CP-element group 21 transition  input  bypass 
    -- predecessors 15 
    -- successors 22 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_304_trigger_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_304_active_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/assign_stmt_304_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_completed_
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/addr_of_303_complete/final_reg_ack
      -- 
    final_reg_ack_4616_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_303_final_reg_ack_0, ack => cp_elements(21)); -- 
    -- CP-element group 22 join  transition  bypass 
    -- predecessors 21 13 
    -- successors 1 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304/$exit
      -- 
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(21);
      predecessors(1) <= cp_elements(13);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(22)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 23 transition  place  input  bypass 
    -- predecessors 1 
    -- successors 24 
    -- members (9) 
      -- 	branch_block_stmt_282/assign_stmt_307__exit__
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327__entry__
      -- 	branch_block_stmt_282/assign_stmt_307/$exit
      -- 	branch_block_stmt_282/assign_stmt_307/assign_stmt_307_trigger_
      -- 	branch_block_stmt_282/assign_stmt_307/assign_stmt_307_active_
      -- 	branch_block_stmt_282/assign_stmt_307/assign_stmt_307_completed_
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_completed_
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_307/simple_obj_ref_306_complete/ack
      -- 
    ack_4630_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_306_inst_ack_0, ack => cp_elements(23)); -- 
    -- CP-element group 24 fork  transition  bypass 
    -- predecessors 23 
    -- successors 25 27 34 36 50 47 43 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/$entry
      -- 
    cp_elements(24) <= cp_elements(23);
    -- CP-element group 25 transition  bypass 
    -- predecessors 24 
    -- successors 26 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_311_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_311_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_310_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_310_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_310_completed_
      -- 
    cp_elements(25) <= cp_elements(24);
    -- CP-element group 26 join  transition  output  bypass 
    -- predecessors 25 30 
    -- successors 31 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/split_req
      -- 
    cpelement_group_26 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(25);
      predecessors(1) <= cp_elements(30);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(26)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(26),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_4668_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(26), ack => ptr_deref_309_gather_scatter_req_0); -- 
    -- CP-element group 27 transition  output  bypass 
    -- predecessors 24 
    -- successors 28 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_308_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_308_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_308_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_addr_resize/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_addr_resize/base_resize_req
      -- 
    cp_elements(27) <= cp_elements(24);
    base_resize_req_4653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(27), ack => ptr_deref_309_base_resize_req_0); -- 
    -- CP-element group 28 transition  input  output  bypass 
    -- predecessors 27 
    -- successors 29 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_address_resized
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_addr_resize/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_plus_offset/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_base_resize_ack_0, ack => cp_elements(28)); -- 
    sum_rename_req_4658_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(28), ack => ptr_deref_309_root_address_inst_req_0); -- 
    -- CP-element group 29 transition  input  output  bypass 
    -- predecessors 28 
    -- successors 30 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_root_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_word_addrgen/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4659_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_root_address_inst_ack_0, ack => cp_elements(29)); -- 
    root_register_req_4663_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(29), ack => ptr_deref_309_addr_0_req_0); -- 
    -- CP-element group 30 transition  input  bypass 
    -- predecessors 29 
    -- successors 26 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_word_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_word_addrgen/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_word_addrgen/root_register_ack
      -- 
    root_register_ack_4664_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_addr_0_ack_0, ack => cp_elements(30)); -- 
    -- CP-element group 31 transition  input  output  bypass 
    -- predecessors 26 
    -- successors 32 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/split_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/word_access_0/rr
      -- 
    split_ack_4669_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_gather_scatter_ack_0, ack => cp_elements(31)); -- 
    rr_4676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(31), ack => ptr_deref_309_store_0_req_0); -- 
    -- CP-element group 32 transition  input  output  bypass 
    -- predecessors 31 
    -- successors 33 
    -- members (9) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/word_access_0/cr
      -- 
    ra_4677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_store_0_ack_0, ack => cp_elements(32)); -- 
    cr_4687_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => ptr_deref_309_store_0_req_1); -- 
    -- CP-element group 33 transition  input  bypass 
    -- predecessors 32 
    -- successors 56 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_311_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_309_complete/word_access/word_access_0/ca
      -- 
    ca_4688_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_309_store_0_ack_1, ack => cp_elements(33)); -- 
    -- CP-element group 34 transition  bypass 
    -- predecessors 24 
    -- successors 35 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_315_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_315_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_314_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_314_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_314_completed_
      -- 
    cp_elements(34) <= cp_elements(24);
    -- CP-element group 35 join  transition  output  bypass 
    -- predecessors 39 34 
    -- successors 40 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/split_req
      -- 
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(39);
      predecessors(1) <= cp_elements(34);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(35)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    split_req_4723_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(35), ack => ptr_deref_313_gather_scatter_req_0); -- 
    -- CP-element group 36 transition  output  bypass 
    -- predecessors 24 
    -- successors 37 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_312_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_312_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_312_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_addr_resize/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_addr_resize/base_resize_req
      -- 
    cp_elements(36) <= cp_elements(24);
    base_resize_req_4708_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(36), ack => ptr_deref_313_base_resize_req_0); -- 
    -- CP-element group 37 transition  input  output  bypass 
    -- predecessors 36 
    -- successors 38 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_address_resized
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_addr_resize/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_plus_offset/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_plus_offset/sum_rename_req
      -- 
    base_resize_ack_4709_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_base_resize_ack_0, ack => cp_elements(37)); -- 
    sum_rename_req_4713_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(37), ack => ptr_deref_313_root_address_inst_req_0); -- 
    -- CP-element group 38 transition  input  output  bypass 
    -- predecessors 37 
    -- successors 39 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_root_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_word_addrgen/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_word_addrgen/root_register_req
      -- 
    sum_rename_ack_4714_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_root_address_inst_ack_0, ack => cp_elements(38)); -- 
    root_register_req_4718_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(38), ack => ptr_deref_313_addr_0_req_0); -- 
    -- CP-element group 39 transition  input  bypass 
    -- predecessors 38 
    -- successors 35 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_word_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_word_addrgen/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_word_addrgen/root_register_ack
      -- 
    root_register_ack_4719_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_addr_0_ack_0, ack => cp_elements(39)); -- 
    -- CP-element group 40 transition  input  output  bypass 
    -- predecessors 35 
    -- successors 41 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/split_ack
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/word_access_0/rr
      -- 
    split_ack_4724_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_gather_scatter_ack_0, ack => cp_elements(40)); -- 
    rr_4731_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(40), ack => ptr_deref_313_store_0_req_0); -- 
    -- CP-element group 41 transition  input  output  bypass 
    -- predecessors 40 
    -- successors 42 
    -- members (9) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/word_access_0/cr
      -- 
    ra_4732_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_store_0_ack_0, ack => cp_elements(41)); -- 
    cr_4742_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => ptr_deref_313_store_0_req_1); -- 
    -- CP-element group 42 transition  input  bypass 
    -- predecessors 41 
    -- successors 56 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_315_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/ptr_deref_313_complete/word_access/word_access_0/ca
      -- 
    ca_4743_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_313_store_0_ack_1, ack => cp_elements(42)); -- 
    -- CP-element group 43 transition  bypass 
    -- predecessors 24 
    -- successors 56 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_active_
      -- 
    cp_elements(43) <= cp_elements(24);
    -- CP-element group 44 join  fork  transition  bypass 
    -- predecessors 49 48 
    -- successors 52 53 
    -- members (8) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_323_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_323_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_323_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_321_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_321_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_321_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_trigger_
      -- 
    cpelement_group_44 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(49);
      predecessors(1) <= cp_elements(48);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(44)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(44),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 45 transition  output  bypass 
    -- predecessors 47 
    -- successors 48 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_sample_start_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Sample/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Sample/rr
      -- 
    cp_elements(45) <= cp_elements(47);
    rr_4760_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(45), ack => binary_320_inst_req_0); -- 
    -- CP-element group 46 transition  output  bypass 
    -- predecessors 47 
    -- successors 49 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_update_start_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Update/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Update/cr
      -- 
    cp_elements(46) <= cp_elements(47);
    cr_4765_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(46), ack => binary_320_inst_req_1); -- 
    -- CP-element group 47 fork  transition  bypass 
    -- predecessors 24 
    -- successors 46 45 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_317_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_317_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/simple_obj_ref_317_completed_
      -- 
    cp_elements(47) <= cp_elements(24);
    -- CP-element group 48 transition  input  bypass 
    -- predecessors 45 
    -- successors 44 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_sample_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Sample/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Sample/ra
      -- 
    ra_4761_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_320_inst_ack_0, ack => cp_elements(48)); -- 
    -- CP-element group 49 transition  input  bypass 
    -- predecessors 46 
    -- successors 44 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_update_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Update/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_320_Update/ca
      -- 
    ca_4766_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_320_inst_ack_1, ack => cp_elements(49)); -- 
    -- CP-element group 50 transition  bypass 
    -- predecessors 24 
    -- successors 56 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_active_
      -- 
    cp_elements(50) <= cp_elements(24);
    -- CP-element group 51 join  transition  bypass 
    -- predecessors 54 55 
    -- successors 56 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_327_trigger_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_327_active_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/assign_stmt_327_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_completed_
      -- 
    cpelement_group_51 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(54);
      predecessors(1) <= cp_elements(55);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(51)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(51),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 52 transition  output  bypass 
    -- predecessors 44 
    -- successors 54 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Sample/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Sample/rr
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_sample_start_
      -- 
    cp_elements(52) <= cp_elements(44);
    rr_4783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(52), ack => binary_326_inst_req_0); -- 
    -- CP-element group 53 transition  output  bypass 
    -- predecessors 44 
    -- successors 55 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Update/cr
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Update/$entry
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_update_start_
      -- 
    cp_elements(53) <= cp_elements(44);
    cr_4788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => binary_326_inst_req_1); -- 
    -- CP-element group 54 transition  input  bypass 
    -- predecessors 52 
    -- successors 51 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Sample/ra
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Sample/$exit
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_sample_completed_
      -- 
    ra_4784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_326_inst_ack_0, ack => cp_elements(54)); -- 
    -- CP-element group 55 transition  input  bypass 
    -- predecessors 53 
    -- successors 51 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_update_completed_
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Update/ca
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/binary_326_Update/$exit
      -- 
    ca_4789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_326_inst_ack_1, ack => cp_elements(55)); -- 
    -- CP-element group 56 join  transition  bypass 
    -- predecessors 33 42 51 50 43 
    -- successors 2 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_311_to_assign_stmt_327/$exit
      -- 
    cpelement_group_56 : Block -- 
      signal predecessors: BooleanArray(4 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(33);
      predecessors(1) <= cp_elements(42);
      predecessors(2) <= cp_elements(51);
      predecessors(3) <= cp_elements(50);
      predecessors(4) <= cp_elements(43);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(56)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(56),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 57 transition  bypass 
    -- predecessors 2 
    -- successors 58 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_328_dead_link/$entry
      -- 
    cp_elements(57) <= cp_elements(2);
    -- CP-element group 58 transition  dead  bypass 
    -- predecessors 57 
    -- successors 59 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_328_dead_link/dead_transition
      -- 
    cp_elements(58) <= false;
    -- CP-element group 59 transition  place  bypass 
    -- predecessors 58 
    -- successors 112 
    -- members (4) 
      -- 	branch_block_stmt_282/if_stmt_328_dead_link/$exit
      -- 	branch_block_stmt_282/if_stmt_328__exit__
      -- 	branch_block_stmt_282/merge_stmt_334__entry__
      -- 	branch_block_stmt_282/merge_stmt_334_dead_link/$entry
      -- 
    cp_elements(59) <= cp_elements(58);
    -- CP-element group 60 transition  output  bypass 
    -- predecessors 2 
    -- successors 61 
    -- members (3) 
      -- 	branch_block_stmt_282/if_stmt_328_eval_test/$entry
      -- 	branch_block_stmt_282/if_stmt_328_eval_test/$exit
      -- 	branch_block_stmt_282/if_stmt_328_eval_test/branch_req
      -- 
    cp_elements(60) <= cp_elements(2);
    branch_req_4797_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(60), ack => if_stmt_328_branch_req_0); -- 
    -- CP-element group 61 branch  place  bypass 
    -- predecessors 60 
    -- successors 64 62 
    -- members (1) 
      -- 	branch_block_stmt_282/simple_obj_ref_329_place
      -- 
    cp_elements(61) <= cp_elements(60);
    -- CP-element group 62 transition  bypass 
    -- predecessors 61 
    -- successors 63 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_328_if_link/$entry
      -- 
    cp_elements(62) <= cp_elements(61);
    -- CP-element group 63 transition  place  input  output  bypass 
    -- predecessors 62 
    -- successors 66 
    -- members (15) 
      -- 	branch_block_stmt_282/sendResultx_xexit_getDatax_xexit
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_start/crr
      -- 	branch_block_stmt_282/if_stmt_328_if_link/$exit
      -- 	branch_block_stmt_282/if_stmt_328_if_link/if_choice_transition
      -- 	branch_block_stmt_282/call_stmt_345/$entry
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_start/$entry
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_trigger_
      -- 	branch_block_stmt_282/merge_stmt_344__exit__
      -- 	branch_block_stmt_282/call_stmt_345__entry__
      -- 	branch_block_stmt_282/sendResultx_xexit_getDatax_xexit_PhiReq/$entry
      -- 	branch_block_stmt_282/sendResultx_xexit_getDatax_xexit_PhiReq/$exit
      -- 	branch_block_stmt_282/merge_stmt_344_PhiReqMerge
      -- 	branch_block_stmt_282/merge_stmt_344_PhiAck/$entry
      -- 	branch_block_stmt_282/merge_stmt_344_PhiAck/$exit
      -- 	branch_block_stmt_282/merge_stmt_344_PhiAck/dummy
      -- 
    if_choice_transition_4802_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_328_branch_ack_1, ack => cp_elements(63)); -- 
    crr_4819_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(63), ack => call_stmt_345_call_req_0); -- 
    -- CP-element group 64 transition  bypass 
    -- predecessors 61 
    -- successors 65 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_328_else_link/$entry
      -- 
    cp_elements(64) <= cp_elements(61);
    -- CP-element group 65 transition  place  input  output  bypass 
    -- predecessors 64 
    -- successors 114 
    -- members (8) 
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge
      -- 	branch_block_stmt_282/if_stmt_328_else_link/$exit
      -- 	branch_block_stmt_282/if_stmt_328_else_link/else_choice_transition
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/$entry
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/$entry
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/$entry
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$entry
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/req
      -- 
    else_choice_transition_4806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_328_branch_ack_0, ack => cp_elements(65)); -- 
    req_5064_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(65), ack => type_cast_338_inst_req_0); -- 
    -- CP-element group 66 transition  input  output  bypass 
    -- predecessors 63 
    -- successors 67 
    -- members (5) 
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_complete/ccr
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_start/cra
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_complete/$entry
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_start/$exit
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_active_
      -- 
    cra_4820_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_345_call_ack_0, ack => cp_elements(66)); -- 
    ccr_4824_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(66), ack => call_stmt_345_call_req_1); -- 
    -- CP-element group 67 transition  place  input  output  bypass 
    -- predecessors 66 
    -- successors 119 
    -- members (18) 
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_complete/$exit
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_complete/cca
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_call_complete
      -- 	branch_block_stmt_282/call_stmt_345/call_stmt_345_completed_
      -- 	branch_block_stmt_282/call_stmt_345/$exit
      -- 	branch_block_stmt_282/call_stmt_345__exit__
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/$entry
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/$exit
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/$entry
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/$exit
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/$entry
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/$exit
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/req
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/ack
      -- 	branch_block_stmt_282/getDatax_xexit_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_req
      -- 
    cca_4825_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_345_call_ack_1, ack => cp_elements(67)); -- 
    phi_stmt_348_req_5124_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(67), ack => phi_stmt_348_req_0); -- 
    -- CP-element group 68 fork  transition  bypass 
    -- predecessors 121 
    -- successors 69 71 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/$entry
      -- 
    cp_elements(68) <= cp_elements(121);
    -- CP-element group 69 transition  bypass 
    -- predecessors 68 
    -- successors 70 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_trigger_
      -- 
    cp_elements(69) <= cp_elements(68);
    -- CP-element group 70 join  transition  output  bypass 
    -- predecessors 69 75 
    -- successors 76 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_complete/final_reg_req
      -- 
    cpelement_group_70 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(69);
      predecessors(1) <= cp_elements(75);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(70)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(70),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    final_reg_req_4866_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(70), ack => addr_of_359_final_reg_req_0); -- 
    -- CP-element group 71 transition  output  bypass 
    -- predecessors 68 
    -- successors 72 
    -- members (6) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_resize_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_357_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_resize_0/index_resize_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_357_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_computed_0
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_357_trigger_
      -- 
    cp_elements(71) <= cp_elements(68);
    index_resize_req_4846_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_358_index_0_resize_req_0); -- 
    -- CP-element group 72 transition  input  output  bypass 
    -- predecessors 71 
    -- successors 73 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_resize_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_scale_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_resized_0
      -- 
    index_resize_ack_4847_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_358_index_0_resize_ack_0, ack => cp_elements(72)); -- 
    scale_rename_req_4851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(72), ack => array_obj_ref_358_index_0_rename_req_0); -- 
    -- CP-element group 73 transition  input  output  bypass 
    -- predecessors 72 
    -- successors 74 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_scale_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_add_indices/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_add_indices/final_index_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_indices_scaled
      -- 
    scale_rename_ack_4852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_358_index_0_rename_ack_0, ack => cp_elements(73)); -- 
    final_index_req_4856_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_358_offset_inst_req_0); -- 
    -- CP-element group 74 transition  input  output  bypass 
    -- predecessors 73 
    -- successors 75 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_base_plus_offset/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_add_indices/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_add_indices/final_index_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_offset_calculated
      -- 
    final_index_ack_4857_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_358_offset_inst_ack_0, ack => cp_elements(74)); -- 
    sum_rename_req_4861_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(74), ack => array_obj_ref_358_root_address_inst_req_0); -- 
    -- CP-element group 75 transition  input  bypass 
    -- predecessors 74 
    -- successors 70 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/array_obj_ref_358_root_address_calculated
      -- 
    sum_rename_ack_4862_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_358_root_address_inst_ack_0, ack => cp_elements(75)); -- 
    -- CP-element group 76 transition  input  output  bypass 
    -- predecessors 70 
    -- successors 77 
    -- members (12) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_360_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_360_trigger_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_addr_resize/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_360_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_362_trigger_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_362_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/simple_obj_ref_362_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/addr_of_359_complete/final_reg_ack
      -- 
    final_reg_ack_4867_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_359_final_reg_ack_0, ack => cp_elements(76)); -- 
    base_resize_req_4884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(76), ack => ptr_deref_363_base_resize_req_0); -- 
    -- CP-element group 77 transition  input  output  bypass 
    -- predecessors 76 
    -- successors 78 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_addr_resize/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_address_resized
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_plus_offset/$entry
      -- 
    base_resize_ack_4885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_base_resize_ack_0, ack => cp_elements(77)); -- 
    sum_rename_req_4889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => ptr_deref_363_root_address_inst_req_0); -- 
    -- CP-element group 78 transition  input  output  bypass 
    -- predecessors 77 
    -- successors 79 
    -- members (5) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_root_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_plus_offset/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_word_addrgen/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_word_addrgen/root_register_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_root_address_inst_ack_0, ack => cp_elements(78)); -- 
    root_register_req_4894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(78), ack => ptr_deref_363_addr_0_req_0); -- 
    -- CP-element group 79 transition  input  output  bypass 
    -- predecessors 78 
    -- successors 80 
    -- members (8) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_word_address_calculated
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_trigger_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_word_addrgen/root_register_ack
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_word_addrgen/$exit
      -- 
    root_register_ack_4895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_addr_0_ack_0, ack => cp_elements(79)); -- 
    rr_4905_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => ptr_deref_363_load_0_req_0); -- 
    -- CP-element group 80 transition  input  output  bypass 
    -- predecessors 79 
    -- successors 81 
    -- members (9) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_request/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/word_access_0/$entry
      -- 
    ra_4906_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_load_0_ack_0, ack => cp_elements(80)); -- 
    cr_4916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(80), ack => ptr_deref_363_load_0_req_1); -- 
    -- CP-element group 81 transition  input  output  bypass 
    -- predecessors 80 
    -- successors 82 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/merge_req
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/word_access/word_access_0/$exit
      -- 
    ca_4917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_load_0_ack_1, ack => cp_elements(81)); -- 
    merge_req_4918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(81), ack => ptr_deref_363_gather_scatter_req_0); -- 
    -- CP-element group 82 transition  place  input  output  bypass 
    -- predecessors 81 
    -- successors 83 
    -- members (18) 
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/$exit
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_364_trigger_
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_complete/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/merge_ack
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_366_trigger_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_364_active_
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_complete/pipe_wreq
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_trigger_
      -- 	branch_block_stmt_282/assign_stmt_367/$entry
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/ptr_deref_363_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_366_active_
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_366_completed_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364/assign_stmt_364_completed_
      -- 	branch_block_stmt_282/assign_stmt_367/assign_stmt_367_trigger_
      -- 	branch_block_stmt_282/assign_stmt_367/assign_stmt_367_active_
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364__exit__
      -- 	branch_block_stmt_282/assign_stmt_367__entry__
      -- 
    merge_ack_4919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_363_gather_scatter_ack_0, ack => cp_elements(82)); -- 
    pipe_wreq_4935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(82), ack => simple_obj_ref_365_inst_req_0); -- 
    -- CP-element group 83 transition  place  input  bypass 
    -- predecessors 82 
    -- successors 84 
    -- members (8) 
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_complete/$exit
      -- 	branch_block_stmt_282/assign_stmt_367/assign_stmt_367_completed_
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_complete/pipe_wack
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_active_
      -- 	branch_block_stmt_282/assign_stmt_367/simple_obj_ref_365_completed_
      -- 	branch_block_stmt_282/assign_stmt_367/$exit
      -- 	branch_block_stmt_282/assign_stmt_367__exit__
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379__entry__
      -- 
    pipe_wack_4936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_365_inst_ack_0, ack => cp_elements(83)); -- 
    -- CP-element group 84 fork  transition  bypass 
    -- predecessors 83 
    -- successors 85 89 92 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/$entry
      -- 
    cp_elements(84) <= cp_elements(83);
    -- CP-element group 85 transition  bypass 
    -- predecessors 84 
    -- successors 98 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_active_
      -- 
    cp_elements(85) <= cp_elements(84);
    -- CP-element group 86 join  fork  transition  bypass 
    -- predecessors 90 91 
    -- successors 94 95 
    -- members (8) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_373_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_375_active_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_375_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_373_trigger_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_373_active_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_375_trigger_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_trigger_
      -- 
    cpelement_group_86 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(90);
      predecessors(1) <= cp_elements(91);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(86)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(86),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 87 transition  output  bypass 
    -- predecessors 89 
    -- successors 90 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Sample/rr
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_sample_start_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Sample/$entry
      -- 
    cp_elements(87) <= cp_elements(89);
    rr_4956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(87), ack => binary_372_inst_req_0); -- 
    -- CP-element group 88 transition  output  bypass 
    -- predecessors 89 
    -- successors 91 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_update_start_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Update/$entry
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Update/cr
      -- 
    cp_elements(88) <= cp_elements(89);
    cr_4961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(88), ack => binary_372_inst_req_1); -- 
    -- CP-element group 89 fork  transition  bypass 
    -- predecessors 84 
    -- successors 87 88 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_trigger_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_369_active_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_369_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/simple_obj_ref_369_trigger_
      -- 
    cp_elements(89) <= cp_elements(84);
    -- CP-element group 90 transition  input  bypass 
    -- predecessors 87 
    -- successors 86 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Sample/$exit
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_sample_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Sample/ra
      -- 
    ra_4957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_372_inst_ack_0, ack => cp_elements(90)); -- 
    -- CP-element group 91 transition  input  bypass 
    -- predecessors 88 
    -- successors 86 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Update/ca
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_update_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_372_Update/$exit
      -- 
    ca_4962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_372_inst_ack_1, ack => cp_elements(91)); -- 
    -- CP-element group 92 transition  bypass 
    -- predecessors 84 
    -- successors 98 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_active_
      -- 
    cp_elements(92) <= cp_elements(84);
    -- CP-element group 93 join  transition  bypass 
    -- predecessors 96 97 
    -- successors 98 
    -- members (4) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_379_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_379_trigger_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/assign_stmt_379_active_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_completed_
      -- 
    cpelement_group_93 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(96);
      predecessors(1) <= cp_elements(97);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(93)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(93),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 94 transition  output  bypass 
    -- predecessors 86 
    -- successors 96 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_sample_start_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Sample/$entry
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Sample/rr
      -- 
    cp_elements(94) <= cp_elements(86);
    rr_4979_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(94), ack => binary_378_inst_req_0); -- 
    -- CP-element group 95 transition  output  bypass 
    -- predecessors 86 
    -- successors 97 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_update_start_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Update/$entry
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Update/cr
      -- 
    cp_elements(95) <= cp_elements(86);
    cr_4984_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => binary_378_inst_req_1); -- 
    -- CP-element group 96 transition  input  bypass 
    -- predecessors 94 
    -- successors 93 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_sample_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Sample/$exit
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Sample/ra
      -- 
    ra_4980_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_378_inst_ack_0, ack => cp_elements(96)); -- 
    -- CP-element group 97 transition  input  bypass 
    -- predecessors 95 
    -- successors 93 
    -- members (3) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_update_completed_
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Update/$exit
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/binary_378_Update/ca
      -- 
    ca_4985_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_378_inst_ack_1, ack => cp_elements(97)); -- 
    -- CP-element group 98 join  transition  bypass 
    -- predecessors 85 92 93 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_282/assign_stmt_373_to_assign_stmt_379/$exit
      -- 
    cpelement_group_98 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(85);
      predecessors(1) <= cp_elements(92);
      predecessors(2) <= cp_elements(93);
      jNoI: join -- 
        generic map(place_capacity => 1,
        bypass => true,
        name => " cp_elements(98)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(98),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 99 transition  bypass 
    -- predecessors 4 
    -- successors 100 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_380_dead_link/$entry
      -- 
    cp_elements(99) <= cp_elements(4);
    -- CP-element group 100 transition  dead  bypass 
    -- predecessors 99 
    -- successors 101 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_380_dead_link/dead_transition
      -- 
    cp_elements(100) <= false;
    -- CP-element group 101 transition  place  bypass 
    -- predecessors 100 
    -- successors 
    -- members (5) 
      -- 	$exit
      -- 	branch_block_stmt_282/$exit
      -- 	branch_block_stmt_282/branch_block_stmt_282__exit__
      -- 	branch_block_stmt_282/if_stmt_380__exit__
      -- 	branch_block_stmt_282/if_stmt_380_dead_link/$exit
      -- 
    cp_elements(101) <= cp_elements(100);
    -- CP-element group 102 transition  output  bypass 
    -- predecessors 4 
    -- successors 103 
    -- members (3) 
      -- 	branch_block_stmt_282/if_stmt_380_eval_test/$entry
      -- 	branch_block_stmt_282/if_stmt_380_eval_test/$exit
      -- 	branch_block_stmt_282/if_stmt_380_eval_test/branch_req
      -- 
    cp_elements(102) <= cp_elements(4);
    branch_req_4993_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(102), ack => if_stmt_380_branch_req_0); -- 
    -- CP-element group 103 branch  place  bypass 
    -- predecessors 102 
    -- successors 104 106 
    -- members (1) 
      -- 	branch_block_stmt_282/simple_obj_ref_381_place
      -- 
    cp_elements(103) <= cp_elements(102);
    -- CP-element group 104 transition  bypass 
    -- predecessors 103 
    -- successors 105 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_380_if_link/$entry
      -- 
    cp_elements(104) <= cp_elements(103);
    -- CP-element group 105 transition  place  input  output  bypass 
    -- predecessors 104 
    -- successors 115 
    -- members (22) 
      -- 	branch_block_stmt_282/merge_stmt_284__exit__
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge
      -- 	branch_block_stmt_282/if_stmt_380_if_link/$exit
      -- 	branch_block_stmt_282/if_stmt_380_if_link/if_choice_transition
      -- 	branch_block_stmt_282/bb_5_sendResultx_xexitx_xloopexit
      -- 	branch_block_stmt_282/bb_5_sendResultx_xexitx_xloopexit_PhiReq/$entry
      -- 	branch_block_stmt_282/bb_5_sendResultx_xexitx_xloopexit_PhiReq/$exit
      -- 	branch_block_stmt_282/merge_stmt_284_PhiReqMerge
      -- 	branch_block_stmt_282/merge_stmt_284_PhiAck/$entry
      -- 	branch_block_stmt_282/merge_stmt_284_PhiAck/$exit
      -- 	branch_block_stmt_282/merge_stmt_284_PhiAck/dummy
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$entry
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/req
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/ack
      -- 	branch_block_stmt_282/sendResultx_xexitx_xloopexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_req
      -- 
    if_choice_transition_4998_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_380_branch_ack_1, ack => cp_elements(105)); -- 
    phi_stmt_335_req_5081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(105), ack => phi_stmt_335_req_1); -- 
    -- CP-element group 106 transition  bypass 
    -- predecessors 103 
    -- successors 107 
    -- members (1) 
      -- 	branch_block_stmt_282/if_stmt_380_else_link/$entry
      -- 
    cp_elements(106) <= cp_elements(103);
    -- CP-element group 107 transition  place  input  output  bypass 
    -- predecessors 106 
    -- successors 118 
    -- members (8) 
      -- 	branch_block_stmt_282/if_stmt_380_else_link/$exit
      -- 	branch_block_stmt_282/if_stmt_380_else_link/else_choice_transition
      -- 	branch_block_stmt_282/bb_5_bb_5
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/$entry
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/$entry
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/$entry
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/$entry
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/req
      -- 
    else_choice_transition_5002_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_380_branch_ack_0, ack => cp_elements(107)); -- 
    req_5107_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(107), ack => type_cast_354_inst_req_0); -- 
    -- CP-element group 108 transition  input  output  bypass 
    -- predecessors 3 
    -- successors 109 
    -- members (6) 
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/$exit
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_sources/type_cast_293/ack
      -- 	branch_block_stmt_282/sendResultx_xexitx_xbackedge_sendResultx_xexit_PhiReq/phi_stmt_287/phi_stmt_287_req
      -- 
    ack_5041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_293_inst_ack_0, ack => cp_elements(108)); -- 
    phi_stmt_287_req_5042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => phi_stmt_287_req_1); -- 
    -- CP-element group 109 merge  place  bypass 
    -- predecessors 108 0 
    -- successors 110 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_286_PhiReqMerge
      -- 
    cp_elements(109) <= OrReduce(cp_elements(108) & cp_elements(0));
    -- CP-element group 110 transition  bypass 
    -- predecessors 109 
    -- successors 111 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_286_PhiAck/$entry
      -- 
    cp_elements(110) <= cp_elements(109);
    -- CP-element group 111 transition  place  input  bypass 
    -- predecessors 110 
    -- successors 5 
    -- members (4) 
      -- 	branch_block_stmt_282/merge_stmt_286__exit__
      -- 	branch_block_stmt_282/assign_stmt_299_to_assign_stmt_304__entry__
      -- 	branch_block_stmt_282/merge_stmt_286_PhiAck/$exit
      -- 	branch_block_stmt_282/merge_stmt_286_PhiAck/phi_stmt_287_ack
      -- 
    phi_stmt_287_ack_5047_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_287_ack_0, ack => cp_elements(111)); -- 
    -- CP-element group 112 transition  dead  bypass 
    -- predecessors 59 
    -- successors 113 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_334_dead_link/dead_transition
      -- 
    cp_elements(112) <= false;
    -- CP-element group 113 transition  bypass 
    -- predecessors 112 
    -- successors 3 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_334_dead_link/$exit
      -- 
    cp_elements(113) <= cp_elements(112);
    -- CP-element group 114 transition  input  output  bypass 
    -- predecessors 65 
    -- successors 115 
    -- members (6) 
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/$exit
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/$exit
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/$exit
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/$exit
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_sources/type_cast_338/ack
      -- 	branch_block_stmt_282/sendResultx_xexit_sendResultx_xexitx_xbackedge_PhiReq/phi_stmt_335/phi_stmt_335_req
      -- 
    ack_5065_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_338_inst_ack_0, ack => cp_elements(114)); -- 
    phi_stmt_335_req_5066_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(114), ack => phi_stmt_335_req_0); -- 
    -- CP-element group 115 merge  place  bypass 
    -- predecessors 105 114 
    -- successors 116 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_334_PhiReqMerge
      -- 
    cp_elements(115) <= OrReduce(cp_elements(105) & cp_elements(114));
    -- CP-element group 116 transition  bypass 
    -- predecessors 115 
    -- successors 117 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_334_PhiAck/$entry
      -- 
    cp_elements(116) <= cp_elements(115);
    -- CP-element group 117 transition  input  bypass 
    -- predecessors 116 
    -- successors 3 
    -- members (2) 
      -- 	branch_block_stmt_282/merge_stmt_334_PhiAck/$exit
      -- 	branch_block_stmt_282/merge_stmt_334_PhiAck/phi_stmt_335_ack
      -- 
    phi_stmt_335_ack_5086_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_335_ack_0, ack => cp_elements(117)); -- 
    -- CP-element group 118 transition  input  output  bypass 
    -- predecessors 107 
    -- successors 119 
    -- members (6) 
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/$exit
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/$exit
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/$exit
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/$exit
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_sources/type_cast_354/ack
      -- 	branch_block_stmt_282/bb_5_bb_5_PhiReq/phi_stmt_348/phi_stmt_348_req
      -- 
    ack_5108_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_354_inst_ack_0, ack => cp_elements(118)); -- 
    phi_stmt_348_req_5109_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => phi_stmt_348_req_1); -- 
    -- CP-element group 119 merge  place  bypass 
    -- predecessors 118 67 
    -- successors 120 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_347_PhiReqMerge
      -- 
    cp_elements(119) <= OrReduce(cp_elements(118) & cp_elements(67));
    -- CP-element group 120 transition  bypass 
    -- predecessors 119 
    -- successors 121 
    -- members (1) 
      -- 	branch_block_stmt_282/merge_stmt_347_PhiAck/$entry
      -- 
    cp_elements(120) <= cp_elements(119);
    -- CP-element group 121 transition  place  input  bypass 
    -- predecessors 120 
    -- successors 68 
    -- members (4) 
      -- 	branch_block_stmt_282/merge_stmt_347__exit__
      -- 	branch_block_stmt_282/assign_stmt_360_to_assign_stmt_364__entry__
      -- 	branch_block_stmt_282/merge_stmt_347_PhiAck/$exit
      -- 	branch_block_stmt_282/merge_stmt_347_PhiAck/phi_stmt_348_ack
      -- 
    phi_stmt_348_ack_5129_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_348_ack_0, ack => cp_elements(121)); -- 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_297_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_297_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_297_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_297_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_302_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_302_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_302_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_302_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_358_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_358_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_358_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_358_root_address : std_logic_vector(6 downto 0);
    signal exitcond1_379 : std_logic_vector(0 downto 0);
    signal exitcondx_xi_327 : std_logic_vector(0 downto 0);
    signal iNsTr_10_364 : std_logic_vector(31 downto 0);
    signal iNsTr_13_373 : std_logic_vector(31 downto 0);
    signal iNsTr_2_307 : std_logic_vector(31 downto 0);
    signal iNsTr_5_321 : std_logic_vector(31 downto 0);
    signal idxx_x01x_xi1_348 : std_logic_vector(31 downto 0);
    signal idxx_x01x_xi_287 : std_logic_vector(31 downto 0);
    signal idxx_x01x_xix_xbe_335 : std_logic_vector(31 downto 0);
    signal ptr_deref_309_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_309_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_309_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_309_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_309_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_309_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_313_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_313_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_313_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_313_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_313_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_313_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_363_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_363_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_363_word_offset_0 : std_logic_vector(6 downto 0);
    signal scevgep2x_xi_304 : std_logic_vector(31 downto 0);
    signal scevgepx_xi2_360 : std_logic_vector(31 downto 0);
    signal scevgepx_xi_299 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_296_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_296_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_301_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_301_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_357_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_357_scaled : std_logic_vector(6 downto 0);
    signal type_cast_291_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_293_wire : std_logic_vector(31 downto 0);
    signal type_cast_319_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_325_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_338_wire : std_logic_vector(31 downto 0);
    signal type_cast_341_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_352_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_354_wire : std_logic_vector(31 downto 0);
    signal type_cast_371_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_377_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_297_offset_scale_factor_0 <= "0000001";
    array_obj_ref_297_resized_base_address <= "0000000";
    array_obj_ref_302_offset_scale_factor_0 <= "0000001";
    array_obj_ref_302_resized_base_address <= "0000000";
    array_obj_ref_358_offset_scale_factor_0 <= "0000001";
    array_obj_ref_358_resized_base_address <= "0000000";
    ptr_deref_309_word_offset_0 <= "0000000";
    ptr_deref_313_word_offset_0 <= "0000000";
    ptr_deref_363_word_offset_0 <= "0000000";
    type_cast_291_wire_constant <= "00000000000000000000000000000000";
    type_cast_319_wire_constant <= "00000000000000000000000000000001";
    type_cast_325_wire_constant <= "00000000000000000000000001000000";
    type_cast_341_wire_constant <= "00000000000000000000000000000000";
    type_cast_352_wire_constant <= "00000000000000000000000000000000";
    type_cast_371_wire_constant <= "00000000000000000000000000000001";
    type_cast_377_wire_constant <= "00000000000000000000000001000000";
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_287_req_0," req0 phi_stmt_287");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_287_req_1," req1 phi_stmt_287");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_287_ack_0," ack0 phi_stmt_287");
    phi_stmt_287: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_291_wire_constant & type_cast_293_wire;
      req <= phi_stmt_287_req_0 & phi_stmt_287_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_287_ack_0,
          idata => idata,
          odata => idxx_x01x_xi_287,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_287
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_335_req_0," req0 phi_stmt_335");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_335_req_1," req1 phi_stmt_335");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_335_ack_0," ack0 phi_stmt_335");
    phi_stmt_335: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_338_wire & type_cast_341_wire_constant;
      req <= phi_stmt_335_req_0 & phi_stmt_335_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_335_ack_0,
          idata => idata,
          odata => idxx_x01x_xix_xbe_335,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_335
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_348_req_0," req0 phi_stmt_348");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_348_req_1," req1 phi_stmt_348");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_348_ack_0," ack0 phi_stmt_348");
    phi_stmt_348: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_352_wire_constant & type_cast_354_wire;
      req <= phi_stmt_348_req_0 & phi_stmt_348_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_348_ack_0,
          idata => idata,
          odata => idxx_x01x_xi1_348,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_348
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_298_final_reg_req_0,addr_of_298_final_reg_ack_0,sl_one,"addr_of_298_final_reg ",false,array_obj_ref_297_root_address,
    false,scevgepx_xi_299);
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_298_final_reg_req_0;
      addr_of_298_final_reg_ack_0 <= ack; 
      addr_of_298_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_297_root_address, dout => scevgepx_xi_299, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_303_final_reg_req_0,addr_of_303_final_reg_ack_0,sl_one,"addr_of_303_final_reg ",false,array_obj_ref_302_root_address,
    false,scevgep2x_xi_304);
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_303_final_reg_req_0;
      addr_of_303_final_reg_ack_0 <= ack; 
      addr_of_303_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_302_root_address, dout => scevgep2x_xi_304, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_359_final_reg_req_0,addr_of_359_final_reg_ack_0,sl_one,"addr_of_359_final_reg ",false,array_obj_ref_358_root_address,
    false,scevgepx_xi2_360);
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_359_final_reg_req_0;
      addr_of_359_final_reg_ack_0 <= ack; 
      addr_of_359_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_358_root_address, dout => scevgepx_xi2_360, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_293_inst_req_0,type_cast_293_inst_ack_0,sl_one,"type_cast_293_inst ",false,idxx_x01x_xix_xbe_335,
    false,type_cast_293_wire);
    register_block_3 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_293_inst_req_0;
      type_cast_293_inst_ack_0 <= ack; 
      type_cast_293_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => idxx_x01x_xix_xbe_335, dout => type_cast_293_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_338_inst_req_0,type_cast_338_inst_ack_0,sl_one,"type_cast_338_inst ",false,iNsTr_5_321,
    false,type_cast_338_wire);
    register_block_4 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_338_inst_req_0;
      type_cast_338_inst_ack_0 <= ack; 
      type_cast_338_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_5_321, dout => type_cast_338_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_354_inst_req_0,type_cast_354_inst_ack_0,sl_one,"type_cast_354_inst ",false,iNsTr_13_373,
    false,type_cast_354_wire);
    register_block_5 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_354_inst_req_0;
      type_cast_354_inst_ack_0 <= ack; 
      type_cast_354_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => iNsTr_13_373, dout => type_cast_354_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_297_index_0_rename_req_0,array_obj_ref_297_index_0_rename_ack_0,sl_one,"array_obj_ref_297_index_0_rename ",false,simple_obj_ref_296_resized,
    false,simple_obj_ref_296_scaled);
    array_obj_ref_297_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_297_index_0_rename_ack_0 <= array_obj_ref_297_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_296_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_296_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_297_index_0_resize_req_0,array_obj_ref_297_index_0_resize_ack_0,sl_one,"array_obj_ref_297_index_0_resize ",false,idxx_x01x_xi_287,
    false,simple_obj_ref_296_resized);
    array_obj_ref_297_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_297_index_0_resize_ack_0 <= array_obj_ref_297_index_0_resize_req_0;
      in_aggregated_sig <= idxx_x01x_xi_287;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_296_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_297_offset_inst_req_0,array_obj_ref_297_offset_inst_ack_0,sl_one,"array_obj_ref_297_offset_inst ",false,simple_obj_ref_296_scaled,
    false,array_obj_ref_297_final_offset);
    array_obj_ref_297_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_297_offset_inst_ack_0 <= array_obj_ref_297_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_296_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_297_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_297_root_address_inst_req_0,array_obj_ref_297_root_address_inst_ack_0,sl_one,"array_obj_ref_297_root_address_inst ",false,array_obj_ref_297_final_offset,
    false,array_obj_ref_297_root_address);
    array_obj_ref_297_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_297_root_address_inst_ack_0 <= array_obj_ref_297_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_297_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_297_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_302_index_0_rename_req_0,array_obj_ref_302_index_0_rename_ack_0,sl_one,"array_obj_ref_302_index_0_rename ",false,simple_obj_ref_301_resized,
    false,simple_obj_ref_301_scaled);
    array_obj_ref_302_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_302_index_0_rename_ack_0 <= array_obj_ref_302_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_301_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_301_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_302_index_0_resize_req_0,array_obj_ref_302_index_0_resize_ack_0,sl_one,"array_obj_ref_302_index_0_resize ",false,idxx_x01x_xi_287,
    false,simple_obj_ref_301_resized);
    array_obj_ref_302_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_302_index_0_resize_ack_0 <= array_obj_ref_302_index_0_resize_req_0;
      in_aggregated_sig <= idxx_x01x_xi_287;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_301_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_302_offset_inst_req_0,array_obj_ref_302_offset_inst_ack_0,sl_one,"array_obj_ref_302_offset_inst ",false,simple_obj_ref_301_scaled,
    false,array_obj_ref_302_final_offset);
    array_obj_ref_302_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_302_offset_inst_ack_0 <= array_obj_ref_302_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_301_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_302_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_302_root_address_inst_req_0,array_obj_ref_302_root_address_inst_ack_0,sl_one,"array_obj_ref_302_root_address_inst ",false,array_obj_ref_302_final_offset,
    false,array_obj_ref_302_root_address);
    array_obj_ref_302_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_302_root_address_inst_ack_0 <= array_obj_ref_302_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_302_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_302_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_358_index_0_rename_req_0,array_obj_ref_358_index_0_rename_ack_0,sl_one,"array_obj_ref_358_index_0_rename ",false,simple_obj_ref_357_resized,
    false,simple_obj_ref_357_scaled);
    array_obj_ref_358_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_358_index_0_rename_ack_0 <= array_obj_ref_358_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_357_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_357_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_358_index_0_resize_req_0,array_obj_ref_358_index_0_resize_ack_0,sl_one,"array_obj_ref_358_index_0_resize ",false,idxx_x01x_xi1_348,
    false,simple_obj_ref_357_resized);
    array_obj_ref_358_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_358_index_0_resize_ack_0 <= array_obj_ref_358_index_0_resize_req_0;
      in_aggregated_sig <= idxx_x01x_xi1_348;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_357_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_358_offset_inst_req_0,array_obj_ref_358_offset_inst_ack_0,sl_one,"array_obj_ref_358_offset_inst ",false,simple_obj_ref_357_scaled,
    false,array_obj_ref_358_final_offset);
    array_obj_ref_358_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_358_offset_inst_ack_0 <= array_obj_ref_358_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_357_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_358_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_358_root_address_inst_req_0,array_obj_ref_358_root_address_inst_ack_0,sl_one,"array_obj_ref_358_root_address_inst ",false,array_obj_ref_358_final_offset,
    false,array_obj_ref_358_root_address);
    array_obj_ref_358_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_358_root_address_inst_ack_0 <= array_obj_ref_358_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_358_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_358_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_309_addr_0_req_0,ptr_deref_309_addr_0_ack_0,sl_one,"ptr_deref_309_addr_0 ",false,ptr_deref_309_root_address,
    false,ptr_deref_309_word_address_0);
    ptr_deref_309_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_309_addr_0_ack_0 <= ptr_deref_309_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_309_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_309_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_309_base_resize_req_0,ptr_deref_309_base_resize_ack_0,sl_one,"ptr_deref_309_base_resize ",false,scevgepx_xi_299,
    false,ptr_deref_309_resized_base_address);
    ptr_deref_309_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_309_base_resize_ack_0 <= ptr_deref_309_base_resize_req_0;
      in_aggregated_sig <= scevgepx_xi_299;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_309_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_309_gather_scatter_req_0,ptr_deref_309_gather_scatter_ack_0,sl_one,"ptr_deref_309_gather_scatter ",false,iNsTr_2_307,
    false,ptr_deref_309_data_0);
    ptr_deref_309_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_309_gather_scatter_ack_0 <= ptr_deref_309_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_2_307;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_309_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_309_root_address_inst_req_0,ptr_deref_309_root_address_inst_ack_0,sl_one,"ptr_deref_309_root_address_inst ",false,ptr_deref_309_resized_base_address,
    false,ptr_deref_309_root_address);
    ptr_deref_309_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_309_root_address_inst_ack_0 <= ptr_deref_309_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_309_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_309_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_313_addr_0_req_0,ptr_deref_313_addr_0_ack_0,sl_one,"ptr_deref_313_addr_0 ",false,ptr_deref_313_root_address,
    false,ptr_deref_313_word_address_0);
    ptr_deref_313_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_313_addr_0_ack_0 <= ptr_deref_313_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_313_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_313_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_313_base_resize_req_0,ptr_deref_313_base_resize_ack_0,sl_one,"ptr_deref_313_base_resize ",false,scevgep2x_xi_304,
    false,ptr_deref_313_resized_base_address);
    ptr_deref_313_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_313_base_resize_ack_0 <= ptr_deref_313_base_resize_req_0;
      in_aggregated_sig <= scevgep2x_xi_304;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_313_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_313_gather_scatter_req_0,ptr_deref_313_gather_scatter_ack_0,sl_one,"ptr_deref_313_gather_scatter ",false,iNsTr_2_307,
    false,ptr_deref_313_data_0);
    ptr_deref_313_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_313_gather_scatter_ack_0 <= ptr_deref_313_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_2_307;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_313_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_313_root_address_inst_req_0,ptr_deref_313_root_address_inst_ack_0,sl_one,"ptr_deref_313_root_address_inst ",false,ptr_deref_313_resized_base_address,
    false,ptr_deref_313_root_address);
    ptr_deref_313_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_313_root_address_inst_ack_0 <= ptr_deref_313_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_313_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_313_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_363_addr_0_req_0,ptr_deref_363_addr_0_ack_0,sl_one,"ptr_deref_363_addr_0 ",false,ptr_deref_363_root_address,
    false,ptr_deref_363_word_address_0);
    ptr_deref_363_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_363_addr_0_ack_0 <= ptr_deref_363_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_363_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_363_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_363_base_resize_req_0,ptr_deref_363_base_resize_ack_0,sl_one,"ptr_deref_363_base_resize ",false,scevgepx_xi2_360,
    false,ptr_deref_363_resized_base_address);
    ptr_deref_363_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_363_base_resize_ack_0 <= ptr_deref_363_base_resize_req_0;
      in_aggregated_sig <= scevgepx_xi2_360;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_363_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_363_gather_scatter_req_0,ptr_deref_363_gather_scatter_ack_0,sl_one,"ptr_deref_363_gather_scatter ",false,ptr_deref_363_data_0,
    false,iNsTr_10_364);
    ptr_deref_363_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_363_gather_scatter_ack_0 <= ptr_deref_363_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_363_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_10_364 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_363_root_address_inst_req_0,ptr_deref_363_root_address_inst_ack_0,sl_one,"ptr_deref_363_root_address_inst ",false,ptr_deref_363_resized_base_address,
    false,ptr_deref_363_root_address);
    ptr_deref_363_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_363_root_address_inst_ack_0 <= ptr_deref_363_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_363_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_363_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_328_branch_req_0," req0 if_stmt_328_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_328_branch_ack_0," ack0 if_stmt_328_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_328_branch_ack_1," ack1 if_stmt_328_branch");
    if_stmt_328_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcondx_xi_327;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_328_branch_req_0,
          ack0 => if_stmt_328_branch_ack_0,
          ack1 => if_stmt_328_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_380_branch_req_0," req0 if_stmt_380_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_380_branch_ack_0," ack0 if_stmt_380_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,if_stmt_380_branch_ack_1," ack1 if_stmt_380_branch");
    if_stmt_380_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= exitcond1_379;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_380_branch_req_0,
          ack0 => if_stmt_380_branch_ack_0,
          ack1 => if_stmt_380_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_320_inst_req_0,binary_320_inst_ack_0,binary_320_inst_req_1,binary_320_inst_ack_1,sl_one,"binary_320_inst",false,idxx_x01x_xi_287 & type_cast_319_wire_constant,
    false,iNsTr_5_321);
    -- shared split operator group (0) : binary_320_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= idxx_x01x_xi_287;
      iNsTr_5_321 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_320_inst_req_0;
      reqR(0) <= binary_320_inst_req_1;
      binary_320_inst_ack_0 <= ackL(0); 
      binary_320_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_326_inst_req_0,binary_326_inst_ack_0,binary_326_inst_req_1,binary_326_inst_ack_1,sl_one,"binary_326_inst",false,iNsTr_5_321 & type_cast_325_wire_constant,
    false,exitcondx_xi_327);
    -- shared split operator group (1) : binary_326_inst 
    ApIntEq_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_5_321;
      exitcondx_xi_327 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_326_inst_req_0;
      reqR(0) <= binary_326_inst_req_1;
      binary_326_inst_ack_0 <= ackL(0); 
      binary_326_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_372_inst_req_0,binary_372_inst_ack_0,binary_372_inst_req_1,binary_372_inst_ack_1,sl_one,"binary_372_inst",false,idxx_x01x_xi1_348 & type_cast_371_wire_constant,
    false,iNsTr_13_373);
    -- shared split operator group (2) : binary_372_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= idxx_x01x_xi1_348;
      iNsTr_13_373 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_372_inst_req_0;
      reqR(0) <= binary_372_inst_req_1;
      binary_372_inst_ack_0 <= ackL(0); 
      binary_372_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_378_inst_req_0,binary_378_inst_ack_0,binary_378_inst_req_1,binary_378_inst_ack_1,sl_one,"binary_378_inst",false,iNsTr_13_373 & type_cast_377_wire_constant,
    false,exitcond1_379);
    -- shared split operator group (3) : binary_378_inst 
    ApIntEq_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_13_373;
      exitcond1_379 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_378_inst_req_0;
      reqR(0) <= binary_378_inst_req_1;
      binary_378_inst_ack_0 <= ackL(0); 
      binary_378_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000001000000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_363_load_0_req_0,ptr_deref_363_load_0_ack_0,ptr_deref_363_load_0_req_1,ptr_deref_363_load_0_ack_1,sl_one,"ptr_deref_363_load_0",false,ptr_deref_363_word_address_0,
    false,ptr_deref_363_data_0);
    -- shared load operator group (0) : ptr_deref_363_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(6 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_363_load_0_req_0,
        ptr_deref_363_load_0_ack_0,
        ptr_deref_363_load_0_req_1,
        ptr_deref_363_load_0_ack_1,
        "ptr_deref_363_load_0",
        "memory_space_2" ,
        ptr_deref_363_data_0,
        ptr_deref_363_word_address_0,
        "ptr_deref_363_data_0",
        "ptr_deref_363_word_address_0" -- 
      );
      reqL_unguarded(0) <= ptr_deref_363_load_0_req_0;
      ptr_deref_363_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_363_load_0_req_1;
      ptr_deref_363_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_363_word_address_0;
      ptr_deref_363_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(6 downto 0),
          mtag => memory_space_2_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 1,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_309_store_0_req_0,ptr_deref_309_store_0_ack_0,ptr_deref_309_store_0_req_1,ptr_deref_309_store_0_ack_1,sl_one,"ptr_deref_309_store_0",false,ptr_deref_309_word_address_0 & ptr_deref_309_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_309_store_0_req_0,
      ptr_deref_309_store_0_ack_0,
      ptr_deref_309_store_0_req_1,
      ptr_deref_309_store_0_ack_1,
      "ptr_deref_309_store_0",
      "memory_space_0" ,
      ptr_deref_309_data_0,
      ptr_deref_309_word_address_0,
      "ptr_deref_309_data_0",
      "ptr_deref_309_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_309_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(6 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_309_store_0_req_0;
      ptr_deref_309_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_309_store_0_req_1;
      ptr_deref_309_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_309_word_address_0;
      data_in <= ptr_deref_309_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_0_sr_req(0),
          mack => memory_space_0_sr_ack(0),
          maddr => memory_space_0_sr_addr(6 downto 0),
          mdata => memory_space_0_sr_data(31 downto 0),
          mtag => memory_space_0_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_0_sc_req(0),
          mack => memory_space_0_sc_ack(0),
          mtag => memory_space_0_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_313_store_0_req_0,ptr_deref_313_store_0_ack_0,ptr_deref_313_store_0_req_1,ptr_deref_313_store_0_ack_1,sl_one,"ptr_deref_313_store_0",false,ptr_deref_313_word_address_0 & ptr_deref_313_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_313_store_0_req_0,
      ptr_deref_313_store_0_ack_0,
      ptr_deref_313_store_0_req_1,
      ptr_deref_313_store_0_ack_1,
      "ptr_deref_313_store_0",
      "memory_space_1" ,
      ptr_deref_313_data_0,
      ptr_deref_313_word_address_0,
      "ptr_deref_313_data_0",
      "ptr_deref_313_word_address_0" -- 
    );
    -- shared store operator group (1) : ptr_deref_313_store_0 
    StoreGroup1: Block -- 
      signal addr_in: std_logic_vector(6 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= ptr_deref_313_store_0_req_0;
      ptr_deref_313_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ptr_deref_313_store_0_req_1;
      ptr_deref_313_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_313_word_address_0;
      data_in <= ptr_deref_313_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 1,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_1_sr_req(0),
          mack => memory_space_1_sr_ack(0),
          maddr => memory_space_1_sr_addr(6 downto 0),
          mdata => memory_space_1_sr_data(31 downto 0),
          mtag => memory_space_1_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 1,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_1_sc_req(0),
          mack => memory_space_1_sc_ack(0),
          mtag => memory_space_1_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 1
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_306_inst_req_0,simple_obj_ref_306_inst_ack_0,sl_one,"simple_obj_ref_306_inst  PipeRead from in_data_pipe",true, slv_zero,
    false,iNsTr_2_307);
    -- shared inport operator group (0) : simple_obj_ref_306_inst 
    InportGroup0: Block -- 
      signal data_out: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      -- logging on!
      process(clk)  begin -- 
        if clk'event and clk = '1' then -- 
          if simple_obj_ref_306_inst_ack_0 then -- 
            assert false report " ReadPipe in_data_pipe to wire iNsTr_2_307 value="  &  convert_slv_to_hex_string(data_out(31 downto 0))  severity note; --
          end if;
          --
        end if;
        -- 
      end process;
      req_unguarded(0) <= simple_obj_ref_306_inst_req_0;
      simple_obj_ref_306_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      iNsTr_2_307 <= data_out(31 downto 0);
      in_data_pipe_read_0: InputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (-- 
          req => req , 
          ack => ack , 
          data => data_out, 
          oreq => in_data_pipe_pipe_read_req(0),
          oack => in_data_pipe_pipe_read_ack(0),
          odata => in_data_pipe_pipe_read_data(31 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_365_inst_req_0,simple_obj_ref_365_inst_ack_0,sl_one,"simple_obj_ref_365_inst  PipeWrite to out_data_pipe",false,iNsTr_10_364,
    true, slv_zero);
    -- logging on!
    process(clk)  begin -- 
      if clk'event and clk = '1' then -- 
        if simple_obj_ref_365_inst_ack_0 then -- 
          assert false report " WritePipe out_data_pipe from wire iNsTr_10_364 value="  &  convert_slv_to_hex_string(iNsTr_10_364) severity note; --
        end if;
        --
      end if;
      -- 
    end process;
    -- shared outport operator group (0) : simple_obj_ref_365_inst 
    OutportGroup0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal req, ack : BooleanArray( 0 downto 0);
      signal req_unguarded, ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      req_unguarded(0) <= simple_obj_ref_365_inst_req_0;
      simple_obj_ref_365_inst_ack_0 <= ack_unguarded(0);
      guard_vector(0)  <=  '1';
      gI: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => req_unguarded,
        ackL => ack_unguarded,
        reqR => req,
        ackR => ack,
        guards => guard_vector); -- 
      data_in <= iNsTr_10_364;
      out_data_pipe_write_0: OutputPort -- 
        generic map ( data_width => 32,  num_reqs => 1,  no_arbitration => false)
        port map (--
          req => req , 
          ack => ack , 
          data => data_in, 
          oreq => out_data_pipe_pipe_write_req(0),
          oack => out_data_pipe_pipe_write_ack(0),
          odata => out_data_pipe_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,call_stmt_345_call_req_0,call_stmt_345_call_ack_0,call_stmt_345_call_req_1,call_stmt_345_call_ack_1,sl_one,"call_stmt_345_call",true, slv_zero,
    true, slv_zero);
    -- shared call operator group (0) : call_stmt_345_call 
    x_vectorSum_x_call_group_0: Block -- 
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_345_call_req_0;
      call_stmt_345_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_345_call_req_1;
      call_stmt_345_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 1) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      CallReq: InputMuxBaseNoData -- 
        generic map (  twidth => 1,
        nreqs => 1,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          reqR => x_vectorSum_x_call_reqs(0),
          ackR => x_vectorSum_x_call_acks(0),
          tagR => x_vectorSum_x_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( 
        twidth => 1, nreqs => 1, no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => x_vectorSum_x_return_acks(0), -- cross-over
          ackL => x_vectorSum_x_return_reqs(0), -- cross-over
          tagL => x_vectorSum_x_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity x_vectorSum_x is -- 
  generic (tag_length : integer); 
  port ( -- 
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic;
    memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_1_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
    memory_space_0_lr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_0_lc_tag :  in  std_logic_vector(3 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
  );
  -- 
end entity x_vectorSum_x;
architecture Default of x_vectorSum_x is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal start_req_symbol: Boolean;
  signal start_ack_symbol: Boolean;
  signal fin_req_symbol: Boolean;
  signal fin_ack_symbol: Boolean;
  signal tag_push, tag_pop: std_logic; 
  signal start_ack_sig, fin_ack_sig: std_logic; 
  -- output port buffer signals
  signal x_vectorSum_x_xCP_1292_start: Boolean;
  -- links between control-path and data-path
  signal array_obj_ref_425_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_425_index_0_resize_req_0 : boolean;
  signal array_obj_ref_430_root_address_inst_ack_0 : boolean;
  signal binary_437_inst_ack_1 : boolean;
  signal array_obj_ref_420_offset_inst_req_0 : boolean;
  signal array_obj_ref_420_offset_inst_ack_0 : boolean;
  signal array_obj_ref_551_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_420_root_address_inst_req_0 : boolean;
  signal addr_of_452_final_reg_req_0 : boolean;
  signal array_obj_ref_561_offset_inst_req_0 : boolean;
  signal array_obj_ref_556_offset_inst_req_0 : boolean;
  signal array_obj_ref_556_index_0_resize_req_0 : boolean;
  signal array_obj_ref_446_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_425_offset_inst_ack_0 : boolean;
  signal array_obj_ref_446_index_0_resize_ack_0 : boolean;
  signal binary_458_inst_req_1 : boolean;
  signal addr_of_452_final_reg_ack_0 : boolean;
  signal array_obj_ref_425_index_0_rename_ack_0 : boolean;
  signal addr_of_447_final_reg_ack_0 : boolean;
  signal array_obj_ref_446_root_address_inst_req_0 : boolean;
  signal array_obj_ref_430_offset_inst_ack_0 : boolean;
  signal addr_of_557_final_reg_ack_0 : boolean;
  signal addr_of_567_final_reg_ack_0 : boolean;
  signal array_obj_ref_446_index_0_rename_req_0 : boolean;
  signal addr_of_447_final_reg_req_0 : boolean;
  signal array_obj_ref_425_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_420_index_0_rename_req_0 : boolean;
  signal array_obj_ref_420_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_462_index_0_rename_req_0 : boolean;
  signal array_obj_ref_425_root_address_inst_req_0 : boolean;
  signal array_obj_ref_441_index_0_resize_req_0 : boolean;
  signal binary_458_inst_ack_1 : boolean;
  signal array_obj_ref_446_index_0_resize_req_0 : boolean;
  signal array_obj_ref_441_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_420_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_441_index_0_rename_req_0 : boolean;
  signal array_obj_ref_441_index_0_resize_ack_0 : boolean;
  signal addr_of_426_final_reg_req_0 : boolean;
  signal array_obj_ref_566_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_462_root_address_inst_req_0 : boolean;
  signal array_obj_ref_451_offset_inst_ack_0 : boolean;
  signal array_obj_ref_462_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_425_offset_inst_req_0 : boolean;
  signal array_obj_ref_430_offset_inst_req_0 : boolean;
  signal addr_of_426_final_reg_ack_0 : boolean;
  signal array_obj_ref_451_root_address_inst_req_0 : boolean;
  signal addr_of_442_final_reg_ack_0 : boolean;
  signal array_obj_ref_451_index_0_resize_req_0 : boolean;
  signal array_obj_ref_441_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_446_root_address_inst_ack_0 : boolean;
  signal addr_of_431_final_reg_req_0 : boolean;
  signal addr_of_557_final_reg_req_0 : boolean;
  signal array_obj_ref_551_offset_inst_req_0 : boolean;
  signal binary_437_inst_req_1 : boolean;
  signal array_obj_ref_420_index_0_resize_req_0 : boolean;
  signal addr_of_431_final_reg_ack_0 : boolean;
  signal array_obj_ref_430_root_address_inst_req_0 : boolean;
  signal array_obj_ref_425_index_0_rename_req_0 : boolean;
  signal array_obj_ref_462_index_0_resize_req_0 : boolean;
  signal array_obj_ref_462_offset_inst_ack_0 : boolean;
  signal array_obj_ref_446_offset_inst_req_0 : boolean;
  signal array_obj_ref_462_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_451_index_0_rename_req_0 : boolean;
  signal addr_of_463_final_reg_ack_0 : boolean;
  signal array_obj_ref_451_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_446_offset_inst_ack_0 : boolean;
  signal array_obj_ref_462_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_420_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_451_root_address_inst_ack_0 : boolean;
  signal addr_of_421_final_reg_req_0 : boolean;
  signal addr_of_421_final_reg_ack_0 : boolean;
  signal binary_458_inst_req_0 : boolean;
  signal array_obj_ref_451_index_0_resize_ack_0 : boolean;
  signal binary_458_inst_ack_0 : boolean;
  signal array_obj_ref_441_offset_inst_req_0 : boolean;
  signal array_obj_ref_441_offset_inst_ack_0 : boolean;
  signal array_obj_ref_430_index_0_resize_req_0 : boolean;
  signal array_obj_ref_430_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_430_index_0_rename_req_0 : boolean;
  signal array_obj_ref_430_index_0_rename_ack_0 : boolean;
  signal addr_of_442_final_reg_req_0 : boolean;
  signal addr_of_463_final_reg_req_0 : boolean;
  signal array_obj_ref_451_offset_inst_req_0 : boolean;
  signal array_obj_ref_441_root_address_inst_req_0 : boolean;
  signal array_obj_ref_462_offset_inst_req_0 : boolean;
  signal binary_437_inst_ack_0 : boolean;
  signal binary_437_inst_req_0 : boolean;
  signal array_obj_ref_551_offset_inst_ack_0 : boolean;
  signal array_obj_ref_561_offset_inst_ack_0 : boolean;
  signal array_obj_ref_561_index_0_resize_ack_0 : boolean;
  signal addr_of_552_final_reg_req_0 : boolean;
  signal addr_of_552_final_reg_ack_0 : boolean;
  signal array_obj_ref_566_offset_inst_req_0 : boolean;
  signal array_obj_ref_571_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_551_index_0_resize_req_0 : boolean;
  signal array_obj_ref_556_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_551_index_0_resize_ack_0 : boolean;
  signal ptr_deref_732_gather_scatter_req_0 : boolean;
  signal array_obj_ref_566_index_0_rename_req_0 : boolean;
  signal array_obj_ref_556_offset_inst_ack_0 : boolean;
  signal array_obj_ref_551_index_0_rename_req_0 : boolean;
  signal array_obj_ref_551_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_566_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_556_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_561_root_address_inst_req_0 : boolean;
  signal array_obj_ref_561_root_address_inst_ack_0 : boolean;
  signal addr_of_567_final_reg_req_0 : boolean;
  signal array_obj_ref_551_root_address_inst_req_0 : boolean;
  signal array_obj_ref_561_index_0_resize_req_0 : boolean;
  signal array_obj_ref_566_offset_inst_ack_0 : boolean;
  signal array_obj_ref_566_index_0_resize_req_0 : boolean;
  signal ptr_deref_732_gather_scatter_ack_0 : boolean;
  signal array_obj_ref_556_root_address_inst_req_0 : boolean;
  signal array_obj_ref_556_index_0_rename_req_0 : boolean;
  signal array_obj_ref_561_index_0_rename_req_0 : boolean;
  signal array_obj_ref_571_index_0_rename_req_0 : boolean;
  signal array_obj_ref_556_root_address_inst_ack_0 : boolean;
  signal array_obj_ref_566_root_address_inst_req_0 : boolean;
  signal array_obj_ref_571_offset_inst_req_0 : boolean;
  signal array_obj_ref_561_index_0_rename_ack_0 : boolean;
  signal addr_of_562_final_reg_req_0 : boolean;
  signal addr_of_562_final_reg_ack_0 : boolean;
  signal array_obj_ref_571_index_0_resize_req_0 : boolean;
  signal array_obj_ref_571_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_566_index_0_rename_ack_0 : boolean;
  signal phi_stmt_400_req_0 : boolean;
  signal phi_stmt_400_req_1 : boolean;
  signal phi_stmt_400_ack_0 : boolean;
  signal type_cast_403_inst_req_0 : boolean;
  signal type_cast_403_inst_ack_0 : boolean;
  signal binary_410_inst_req_0 : boolean;
  signal binary_410_inst_ack_0 : boolean;
  signal binary_410_inst_req_1 : boolean;
  signal binary_410_inst_ack_1 : boolean;
  signal binary_416_inst_req_0 : boolean;
  signal binary_416_inst_ack_0 : boolean;
  signal binary_416_inst_req_1 : boolean;
  signal binary_416_inst_ack_1 : boolean;
  signal array_obj_ref_467_index_0_resize_req_0 : boolean;
  signal array_obj_ref_467_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_467_index_0_rename_req_0 : boolean;
  signal array_obj_ref_467_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_467_offset_inst_req_0 : boolean;
  signal array_obj_ref_467_offset_inst_ack_0 : boolean;
  signal array_obj_ref_467_root_address_inst_req_0 : boolean;
  signal array_obj_ref_467_root_address_inst_ack_0 : boolean;
  signal addr_of_468_final_reg_req_0 : boolean;
  signal addr_of_468_final_reg_ack_0 : boolean;
  signal ptr_deref_713_store_0_ack_0 : boolean;
  signal array_obj_ref_472_index_0_resize_req_0 : boolean;
  signal array_obj_ref_472_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_472_index_0_rename_req_0 : boolean;
  signal array_obj_ref_472_index_0_rename_ack_0 : boolean;
  signal ptr_deref_713_store_0_req_0 : boolean;
  signal array_obj_ref_472_offset_inst_req_0 : boolean;
  signal array_obj_ref_472_offset_inst_ack_0 : boolean;
  signal ptr_deref_732_addr_0_req_0 : boolean;
  signal simple_obj_ref_766_inst_req_0 : boolean;
  signal array_obj_ref_472_root_address_inst_req_0 : boolean;
  signal array_obj_ref_472_root_address_inst_ack_0 : boolean;
  signal addr_of_473_final_reg_req_0 : boolean;
  signal addr_of_473_final_reg_ack_0 : boolean;
  signal array_obj_ref_571_offset_inst_ack_0 : boolean;
  signal simple_obj_ref_760_inst_req_0 : boolean;
  signal simple_obj_ref_735_inst_ack_0 : boolean;
  signal ptr_deref_713_gather_scatter_ack_0 : boolean;
  signal binary_479_inst_req_0 : boolean;
  signal binary_479_inst_ack_0 : boolean;
  signal binary_479_inst_req_1 : boolean;
  signal binary_479_inst_ack_1 : boolean;
  signal ptr_deref_713_gather_scatter_req_0 : boolean;
  signal simple_obj_ref_722_inst_req_0 : boolean;
  signal ptr_deref_751_store_0_ack_0 : boolean;
  signal array_obj_ref_483_index_0_resize_req_0 : boolean;
  signal simple_obj_ref_738_inst_ack_0 : boolean;
  signal array_obj_ref_483_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_483_index_0_rename_req_0 : boolean;
  signal array_obj_ref_483_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_483_offset_inst_req_0 : boolean;
  signal array_obj_ref_483_offset_inst_ack_0 : boolean;
  signal array_obj_ref_483_root_address_inst_req_0 : boolean;
  signal array_obj_ref_483_root_address_inst_ack_0 : boolean;
  signal addr_of_484_final_reg_req_0 : boolean;
  signal addr_of_484_final_reg_ack_0 : boolean;
  signal simple_obj_ref_735_inst_req_0 : boolean;
  signal array_obj_ref_488_index_0_resize_req_0 : boolean;
  signal array_obj_ref_488_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_488_index_0_rename_req_0 : boolean;
  signal array_obj_ref_488_index_0_rename_ack_0 : boolean;
  signal simple_obj_ref_719_inst_ack_0 : boolean;
  signal array_obj_ref_488_offset_inst_req_0 : boolean;
  signal array_obj_ref_488_offset_inst_ack_0 : boolean;
  signal array_obj_ref_488_root_address_inst_req_0 : boolean;
  signal array_obj_ref_488_root_address_inst_ack_0 : boolean;
  signal addr_of_489_final_reg_req_0 : boolean;
  signal addr_of_489_final_reg_ack_0 : boolean;
  signal simple_obj_ref_722_inst_ack_0 : boolean;
  signal array_obj_ref_493_index_0_resize_req_0 : boolean;
  signal array_obj_ref_493_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_493_index_0_rename_req_0 : boolean;
  signal array_obj_ref_493_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_493_offset_inst_req_0 : boolean;
  signal array_obj_ref_493_offset_inst_ack_0 : boolean;
  signal array_obj_ref_493_root_address_inst_req_0 : boolean;
  signal array_obj_ref_493_root_address_inst_ack_0 : boolean;
  signal addr_of_494_final_reg_req_0 : boolean;
  signal addr_of_494_final_reg_ack_0 : boolean;
  signal ptr_deref_713_addr_0_ack_0 : boolean;
  signal ptr_deref_751_store_0_req_0 : boolean;
  signal ptr_deref_732_root_address_inst_ack_0 : boolean;
  signal simple_obj_ref_719_inst_req_0 : boolean;
  signal binary_500_inst_req_0 : boolean;
  signal binary_500_inst_ack_0 : boolean;
  signal binary_500_inst_req_1 : boolean;
  signal binary_500_inst_ack_1 : boolean;
  signal ptr_deref_732_store_0_ack_0 : boolean;
  signal array_obj_ref_504_index_0_resize_req_0 : boolean;
  signal array_obj_ref_504_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_504_index_0_rename_req_0 : boolean;
  signal simple_obj_ref_728_inst_req_0 : boolean;
  signal array_obj_ref_504_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_504_offset_inst_req_0 : boolean;
  signal array_obj_ref_504_offset_inst_ack_0 : boolean;
  signal array_obj_ref_504_root_address_inst_req_0 : boolean;
  signal array_obj_ref_504_root_address_inst_ack_0 : boolean;
  signal addr_of_505_final_reg_req_0 : boolean;
  signal addr_of_505_final_reg_ack_0 : boolean;
  signal simple_obj_ref_728_inst_ack_0 : boolean;
  signal array_obj_ref_509_index_0_resize_req_0 : boolean;
  signal array_obj_ref_509_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_509_index_0_rename_req_0 : boolean;
  signal array_obj_ref_509_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_509_offset_inst_req_0 : boolean;
  signal array_obj_ref_509_offset_inst_ack_0 : boolean;
  signal array_obj_ref_509_root_address_inst_req_0 : boolean;
  signal array_obj_ref_509_root_address_inst_ack_0 : boolean;
  signal addr_of_510_final_reg_req_0 : boolean;
  signal addr_of_510_final_reg_ack_0 : boolean;
  signal array_obj_ref_514_index_0_resize_req_0 : boolean;
  signal array_obj_ref_514_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_514_index_0_rename_req_0 : boolean;
  signal array_obj_ref_514_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_514_offset_inst_req_0 : boolean;
  signal array_obj_ref_514_offset_inst_ack_0 : boolean;
  signal array_obj_ref_514_root_address_inst_req_0 : boolean;
  signal array_obj_ref_514_root_address_inst_ack_0 : boolean;
  signal addr_of_515_final_reg_req_0 : boolean;
  signal addr_of_515_final_reg_ack_0 : boolean;
  signal binary_521_inst_req_0 : boolean;
  signal binary_521_inst_ack_0 : boolean;
  signal binary_521_inst_req_1 : boolean;
  signal binary_521_inst_ack_1 : boolean;
  signal array_obj_ref_525_index_0_resize_req_0 : boolean;
  signal array_obj_ref_525_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_525_index_0_rename_req_0 : boolean;
  signal array_obj_ref_525_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_525_offset_inst_req_0 : boolean;
  signal array_obj_ref_525_offset_inst_ack_0 : boolean;
  signal array_obj_ref_525_root_address_inst_req_0 : boolean;
  signal array_obj_ref_525_root_address_inst_ack_0 : boolean;
  signal addr_of_526_final_reg_req_0 : boolean;
  signal addr_of_526_final_reg_ack_0 : boolean;
  signal array_obj_ref_530_index_0_resize_req_0 : boolean;
  signal array_obj_ref_530_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_530_index_0_rename_req_0 : boolean;
  signal array_obj_ref_530_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_530_offset_inst_req_0 : boolean;
  signal array_obj_ref_530_offset_inst_ack_0 : boolean;
  signal array_obj_ref_530_root_address_inst_req_0 : boolean;
  signal array_obj_ref_530_root_address_inst_ack_0 : boolean;
  signal addr_of_531_final_reg_req_0 : boolean;
  signal addr_of_531_final_reg_ack_0 : boolean;
  signal array_obj_ref_535_index_0_resize_req_0 : boolean;
  signal array_obj_ref_535_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_535_index_0_rename_req_0 : boolean;
  signal array_obj_ref_535_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_535_offset_inst_req_0 : boolean;
  signal array_obj_ref_535_offset_inst_ack_0 : boolean;
  signal array_obj_ref_535_root_address_inst_req_0 : boolean;
  signal array_obj_ref_535_root_address_inst_ack_0 : boolean;
  signal addr_of_536_final_reg_req_0 : boolean;
  signal addr_of_536_final_reg_ack_0 : boolean;
  signal binary_542_inst_req_0 : boolean;
  signal binary_542_inst_ack_0 : boolean;
  signal binary_542_inst_req_1 : boolean;
  signal binary_542_inst_ack_1 : boolean;
  signal array_obj_ref_546_index_0_resize_req_0 : boolean;
  signal array_obj_ref_546_index_0_resize_ack_0 : boolean;
  signal array_obj_ref_546_index_0_rename_req_0 : boolean;
  signal array_obj_ref_546_index_0_rename_ack_0 : boolean;
  signal array_obj_ref_546_offset_inst_req_0 : boolean;
  signal array_obj_ref_546_offset_inst_ack_0 : boolean;
  signal array_obj_ref_546_root_address_inst_req_0 : boolean;
  signal array_obj_ref_546_root_address_inst_ack_0 : boolean;
  signal addr_of_547_final_reg_req_0 : boolean;
  signal addr_of_547_final_reg_ack_0 : boolean;
  signal ptr_deref_751_base_resize_ack_0 : boolean;
  signal simple_obj_ref_754_inst_req_0 : boolean;
  signal ptr_deref_751_base_resize_req_0 : boolean;
  signal simple_obj_ref_754_inst_ack_0 : boolean;
  signal array_obj_ref_571_root_address_inst_req_0 : boolean;
  signal array_obj_ref_571_root_address_inst_ack_0 : boolean;
  signal addr_of_572_final_reg_req_0 : boolean;
  signal addr_of_572_final_reg_ack_0 : boolean;
  signal ptr_deref_576_base_resize_req_0 : boolean;
  signal ptr_deref_576_base_resize_ack_0 : boolean;
  signal ptr_deref_576_root_address_inst_req_0 : boolean;
  signal ptr_deref_576_root_address_inst_ack_0 : boolean;
  signal ptr_deref_576_addr_0_req_0 : boolean;
  signal ptr_deref_576_addr_0_ack_0 : boolean;
  signal ptr_deref_576_load_0_req_0 : boolean;
  signal ptr_deref_576_load_0_ack_0 : boolean;
  signal ptr_deref_576_load_0_req_1 : boolean;
  signal ptr_deref_576_load_0_ack_1 : boolean;
  signal ptr_deref_576_gather_scatter_req_0 : boolean;
  signal ptr_deref_576_gather_scatter_ack_0 : boolean;
  signal ptr_deref_580_base_resize_req_0 : boolean;
  signal ptr_deref_580_base_resize_ack_0 : boolean;
  signal ptr_deref_580_root_address_inst_req_0 : boolean;
  signal ptr_deref_580_root_address_inst_ack_0 : boolean;
  signal ptr_deref_580_addr_0_req_0 : boolean;
  signal ptr_deref_580_addr_0_ack_0 : boolean;
  signal ptr_deref_580_load_0_req_0 : boolean;
  signal ptr_deref_580_load_0_ack_0 : boolean;
  signal ptr_deref_580_load_0_req_1 : boolean;
  signal ptr_deref_580_load_0_ack_1 : boolean;
  signal ptr_deref_580_gather_scatter_req_0 : boolean;
  signal ptr_deref_580_gather_scatter_ack_0 : boolean;
  signal binary_585_inst_req_0 : boolean;
  signal binary_585_inst_ack_0 : boolean;
  signal binary_585_inst_req_1 : boolean;
  signal binary_585_inst_ack_1 : boolean;
  signal ptr_deref_713_store_0_req_1 : boolean;
  signal ptr_deref_713_store_0_ack_1 : boolean;
  signal ptr_deref_589_base_resize_req_0 : boolean;
  signal ptr_deref_589_base_resize_ack_0 : boolean;
  signal ptr_deref_589_root_address_inst_req_0 : boolean;
  signal ptr_deref_589_root_address_inst_ack_0 : boolean;
  signal ptr_deref_589_addr_0_req_0 : boolean;
  signal ptr_deref_589_addr_0_ack_0 : boolean;
  signal ptr_deref_589_load_0_req_0 : boolean;
  signal ptr_deref_589_load_0_ack_0 : boolean;
  signal simple_obj_ref_747_inst_req_0 : boolean;
  signal ptr_deref_589_load_0_req_1 : boolean;
  signal ptr_deref_589_load_0_ack_1 : boolean;
  signal ptr_deref_589_gather_scatter_req_0 : boolean;
  signal ptr_deref_589_gather_scatter_ack_0 : boolean;
  signal ptr_deref_751_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_757_inst_ack_0 : boolean;
  signal ptr_deref_732_store_0_req_0 : boolean;
  signal ptr_deref_593_base_resize_req_0 : boolean;
  signal ptr_deref_593_base_resize_ack_0 : boolean;
  signal ptr_deref_593_root_address_inst_req_0 : boolean;
  signal ptr_deref_593_root_address_inst_ack_0 : boolean;
  signal ptr_deref_593_addr_0_req_0 : boolean;
  signal simple_obj_ref_747_inst_ack_0 : boolean;
  signal ptr_deref_593_addr_0_ack_0 : boolean;
  signal ptr_deref_593_load_0_req_0 : boolean;
  signal ptr_deref_593_load_0_ack_0 : boolean;
  signal ptr_deref_593_load_0_req_1 : boolean;
  signal ptr_deref_593_load_0_ack_1 : boolean;
  signal ptr_deref_593_gather_scatter_req_0 : boolean;
  signal ptr_deref_593_gather_scatter_ack_0 : boolean;
  signal ptr_deref_732_root_address_inst_req_0 : boolean;
  signal simple_obj_ref_760_inst_ack_0 : boolean;
  signal ptr_deref_751_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_738_inst_req_0 : boolean;
  signal ptr_deref_732_store_0_req_1 : boolean;
  signal simple_obj_ref_716_inst_req_0 : boolean;
  signal simple_obj_ref_716_inst_ack_0 : boolean;
  signal binary_598_inst_req_0 : boolean;
  signal binary_598_inst_ack_0 : boolean;
  signal binary_598_inst_req_1 : boolean;
  signal binary_598_inst_ack_1 : boolean;
  signal ptr_deref_751_gather_scatter_req_0 : boolean;
  signal ptr_deref_602_base_resize_req_0 : boolean;
  signal ptr_deref_602_base_resize_ack_0 : boolean;
  signal ptr_deref_732_addr_0_ack_0 : boolean;
  signal ptr_deref_602_root_address_inst_req_0 : boolean;
  signal ptr_deref_602_root_address_inst_ack_0 : boolean;
  signal ptr_deref_602_addr_0_req_0 : boolean;
  signal ptr_deref_602_addr_0_ack_0 : boolean;
  signal simple_obj_ref_741_inst_req_0 : boolean;
  signal ptr_deref_602_load_0_req_0 : boolean;
  signal ptr_deref_602_load_0_ack_0 : boolean;
  signal ptr_deref_602_load_0_req_1 : boolean;
  signal ptr_deref_602_load_0_ack_1 : boolean;
  signal ptr_deref_602_gather_scatter_req_0 : boolean;
  signal ptr_deref_602_gather_scatter_ack_0 : boolean;
  signal simple_obj_ref_744_inst_req_0 : boolean;
  signal simple_obj_ref_744_inst_ack_0 : boolean;
  signal simple_obj_ref_757_inst_req_0 : boolean;
  signal ptr_deref_732_store_0_ack_1 : boolean;
  signal ptr_deref_606_base_resize_req_0 : boolean;
  signal ptr_deref_606_base_resize_ack_0 : boolean;
  signal ptr_deref_606_root_address_inst_req_0 : boolean;
  signal ptr_deref_606_root_address_inst_ack_0 : boolean;
  signal ptr_deref_606_addr_0_req_0 : boolean;
  signal ptr_deref_606_addr_0_ack_0 : boolean;
  signal simple_obj_ref_741_inst_ack_0 : boolean;
  signal ptr_deref_606_load_0_req_0 : boolean;
  signal ptr_deref_606_load_0_ack_0 : boolean;
  signal ptr_deref_606_load_0_req_1 : boolean;
  signal ptr_deref_606_load_0_ack_1 : boolean;
  signal ptr_deref_606_gather_scatter_req_0 : boolean;
  signal ptr_deref_606_gather_scatter_ack_0 : boolean;
  signal ptr_deref_732_base_resize_req_0 : boolean;
  signal ptr_deref_732_base_resize_ack_0 : boolean;
  signal binary_611_inst_req_0 : boolean;
  signal binary_611_inst_ack_0 : boolean;
  signal binary_611_inst_req_1 : boolean;
  signal binary_611_inst_ack_1 : boolean;
  signal ptr_deref_615_base_resize_req_0 : boolean;
  signal ptr_deref_615_base_resize_ack_0 : boolean;
  signal ptr_deref_615_root_address_inst_req_0 : boolean;
  signal ptr_deref_615_root_address_inst_ack_0 : boolean;
  signal ptr_deref_615_addr_0_req_0 : boolean;
  signal ptr_deref_615_addr_0_ack_0 : boolean;
  signal ptr_deref_615_load_0_req_0 : boolean;
  signal ptr_deref_615_load_0_ack_0 : boolean;
  signal ptr_deref_615_load_0_req_1 : boolean;
  signal ptr_deref_615_load_0_ack_1 : boolean;
  signal ptr_deref_615_gather_scatter_req_0 : boolean;
  signal ptr_deref_615_gather_scatter_ack_0 : boolean;
  signal ptr_deref_619_base_resize_req_0 : boolean;
  signal ptr_deref_619_base_resize_ack_0 : boolean;
  signal ptr_deref_619_root_address_inst_req_0 : boolean;
  signal ptr_deref_619_root_address_inst_ack_0 : boolean;
  signal ptr_deref_619_addr_0_req_0 : boolean;
  signal ptr_deref_619_addr_0_ack_0 : boolean;
  signal ptr_deref_619_load_0_req_0 : boolean;
  signal ptr_deref_619_load_0_ack_0 : boolean;
  signal ptr_deref_619_load_0_req_1 : boolean;
  signal ptr_deref_619_load_0_ack_1 : boolean;
  signal ptr_deref_619_gather_scatter_req_0 : boolean;
  signal ptr_deref_619_gather_scatter_ack_0 : boolean;
  signal binary_624_inst_req_0 : boolean;
  signal binary_624_inst_ack_0 : boolean;
  signal binary_624_inst_req_1 : boolean;
  signal binary_624_inst_ack_1 : boolean;
  signal ptr_deref_628_base_resize_req_0 : boolean;
  signal ptr_deref_628_base_resize_ack_0 : boolean;
  signal ptr_deref_628_root_address_inst_req_0 : boolean;
  signal ptr_deref_628_root_address_inst_ack_0 : boolean;
  signal ptr_deref_628_addr_0_req_0 : boolean;
  signal ptr_deref_628_addr_0_ack_0 : boolean;
  signal ptr_deref_628_load_0_req_0 : boolean;
  signal ptr_deref_628_load_0_ack_0 : boolean;
  signal ptr_deref_628_load_0_req_1 : boolean;
  signal ptr_deref_628_load_0_ack_1 : boolean;
  signal ptr_deref_628_gather_scatter_req_0 : boolean;
  signal ptr_deref_628_gather_scatter_ack_0 : boolean;
  signal ptr_deref_632_base_resize_req_0 : boolean;
  signal ptr_deref_632_base_resize_ack_0 : boolean;
  signal ptr_deref_632_root_address_inst_req_0 : boolean;
  signal ptr_deref_632_root_address_inst_ack_0 : boolean;
  signal ptr_deref_632_addr_0_req_0 : boolean;
  signal ptr_deref_632_addr_0_ack_0 : boolean;
  signal ptr_deref_632_load_0_req_0 : boolean;
  signal ptr_deref_632_load_0_ack_0 : boolean;
  signal ptr_deref_632_load_0_req_1 : boolean;
  signal ptr_deref_632_load_0_ack_1 : boolean;
  signal ptr_deref_632_gather_scatter_req_0 : boolean;
  signal ptr_deref_632_gather_scatter_ack_0 : boolean;
  signal binary_637_inst_req_0 : boolean;
  signal binary_637_inst_ack_0 : boolean;
  signal binary_637_inst_req_1 : boolean;
  signal binary_637_inst_ack_1 : boolean;
  signal ptr_deref_641_base_resize_req_0 : boolean;
  signal ptr_deref_641_base_resize_ack_0 : boolean;
  signal ptr_deref_641_root_address_inst_req_0 : boolean;
  signal ptr_deref_641_root_address_inst_ack_0 : boolean;
  signal ptr_deref_641_addr_0_req_0 : boolean;
  signal ptr_deref_641_addr_0_ack_0 : boolean;
  signal ptr_deref_641_load_0_req_0 : boolean;
  signal ptr_deref_641_load_0_ack_0 : boolean;
  signal ptr_deref_641_load_0_req_1 : boolean;
  signal ptr_deref_641_load_0_ack_1 : boolean;
  signal ptr_deref_641_gather_scatter_req_0 : boolean;
  signal ptr_deref_641_gather_scatter_ack_0 : boolean;
  signal ptr_deref_645_base_resize_req_0 : boolean;
  signal ptr_deref_645_base_resize_ack_0 : boolean;
  signal ptr_deref_645_root_address_inst_req_0 : boolean;
  signal ptr_deref_645_root_address_inst_ack_0 : boolean;
  signal ptr_deref_645_addr_0_req_0 : boolean;
  signal ptr_deref_645_addr_0_ack_0 : boolean;
  signal ptr_deref_645_load_0_req_0 : boolean;
  signal ptr_deref_645_load_0_ack_0 : boolean;
  signal ptr_deref_645_load_0_req_1 : boolean;
  signal ptr_deref_645_load_0_ack_1 : boolean;
  signal ptr_deref_645_gather_scatter_req_0 : boolean;
  signal ptr_deref_645_gather_scatter_ack_0 : boolean;
  signal binary_650_inst_req_0 : boolean;
  signal binary_650_inst_ack_0 : boolean;
  signal binary_650_inst_req_1 : boolean;
  signal binary_650_inst_ack_1 : boolean;
  signal ptr_deref_654_base_resize_req_0 : boolean;
  signal ptr_deref_654_base_resize_ack_0 : boolean;
  signal ptr_deref_654_root_address_inst_req_0 : boolean;
  signal ptr_deref_654_root_address_inst_ack_0 : boolean;
  signal ptr_deref_654_addr_0_req_0 : boolean;
  signal ptr_deref_654_addr_0_ack_0 : boolean;
  signal ptr_deref_654_load_0_req_0 : boolean;
  signal ptr_deref_654_load_0_ack_0 : boolean;
  signal ptr_deref_654_load_0_req_1 : boolean;
  signal ptr_deref_654_load_0_ack_1 : boolean;
  signal ptr_deref_654_gather_scatter_req_0 : boolean;
  signal ptr_deref_654_gather_scatter_ack_0 : boolean;
  signal ptr_deref_658_base_resize_req_0 : boolean;
  signal ptr_deref_658_base_resize_ack_0 : boolean;
  signal ptr_deref_658_root_address_inst_req_0 : boolean;
  signal ptr_deref_658_root_address_inst_ack_0 : boolean;
  signal ptr_deref_658_addr_0_req_0 : boolean;
  signal ptr_deref_658_addr_0_ack_0 : boolean;
  signal ptr_deref_658_load_0_req_0 : boolean;
  signal ptr_deref_658_load_0_ack_0 : boolean;
  signal ptr_deref_658_load_0_req_1 : boolean;
  signal ptr_deref_658_load_0_ack_1 : boolean;
  signal ptr_deref_658_gather_scatter_req_0 : boolean;
  signal ptr_deref_658_gather_scatter_ack_0 : boolean;
  signal binary_663_inst_req_0 : boolean;
  signal binary_663_inst_ack_0 : boolean;
  signal binary_663_inst_req_1 : boolean;
  signal binary_663_inst_ack_1 : boolean;
  signal ptr_deref_667_base_resize_req_0 : boolean;
  signal ptr_deref_667_base_resize_ack_0 : boolean;
  signal ptr_deref_667_root_address_inst_req_0 : boolean;
  signal ptr_deref_667_root_address_inst_ack_0 : boolean;
  signal ptr_deref_667_addr_0_req_0 : boolean;
  signal ptr_deref_667_addr_0_ack_0 : boolean;
  signal ptr_deref_667_load_0_req_0 : boolean;
  signal ptr_deref_667_load_0_ack_0 : boolean;
  signal ptr_deref_667_load_0_req_1 : boolean;
  signal ptr_deref_667_load_0_ack_1 : boolean;
  signal ptr_deref_667_gather_scatter_req_0 : boolean;
  signal ptr_deref_667_gather_scatter_ack_0 : boolean;
  signal ptr_deref_671_base_resize_req_0 : boolean;
  signal ptr_deref_671_base_resize_ack_0 : boolean;
  signal ptr_deref_671_root_address_inst_req_0 : boolean;
  signal ptr_deref_671_root_address_inst_ack_0 : boolean;
  signal ptr_deref_671_addr_0_req_0 : boolean;
  signal ptr_deref_671_addr_0_ack_0 : boolean;
  signal ptr_deref_671_load_0_req_0 : boolean;
  signal ptr_deref_671_load_0_ack_0 : boolean;
  signal ptr_deref_671_load_0_req_1 : boolean;
  signal ptr_deref_671_load_0_ack_1 : boolean;
  signal ptr_deref_671_gather_scatter_req_0 : boolean;
  signal ptr_deref_671_gather_scatter_ack_0 : boolean;
  signal binary_676_inst_req_0 : boolean;
  signal binary_676_inst_ack_0 : boolean;
  signal binary_676_inst_req_1 : boolean;
  signal binary_676_inst_ack_1 : boolean;
  signal simple_obj_ref_678_inst_req_0 : boolean;
  signal simple_obj_ref_678_inst_ack_0 : boolean;
  signal ptr_deref_751_addr_0_ack_0 : boolean;
  signal simple_obj_ref_681_inst_req_0 : boolean;
  signal simple_obj_ref_681_inst_ack_0 : boolean;
  signal ptr_deref_751_addr_0_req_0 : boolean;
  signal simple_obj_ref_763_inst_ack_0 : boolean;
  signal simple_obj_ref_684_inst_req_0 : boolean;
  signal simple_obj_ref_684_inst_ack_0 : boolean;
  signal simple_obj_ref_766_inst_ack_0 : boolean;
  signal simple_obj_ref_763_inst_req_0 : boolean;
  signal ptr_deref_713_addr_0_req_0 : boolean;
  signal simple_obj_ref_687_inst_req_0 : boolean;
  signal simple_obj_ref_687_inst_ack_0 : boolean;
  signal ptr_deref_713_root_address_inst_ack_0 : boolean;
  signal ptr_deref_713_root_address_inst_req_0 : boolean;
  signal ptr_deref_751_store_0_ack_1 : boolean;
  signal ptr_deref_713_base_resize_ack_0 : boolean;
  signal ptr_deref_713_base_resize_req_0 : boolean;
  signal simple_obj_ref_725_inst_ack_0 : boolean;
  signal simple_obj_ref_725_inst_req_0 : boolean;
  signal ptr_deref_751_store_0_req_1 : boolean;
  signal simple_obj_ref_690_inst_req_0 : boolean;
  signal simple_obj_ref_690_inst_ack_0 : boolean;
  signal ptr_deref_751_root_address_inst_ack_0 : boolean;
  signal ptr_deref_694_base_resize_req_0 : boolean;
  signal ptr_deref_694_base_resize_ack_0 : boolean;
  signal ptr_deref_694_root_address_inst_req_0 : boolean;
  signal ptr_deref_694_root_address_inst_ack_0 : boolean;
  signal ptr_deref_694_addr_0_req_0 : boolean;
  signal ptr_deref_694_addr_0_ack_0 : boolean;
  signal ptr_deref_694_gather_scatter_req_0 : boolean;
  signal ptr_deref_694_gather_scatter_ack_0 : boolean;
  signal ptr_deref_694_store_0_req_0 : boolean;
  signal ptr_deref_694_store_0_ack_0 : boolean;
  signal ptr_deref_694_store_0_req_1 : boolean;
  signal ptr_deref_694_store_0_ack_1 : boolean;
  signal simple_obj_ref_697_inst_req_0 : boolean;
  signal simple_obj_ref_697_inst_ack_0 : boolean;
  signal simple_obj_ref_700_inst_req_0 : boolean;
  signal simple_obj_ref_700_inst_ack_0 : boolean;
  signal simple_obj_ref_703_inst_req_0 : boolean;
  signal simple_obj_ref_703_inst_ack_0 : boolean;
  signal simple_obj_ref_706_inst_req_0 : boolean;
  signal simple_obj_ref_706_inst_ack_0 : boolean;
  signal simple_obj_ref_709_inst_req_0 : boolean;
  signal simple_obj_ref_709_inst_ack_0 : boolean;
  signal ptr_deref_770_base_resize_req_0 : boolean;
  signal ptr_deref_770_base_resize_ack_0 : boolean;
  signal ptr_deref_770_root_address_inst_req_0 : boolean;
  signal ptr_deref_770_root_address_inst_ack_0 : boolean;
  signal ptr_deref_770_addr_0_req_0 : boolean;
  signal ptr_deref_770_addr_0_ack_0 : boolean;
  signal ptr_deref_770_gather_scatter_req_0 : boolean;
  signal ptr_deref_770_gather_scatter_ack_0 : boolean;
  signal ptr_deref_770_store_0_req_0 : boolean;
  signal ptr_deref_770_store_0_ack_0 : boolean;
  signal ptr_deref_770_store_0_req_1 : boolean;
  signal ptr_deref_770_store_0_ack_1 : boolean;
  signal simple_obj_ref_773_inst_req_0 : boolean;
  signal simple_obj_ref_773_inst_ack_0 : boolean;
  signal simple_obj_ref_776_inst_req_0 : boolean;
  signal simple_obj_ref_776_inst_ack_0 : boolean;
  signal simple_obj_ref_779_inst_req_0 : boolean;
  signal simple_obj_ref_779_inst_ack_0 : boolean;
  signal simple_obj_ref_782_inst_req_0 : boolean;
  signal simple_obj_ref_782_inst_ack_0 : boolean;
  signal simple_obj_ref_785_inst_req_0 : boolean;
  signal simple_obj_ref_785_inst_ack_0 : boolean;
  signal ptr_deref_789_base_resize_req_0 : boolean;
  signal ptr_deref_789_base_resize_ack_0 : boolean;
  signal ptr_deref_789_root_address_inst_req_0 : boolean;
  signal ptr_deref_789_root_address_inst_ack_0 : boolean;
  signal ptr_deref_789_addr_0_req_0 : boolean;
  signal ptr_deref_789_addr_0_ack_0 : boolean;
  signal ptr_deref_789_gather_scatter_req_0 : boolean;
  signal ptr_deref_789_gather_scatter_ack_0 : boolean;
  signal ptr_deref_789_store_0_req_0 : boolean;
  signal ptr_deref_789_store_0_ack_0 : boolean;
  signal ptr_deref_789_store_0_req_1 : boolean;
  signal ptr_deref_789_store_0_ack_1 : boolean;
  signal simple_obj_ref_792_inst_req_0 : boolean;
  signal simple_obj_ref_792_inst_ack_0 : boolean;
  signal simple_obj_ref_795_inst_req_0 : boolean;
  signal simple_obj_ref_795_inst_ack_0 : boolean;
  signal simple_obj_ref_798_inst_req_0 : boolean;
  signal simple_obj_ref_798_inst_ack_0 : boolean;
  signal simple_obj_ref_801_inst_req_0 : boolean;
  signal simple_obj_ref_801_inst_ack_0 : boolean;
  signal simple_obj_ref_804_inst_req_0 : boolean;
  signal simple_obj_ref_804_inst_ack_0 : boolean;
  signal ptr_deref_808_base_resize_req_0 : boolean;
  signal ptr_deref_808_base_resize_ack_0 : boolean;
  signal ptr_deref_808_root_address_inst_req_0 : boolean;
  signal ptr_deref_808_root_address_inst_ack_0 : boolean;
  signal ptr_deref_808_addr_0_req_0 : boolean;
  signal ptr_deref_808_addr_0_ack_0 : boolean;
  signal ptr_deref_808_gather_scatter_req_0 : boolean;
  signal ptr_deref_808_gather_scatter_ack_0 : boolean;
  signal ptr_deref_808_store_0_req_0 : boolean;
  signal ptr_deref_808_store_0_ack_0 : boolean;
  signal ptr_deref_808_store_0_req_1 : boolean;
  signal ptr_deref_808_store_0_ack_1 : boolean;
  signal simple_obj_ref_811_inst_req_0 : boolean;
  signal simple_obj_ref_811_inst_ack_0 : boolean;
  signal simple_obj_ref_814_inst_req_0 : boolean;
  signal simple_obj_ref_814_inst_ack_0 : boolean;
  signal simple_obj_ref_817_inst_req_0 : boolean;
  signal simple_obj_ref_817_inst_ack_0 : boolean;
  signal simple_obj_ref_820_inst_req_0 : boolean;
  signal simple_obj_ref_820_inst_ack_0 : boolean;
  signal simple_obj_ref_823_inst_req_0 : boolean;
  signal simple_obj_ref_823_inst_ack_0 : boolean;
  signal ptr_deref_827_base_resize_req_0 : boolean;
  signal ptr_deref_827_base_resize_ack_0 : boolean;
  signal ptr_deref_827_root_address_inst_req_0 : boolean;
  signal ptr_deref_827_root_address_inst_ack_0 : boolean;
  signal ptr_deref_827_addr_0_req_0 : boolean;
  signal ptr_deref_827_addr_0_ack_0 : boolean;
  signal ptr_deref_827_gather_scatter_req_0 : boolean;
  signal ptr_deref_827_gather_scatter_ack_0 : boolean;
  signal ptr_deref_827_store_0_req_0 : boolean;
  signal ptr_deref_827_store_0_ack_0 : boolean;
  signal ptr_deref_827_store_0_req_1 : boolean;
  signal ptr_deref_827_store_0_ack_1 : boolean;
  signal binary_834_inst_req_0 : boolean;
  signal binary_834_inst_ack_0 : boolean;
  signal binary_834_inst_req_1 : boolean;
  signal binary_834_inst_ack_1 : boolean;
  signal binary_840_inst_req_0 : boolean;
  signal binary_840_inst_ack_0 : boolean;
  signal binary_840_inst_req_1 : boolean;
  signal binary_840_inst_ack_1 : boolean;
  signal do_while_stmt_398_branch_req_0 : boolean;
  signal unary_844_inst_req_0 : boolean;
  signal unary_844_inst_ack_0 : boolean;
  signal unary_844_inst_req_1 : boolean;
  signal unary_844_inst_ack_1 : boolean;
  signal do_while_stmt_398_branch_ack_0 : boolean;
  signal do_while_stmt_398_branch_ack_1 : boolean;
  signal phi_stmt_392_req_0 : boolean;
  signal phi_stmt_392_ack_0 : boolean;
  signal global_clock_cycle_count: integer := 0;
  -- 
begin --  
  ---------------------------------------------------------- 
  process(clk)  
  begin -- 
    if(clk'event and clk = '1') then -- 
      if(reset = '1') then -- 
        global_clock_cycle_count <= 0; --
      else -- 
        global_clock_cycle_count <= global_clock_cycle_count + 1; -- 
      end if; --
    end if; --
  end process;
  ---------------------------------------------------------- 
  -- output port buffering assignments
  -- level-to-pulse translation..
  l2pStart: level_to_pulse -- 
    generic map (forward_delay => 0, backward_delay => 0) 
    port map(clk => clk, reset =>reset, lreq => start_req, lack => start_ack_sig, preq => start_req_symbol, pack => start_ack_symbol); -- 
  start_ack <= start_ack_sig; 
  l2pFin: level_to_pulse -- 
    generic map (forward_delay => 0, backward_delay => 0) 
    port map(clk => clk, reset =>reset, lreq => fin_req, lack => fin_ack_sig, preq => fin_req_symbol, pack => fin_ack_symbol); -- 
  fin_ack <= fin_ack_sig; 
  tag_push <= '1' when start_req_symbol else '0'; 
  tag_pop  <= fin_req and fin_ack_sig ; 
  LogCPEvent(clk,reset,global_clock_cycle_count, start_req_symbol,"x_vectorSum_x start_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  start_ack_symbol,"x_vectorSum_x start_ack symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_req_symbol,"x_vectorSum_x fin_req symbol");
  LogCPEvent(clk,reset,global_clock_cycle_count,  fin_ack_symbol,"x_vectorSum_x fin_ack symbol");
  tagQueue: QueueBase generic map(data_width => 2, queue_depth => 2 ) -- 
    port map(pop_req => tag_pop, pop_ack => open, 
    push_req => tag_push, push_ack => open, 
    data_out => tag_out, data_in => tag_in, 
    clk => clk, reset => reset); -- 
  -- the control path
  always_true_symbol <= true; 
  x_vectorSum_x_xCP_1292: Block -- control-path 
    signal cp_elements: BooleanArray(1181 downto 0);
    -- 
  begin -- 
    cp_elements(0) <= start_req_symbol;
    start_ack_symbol <= cp_elements(1180);
    finAckJoin: join2 
    port map(pred0 => fin_req_symbol, pred1 =>cp_elements(1180), symbol_out => fin_ack_symbol, clk => clk, reset => reset);
    -- CP-element group 0 transition  place  output  bypass 
    -- predecessors 
    -- successors 1181 
    -- members (13) 
      -- 	$entry
      -- 	branch_block_stmt_389/$entry
      -- 	branch_block_stmt_389/branch_block_stmt_389__entry__
      -- 	branch_block_stmt_389/bbx_xnph_bb_1
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/$entry
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/$exit
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/phi_stmt_392/$entry
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/phi_stmt_392/$exit
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/phi_stmt_392/phi_stmt_392_sources/$entry
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/phi_stmt_392/phi_stmt_392_sources/$exit
      -- 	branch_block_stmt_389/bbx_xnph_bb_1_PhiReq/phi_stmt_392/phi_stmt_392_req
      -- 	branch_block_stmt_389/merge_stmt_391_PhiReqMerge
      -- 	branch_block_stmt_389/merge_stmt_391_PhiAck/$entry
      -- 
    phi_stmt_392_req_4478_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(0), ack => phi_stmt_392_req_0); -- 
    -- CP-element group 1 merge  place  bypass 
    -- predecessors 
    -- successors 1180 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398__exit__
      -- 
    -- Element group cp_elements(1) is bound as output of CP function.
    -- CP-element group 2 merge  place  bypass 
    -- predecessors 
    -- successors 5 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_back
      -- 
    -- Element group cp_elements(2) is bound as output of CP function.
    -- CP-element group 3 branch  place  bypass 
    -- predecessors 1165 
    -- successors 1176 1178 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/condition_done
      -- 
    cp_elements(3) <= cp_elements(1165);
    -- CP-element group 4 branch  place  bypass 
    -- predecessors 1175 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_body_done
      -- 
    cp_elements(4) <= cp_elements(1175);
    -- CP-element group 5 fork  transition  bypass 
    -- predecessors 2 
    -- successors 10 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/back_edge_to_loop_body
      -- 
    cp_elements(5) <= cp_elements(2);
    -- CP-element group 6 fork  transition  bypass 
    -- predecessors 1181 
    -- successors 13 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/first_time_through_loop_body
      -- 
    cp_elements(6) <= cp_elements(1181);
    -- CP-element group 7 join  fork  transition  bypass 
    -- predecessors 
    -- successors 341 19 45 63 81 99 110 128 146 164 175 370 388 305 877 1143 791 489 507 525 834 705 748 1154 1164 323 359 22 23 34 576 619 662 406 424 435 453 471 193 211 229 240 258 276 294 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/loop_body_start
      -- 
    -- Element group cp_elements(7) is bound as output of CP function.
    -- CP-element group 8 join  transition  bypass 
    -- predecessors 
    -- successors 9 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_req_0_raw
      -- 
    -- Element group cp_elements(8) is bound as output of CP function.
    -- CP-element group 9 transition  output  bypass 
    -- predecessors 8 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_req_0
      -- 
    cp_elements(9) <= cp_elements(8);
    phi_stmt_400_req_0_1324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(9), ack => phi_stmt_400_req_0); -- 
    -- CP-element group 10 fork  transition  bypass 
    -- predecessors 5 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_trigger_from_back_edge_to_loop_body
      -- 
    cp_elements(10) <= cp_elements(5);
    -- CP-element group 11 join  transition  bypass 
    -- predecessors 
    -- successors 12 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_req_1_raw
      -- 
    -- Element group cp_elements(11) is bound as output of CP function.
    -- CP-element group 12 transition  output  bypass 
    -- predecessors 11 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_req_1
      -- 
    cp_elements(12) <= cp_elements(11);
    phi_stmt_400_req_1_1327_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(12), ack => phi_stmt_400_req_1); -- 
    -- CP-element group 13 fork  transition  bypass 
    -- predecessors 6 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_trigger_from_first_time_through_loop_body
      -- 
    cp_elements(13) <= cp_elements(6);
    -- CP-element group 14 join  transition  bypass 
    -- predecessors 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_phi_sequencer_reqs_merged
      -- 
    -- Element group cp_elements(14) is bound as output of CP function.
    -- CP-element group 15 join  fork  transition  bypass 
    -- predecessors 
    -- successors 1149 29 
    -- marked successors 18 22 
    -- members (3) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_phi_sequencer_done
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_completed_
      -- 
    -- Element group cp_elements(15) is bound as output of CP function.
    -- CP-element group 16 transition  input  bypass 
    -- predecessors 
    -- successors 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_ack
      -- 
    phi_stmt_400_ack_1331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_400_ack_0, ack => cp_elements(16)); -- 
    -- CP-element group 17 join  fork  transition  bypass 
    -- predecessors 18 22 
    -- marked predecessors 1146 26 
    -- successors 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_enable_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/phi_stmt_400_trigger_
      -- 
    cpelement_group_17 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(18);
      predecessors(1) <= cp_elements(22);
      marked_predecessors(0) <= cp_elements(1146);
      marked_predecessors(1) <= cp_elements(26);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(17)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(17),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 18 join  transition  bypass 
    -- predecessors 21 
    -- marked predecessors 15 
    -- successors 17 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_completed_
      -- 
    cpelement_group_18 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(21);
      marked_predecessors(0) <= cp_elements(15);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(18)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(18),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 19 join  transition  bypass 
    -- predecessors 7 
    -- marked predecessors 1144 
    -- successors 20 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_402_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_402_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_402_completed_
      -- 
    cpelement_group_19 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(7);
      marked_predecessors(0) <= cp_elements(1144);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(19)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(19),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 20 transition  output  bypass 
    -- predecessors 19 
    -- successors 21 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_complete/req
      -- 
    cp_elements(20) <= cp_elements(19);
    req_1347_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(20), ack => type_cast_403_inst_req_0); -- 
    -- CP-element group 21 transition  input  bypass 
    -- predecessors 20 
    -- successors 18 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/type_cast_403_complete/ack
      -- 
    ack_1348_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_403_inst_ack_0, ack => cp_elements(21)); -- 
    -- CP-element group 22 join  transition  bypass 
    -- predecessors 7 
    -- marked predecessors 15 
    -- successors 17 
    -- members (3) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_404_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_404_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_404_completed_
      -- 
    cpelement_group_22 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(7);
      marked_predecessors(0) <= cp_elements(15);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(22)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(22),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 23 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_active_
      -- 
    cp_elements(23) <= cp_elements(7);
    -- CP-element group 24 join  fork  transition  bypass 
    -- predecessors 26 28 
    -- successors 40 105 170 496 514 532 365 430 235 300 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_411_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_411_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_411_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_completed_
      -- 
    cpelement_group_24 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(26);
      predecessors(1) <= cp_elements(28);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(24)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(24),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 25 join  transition  bypass 
    -- predecessors 29 
    -- marked predecessors 26 
    -- successors 30 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_sample_start_
      -- 
    cpelement_group_25 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(29);
      marked_predecessors(0) <= cp_elements(26);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(25)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(25),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 26 fork  transition  bypass 
    -- predecessors 31 
    -- successors 24 
    -- marked successors 17 25 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_sample_completed_
      -- 
    cp_elements(26) <= cp_elements(31);
    -- CP-element group 27 join  transition  bypass 
    -- predecessors 29 
    -- marked predecessors 37 102 167 491 509 527 362 427 232 297 
    -- successors 32 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_update_start_
      -- 
    cpelement_group_27 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(9 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(29);
      marked_predecessors(0) <= cp_elements(37);
      marked_predecessors(1) <= cp_elements(102);
      marked_predecessors(2) <= cp_elements(167);
      marked_predecessors(3) <= cp_elements(491);
      marked_predecessors(4) <= cp_elements(509);
      marked_predecessors(5) <= cp_elements(527);
      marked_predecessors(6) <= cp_elements(362);
      marked_predecessors(7) <= cp_elements(427);
      marked_predecessors(8) <= cp_elements(232);
      marked_predecessors(9) <= cp_elements(297);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(27)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(27),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 28 transition  bypass 
    -- predecessors 33 
    -- successors 24 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_update_completed_
      -- 
    cp_elements(28) <= cp_elements(33);
    -- CP-element group 29 fork  transition  bypass 
    -- predecessors 15 
    -- successors 25 27 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_407_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_407_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_407_completed_
      -- 
    cp_elements(29) <= cp_elements(15);
    -- CP-element group 30 transition  output  bypass 
    -- predecessors 25 
    -- successors 31 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Sample/rr
      -- 
    cp_elements(30) <= cp_elements(25);
    rr_1368_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(30), ack => binary_410_inst_req_0); -- 
    -- CP-element group 31 transition  input  bypass 
    -- predecessors 30 
    -- successors 26 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Sample/ra
      -- 
    ra_1369_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_410_inst_ack_0, ack => cp_elements(31)); -- 
    -- CP-element group 32 transition  output  bypass 
    -- predecessors 27 
    -- successors 33 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Update/cr
      -- 
    cp_elements(32) <= cp_elements(27);
    cr_1373_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(32), ack => binary_410_inst_req_1); -- 
    -- CP-element group 33 transition  input  bypass 
    -- predecessors 32 
    -- successors 28 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_410_Update/ca
      -- 
    ca_1374_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_410_inst_ack_1, ack => cp_elements(33)); -- 
    -- CP-element group 34 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_active_
      -- 
    cp_elements(34) <= cp_elements(7);
    -- CP-element group 35 join  fork  transition  bypass 
    -- predecessors 37 39 
    -- successors 52 70 88 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_417_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_417_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_417_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_completed_
      -- 
    cpelement_group_35 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(37);
      predecessors(1) <= cp_elements(39);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(35)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(35),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 36 join  transition  bypass 
    -- predecessors 40 
    -- marked predecessors 37 
    -- successors 41 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_sample_start_
      -- 
    cpelement_group_36 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(40);
      marked_predecessors(0) <= cp_elements(37);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(36)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(36),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 37 fork  transition  bypass 
    -- predecessors 42 
    -- successors 35 
    -- marked successors 36 27 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_sample_completed_
      -- 
    cp_elements(37) <= cp_elements(42);
    -- CP-element group 38 join  transition  bypass 
    -- predecessors 40 
    -- marked predecessors 47 65 83 
    -- successors 43 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_update_start_
      -- 
    cpelement_group_38 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(40);
      marked_predecessors(0) <= cp_elements(47);
      marked_predecessors(1) <= cp_elements(65);
      marked_predecessors(2) <= cp_elements(83);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(38)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(38),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 39 transition  bypass 
    -- predecessors 44 
    -- successors 35 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_update_completed_
      -- 
    cp_elements(39) <= cp_elements(44);
    -- CP-element group 40 fork  transition  bypass 
    -- predecessors 24 
    -- successors 36 38 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_413_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_413_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_413_completed_
      -- 
    cp_elements(40) <= cp_elements(24);
    -- CP-element group 41 transition  output  bypass 
    -- predecessors 36 
    -- successors 42 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Sample/rr
      -- 
    cp_elements(41) <= cp_elements(36);
    rr_1391_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(41), ack => binary_416_inst_req_0); -- 
    -- CP-element group 42 transition  input  bypass 
    -- predecessors 41 
    -- successors 37 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Sample/ra
      -- 
    ra_1392_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_416_inst_ack_0, ack => cp_elements(42)); -- 
    -- CP-element group 43 transition  output  bypass 
    -- predecessors 38 
    -- successors 44 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Update/cr
      -- 
    cp_elements(43) <= cp_elements(38);
    cr_1396_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(43), ack => binary_416_inst_req_1); -- 
    -- CP-element group 44 transition  input  bypass 
    -- predecessors 43 
    -- successors 39 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_416_Update/ca
      -- 
    ca_1397_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_416_inst_ack_1, ack => cp_elements(44)); -- 
    -- CP-element group 45 transition  bypass 
    -- predecessors 7 
    -- successors 46 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_trigger_
      -- 
    cp_elements(45) <= cp_elements(7);
    -- CP-element group 46 join  transition  bypass 
    -- predecessors 45 48 
    -- marked predecessors 1111 
    -- successors 61 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_active_
      -- 
    cpelement_group_46 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(45);
      predecessors(1) <= cp_elements(48);
      marked_predecessors(0) <= cp_elements(1111);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(46)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(46),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 47 join  fork  transition  bypass 
    -- predecessors 62 
    -- marked predecessors 1114 
    -- successors 1112 
    -- marked successors 38 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_422_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_422_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_422_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_812_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_812_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_812_completed_
      -- 
    cpelement_group_47 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(62);
      marked_predecessors(0) <= cp_elements(1114);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(47)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(47),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 48 transition  bypass 
    -- predecessors 60 
    -- successors 46 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_root_address_calculated
      -- 
    cp_elements(48) <= cp_elements(60);
    -- CP-element group 49 transition  bypass 
    -- predecessors 56 
    -- successors 57 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_indices_scaled
      -- 
    cp_elements(49) <= cp_elements(56);
    -- CP-element group 50 transition  bypass 
    -- predecessors 58 
    -- successors 59 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_offset_calculated
      -- 
    cp_elements(50) <= cp_elements(58);
    -- CP-element group 51 transition  bypass 
    -- predecessors 54 
    -- successors 55 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_resized_0
      -- 
    cp_elements(51) <= cp_elements(54);
    -- CP-element group 52 transition  bypass 
    -- predecessors 35 
    -- successors 53 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_419_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_419_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_419_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_computed_0
      -- 
    cp_elements(52) <= cp_elements(35);
    -- CP-element group 53 transition  output  bypass 
    -- predecessors 52 
    -- successors 54 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_resize_0/index_resize_req
      -- 
    cp_elements(53) <= cp_elements(52);
    index_resize_req_1415_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(53), ack => array_obj_ref_420_index_0_resize_req_0); -- 
    -- CP-element group 54 transition  input  bypass 
    -- predecessors 53 
    -- successors 51 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_resize_0/$exit
      -- 
    index_resize_ack_1416_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_420_index_0_resize_ack_0, ack => cp_elements(54)); -- 
    -- CP-element group 55 transition  output  bypass 
    -- predecessors 51 
    -- successors 56 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_scale_0/$entry
      -- 
    cp_elements(55) <= cp_elements(51);
    scale_rename_req_1420_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(55), ack => array_obj_ref_420_index_0_rename_req_0); -- 
    -- CP-element group 56 transition  input  bypass 
    -- predecessors 55 
    -- successors 49 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1421_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_420_index_0_rename_ack_0, ack => cp_elements(56)); -- 
    -- CP-element group 57 transition  output  bypass 
    -- predecessors 49 
    -- successors 58 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_add_indices/$entry
      -- 
    cp_elements(57) <= cp_elements(49);
    final_index_req_1425_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(57), ack => array_obj_ref_420_offset_inst_req_0); -- 
    -- CP-element group 58 transition  input  bypass 
    -- predecessors 57 
    -- successors 50 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_add_indices/final_index_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_add_indices/$exit
      -- 
    final_index_ack_1426_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_420_offset_inst_ack_0, ack => cp_elements(58)); -- 
    -- CP-element group 59 transition  output  bypass 
    -- predecessors 50 
    -- successors 60 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_base_plus_offset/sum_rename_req
      -- 
    cp_elements(59) <= cp_elements(50);
    sum_rename_req_1430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(59), ack => array_obj_ref_420_root_address_inst_req_0); -- 
    -- CP-element group 60 transition  input  bypass 
    -- predecessors 59 
    -- successors 48 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_420_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_420_root_address_inst_ack_0, ack => cp_elements(60)); -- 
    -- CP-element group 61 transition  output  bypass 
    -- predecessors 46 
    -- successors 62 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_complete/final_reg_req
      -- 
    cp_elements(61) <= cp_elements(46);
    final_reg_req_1435_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(61), ack => addr_of_421_final_reg_req_0); -- 
    -- CP-element group 62 transition  input  bypass 
    -- predecessors 61 
    -- successors 47 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_421_complete/final_reg_ack
      -- 
    final_reg_ack_1436_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_421_final_reg_ack_0, ack => cp_elements(62)); -- 
    -- CP-element group 63 transition  bypass 
    -- predecessors 7 
    -- successors 64 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_trigger_
      -- 
    cp_elements(63) <= cp_elements(7);
    -- CP-element group 64 join  transition  bypass 
    -- predecessors 63 66 
    -- marked predecessors 860 
    -- successors 79 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_active_
      -- 
    cpelement_group_64 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(63);
      predecessors(1) <= cp_elements(66);
      marked_predecessors(0) <= cp_elements(860);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(64)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(64),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 65 fork  transition  bypass 
    -- predecessors 80 
    -- successors 865 
    -- marked successors 38 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_427_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_427_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_427_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_670_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_670_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_670_completed_
      -- 
    cp_elements(65) <= cp_elements(80);
    -- CP-element group 66 transition  bypass 
    -- predecessors 78 
    -- successors 64 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_root_address_calculated
      -- 
    cp_elements(66) <= cp_elements(78);
    -- CP-element group 67 transition  bypass 
    -- predecessors 74 
    -- successors 75 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_indices_scaled
      -- 
    cp_elements(67) <= cp_elements(74);
    -- CP-element group 68 transition  bypass 
    -- predecessors 76 
    -- successors 77 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_offset_calculated
      -- 
    cp_elements(68) <= cp_elements(76);
    -- CP-element group 69 transition  bypass 
    -- predecessors 72 
    -- successors 73 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_resized_0
      -- 
    cp_elements(69) <= cp_elements(72);
    -- CP-element group 70 transition  bypass 
    -- predecessors 35 
    -- successors 71 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_424_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_424_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_424_completed_
      -- 
    cp_elements(70) <= cp_elements(35);
    -- CP-element group 71 transition  output  bypass 
    -- predecessors 70 
    -- successors 72 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_resize_0/index_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_resize_0/$entry
      -- 
    cp_elements(71) <= cp_elements(70);
    index_resize_req_1454_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(71), ack => array_obj_ref_425_index_0_resize_req_0); -- 
    -- CP-element group 72 transition  input  bypass 
    -- predecessors 71 
    -- successors 69 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_resize_0/$exit
      -- 
    index_resize_ack_1455_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_425_index_0_resize_ack_0, ack => cp_elements(72)); -- 
    -- CP-element group 73 transition  output  bypass 
    -- predecessors 69 
    -- successors 74 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_scale_0/scale_rename_req
      -- 
    cp_elements(73) <= cp_elements(69);
    scale_rename_req_1459_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(73), ack => array_obj_ref_425_index_0_rename_req_0); -- 
    -- CP-element group 74 transition  input  bypass 
    -- predecessors 73 
    -- successors 67 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_index_scale_0/$exit
      -- 
    scale_rename_ack_1460_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_425_index_0_rename_ack_0, ack => cp_elements(74)); -- 
    -- CP-element group 75 transition  output  bypass 
    -- predecessors 67 
    -- successors 76 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_add_indices/final_index_req
      -- 
    cp_elements(75) <= cp_elements(67);
    final_index_req_1464_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(75), ack => array_obj_ref_425_offset_inst_req_0); -- 
    -- CP-element group 76 transition  input  bypass 
    -- predecessors 75 
    -- successors 68 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_add_indices/final_index_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_add_indices/$exit
      -- 
    final_index_ack_1465_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_425_offset_inst_ack_0, ack => cp_elements(76)); -- 
    -- CP-element group 77 transition  output  bypass 
    -- predecessors 68 
    -- successors 78 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_base_plus_offset/$entry
      -- 
    cp_elements(77) <= cp_elements(68);
    sum_rename_req_1469_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(77), ack => array_obj_ref_425_root_address_inst_req_0); -- 
    -- CP-element group 78 transition  input  bypass 
    -- predecessors 77 
    -- successors 66 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_425_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1470_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_425_root_address_inst_ack_0, ack => cp_elements(78)); -- 
    -- CP-element group 79 transition  output  bypass 
    -- predecessors 64 
    -- successors 80 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_complete/final_reg_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_complete/$entry
      -- 
    cp_elements(79) <= cp_elements(64);
    final_reg_req_1474_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(79), ack => addr_of_426_final_reg_req_0); -- 
    -- CP-element group 80 transition  input  bypass 
    -- predecessors 79 
    -- successors 65 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_426_complete/final_reg_ack
      -- 
    final_reg_ack_1475_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_426_final_reg_ack_0, ack => cp_elements(80)); -- 
    -- CP-element group 81 transition  bypass 
    -- predecessors 7 
    -- successors 82 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_trigger_
      -- 
    cp_elements(81) <= cp_elements(7);
    -- CP-element group 82 join  transition  bypass 
    -- predecessors 81 84 
    -- marked predecessors 844 
    -- successors 97 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_active_
      -- 
    cpelement_group_82 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(81);
      predecessors(1) <= cp_elements(84);
      marked_predecessors(0) <= cp_elements(844);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(82)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(82),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 83 fork  transition  bypass 
    -- predecessors 98 
    -- successors 849 
    -- marked successors 38 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_432_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_432_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_432_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_666_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_666_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_666_completed_
      -- 
    cp_elements(83) <= cp_elements(98);
    -- CP-element group 84 transition  bypass 
    -- predecessors 96 
    -- successors 82 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_root_address_calculated
      -- 
    cp_elements(84) <= cp_elements(96);
    -- CP-element group 85 transition  bypass 
    -- predecessors 92 
    -- successors 93 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_indices_scaled
      -- 
    cp_elements(85) <= cp_elements(92);
    -- CP-element group 86 transition  bypass 
    -- predecessors 94 
    -- successors 95 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_offset_calculated
      -- 
    cp_elements(86) <= cp_elements(94);
    -- CP-element group 87 transition  bypass 
    -- predecessors 90 
    -- successors 91 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_resized_0
      -- 
    cp_elements(87) <= cp_elements(90);
    -- CP-element group 88 transition  bypass 
    -- predecessors 35 
    -- successors 89 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_429_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_429_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_429_completed_
      -- 
    cp_elements(88) <= cp_elements(35);
    -- CP-element group 89 transition  output  bypass 
    -- predecessors 88 
    -- successors 90 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_resize_0/index_resize_req
      -- 
    cp_elements(89) <= cp_elements(88);
    index_resize_req_1493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(89), ack => array_obj_ref_430_index_0_resize_req_0); -- 
    -- CP-element group 90 transition  input  bypass 
    -- predecessors 89 
    -- successors 87 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_0_resize_ack_0, ack => cp_elements(90)); -- 
    -- CP-element group 91 transition  output  bypass 
    -- predecessors 87 
    -- successors 92 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_scale_0/scale_rename_req
      -- 
    cp_elements(91) <= cp_elements(87);
    scale_rename_req_1498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(91), ack => array_obj_ref_430_index_0_rename_req_0); -- 
    -- CP-element group 92 transition  input  bypass 
    -- predecessors 91 
    -- successors 85 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_index_0_rename_ack_0, ack => cp_elements(92)); -- 
    -- CP-element group 93 transition  output  bypass 
    -- predecessors 85 
    -- successors 94 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_add_indices/$entry
      -- 
    cp_elements(93) <= cp_elements(85);
    final_index_req_1503_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(93), ack => array_obj_ref_430_offset_inst_req_0); -- 
    -- CP-element group 94 transition  input  bypass 
    -- predecessors 93 
    -- successors 86 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_add_indices/final_index_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_add_indices/$exit
      -- 
    final_index_ack_1504_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_offset_inst_ack_0, ack => cp_elements(94)); -- 
    -- CP-element group 95 transition  output  bypass 
    -- predecessors 86 
    -- successors 96 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_base_plus_offset/$entry
      -- 
    cp_elements(95) <= cp_elements(86);
    sum_rename_req_1508_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(95), ack => array_obj_ref_430_root_address_inst_req_0); -- 
    -- CP-element group 96 transition  input  bypass 
    -- predecessors 95 
    -- successors 84 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_430_base_plus_offset/$exit
      -- 
    sum_rename_ack_1509_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_430_root_address_inst_ack_0, ack => cp_elements(96)); -- 
    -- CP-element group 97 transition  output  bypass 
    -- predecessors 82 
    -- successors 98 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_complete/final_reg_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_complete/$entry
      -- 
    cp_elements(97) <= cp_elements(82);
    final_reg_req_1513_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(97), ack => addr_of_431_final_reg_req_0); -- 
    -- CP-element group 98 transition  input  bypass 
    -- predecessors 97 
    -- successors 83 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_431_complete/final_reg_ack
      -- 
    final_reg_ack_1514_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_431_final_reg_ack_0, ack => cp_elements(98)); -- 
    -- CP-element group 99 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_active_
      -- 
    cp_elements(99) <= cp_elements(7);
    -- CP-element group 100 join  fork  transition  bypass 
    -- predecessors 102 104 
    -- successors 117 135 153 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_438_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_438_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_438_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_completed_
      -- 
    cpelement_group_100 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(102);
      predecessors(1) <= cp_elements(104);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(100)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(100),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 101 join  transition  bypass 
    -- predecessors 105 
    -- marked predecessors 102 
    -- successors 106 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_sample_start_
      -- 
    cpelement_group_101 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(105);
      marked_predecessors(0) <= cp_elements(102);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(101)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(101),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 102 fork  transition  bypass 
    -- predecessors 107 
    -- successors 100 
    -- marked successors 101 27 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_sample_completed_
      -- 
    cp_elements(102) <= cp_elements(107);
    -- CP-element group 103 join  transition  bypass 
    -- predecessors 105 
    -- marked predecessors 112 130 148 
    -- successors 108 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_update_start_
      -- 
    cpelement_group_103 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(105);
      marked_predecessors(0) <= cp_elements(112);
      marked_predecessors(1) <= cp_elements(130);
      marked_predecessors(2) <= cp_elements(148);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(103)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(103),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 104 transition  bypass 
    -- predecessors 109 
    -- successors 100 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_update_completed_
      -- 
    cp_elements(104) <= cp_elements(109);
    -- CP-element group 105 fork  transition  bypass 
    -- predecessors 24 
    -- successors 101 103 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_434_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_434_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_434_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_trigger_
      -- 
    cp_elements(105) <= cp_elements(24);
    -- CP-element group 106 transition  output  bypass 
    -- predecessors 101 
    -- successors 107 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Sample/rr
      -- 
    cp_elements(106) <= cp_elements(101);
    rr_1531_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(106), ack => binary_437_inst_req_0); -- 
    -- CP-element group 107 transition  input  bypass 
    -- predecessors 106 
    -- successors 102 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Sample/ra
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Sample/$exit
      -- 
    ra_1532_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_437_inst_ack_0, ack => cp_elements(107)); -- 
    -- CP-element group 108 transition  output  bypass 
    -- predecessors 103 
    -- successors 109 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Update/cr
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Update/$entry
      -- 
    cp_elements(108) <= cp_elements(103);
    cr_1536_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(108), ack => binary_437_inst_req_1); -- 
    -- CP-element group 109 transition  input  bypass 
    -- predecessors 108 
    -- successors 104 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Update/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_437_Update/$exit
      -- 
    ca_1537_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_437_inst_ack_1, ack => cp_elements(109)); -- 
    -- CP-element group 110 transition  bypass 
    -- predecessors 7 
    -- successors 111 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_trigger_
      -- 
    cp_elements(110) <= cp_elements(7);
    -- CP-element group 111 join  transition  bypass 
    -- predecessors 110 113 
    -- marked predecessors 1079 
    -- successors 126 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_active_
      -- 
    cpelement_group_111 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(110);
      predecessors(1) <= cp_elements(113);
      marked_predecessors(0) <= cp_elements(1079);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(111)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 112 join  fork  transition  bypass 
    -- predecessors 127 
    -- marked predecessors 1082 
    -- successors 1080 
    -- marked successors 103 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_443_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_443_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_443_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_793_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_793_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_793_completed_
      -- 
    cpelement_group_112 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(127);
      marked_predecessors(0) <= cp_elements(1082);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(112)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(112),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 113 transition  bypass 
    -- predecessors 125 
    -- successors 111 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_root_address_calculated
      -- 
    cp_elements(113) <= cp_elements(125);
    -- CP-element group 114 transition  bypass 
    -- predecessors 121 
    -- successors 122 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_indices_scaled
      -- 
    cp_elements(114) <= cp_elements(121);
    -- CP-element group 115 transition  bypass 
    -- predecessors 123 
    -- successors 124 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_offset_calculated
      -- 
    cp_elements(115) <= cp_elements(123);
    -- CP-element group 116 transition  bypass 
    -- predecessors 119 
    -- successors 120 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_resized_0
      -- 
    cp_elements(116) <= cp_elements(119);
    -- CP-element group 117 transition  bypass 
    -- predecessors 100 
    -- successors 118 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_440_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_440_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_440_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_computed_0
      -- 
    cp_elements(117) <= cp_elements(100);
    -- CP-element group 118 transition  output  bypass 
    -- predecessors 117 
    -- successors 119 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_resize_0/index_resize_req
      -- 
    cp_elements(118) <= cp_elements(117);
    index_resize_req_1555_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(118), ack => array_obj_ref_441_index_0_resize_req_0); -- 
    -- CP-element group 119 transition  input  bypass 
    -- predecessors 118 
    -- successors 116 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1556_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_441_index_0_resize_ack_0, ack => cp_elements(119)); -- 
    -- CP-element group 120 transition  output  bypass 
    -- predecessors 116 
    -- successors 121 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_scale_0/scale_rename_req
      -- 
    cp_elements(120) <= cp_elements(116);
    scale_rename_req_1560_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(120), ack => array_obj_ref_441_index_0_rename_req_0); -- 
    -- CP-element group 121 transition  input  bypass 
    -- predecessors 120 
    -- successors 114 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1561_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_441_index_0_rename_ack_0, ack => cp_elements(121)); -- 
    -- CP-element group 122 transition  output  bypass 
    -- predecessors 114 
    -- successors 123 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_add_indices/final_index_req
      -- 
    cp_elements(122) <= cp_elements(114);
    final_index_req_1565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(122), ack => array_obj_ref_441_offset_inst_req_0); -- 
    -- CP-element group 123 transition  input  bypass 
    -- predecessors 122 
    -- successors 115 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_add_indices/final_index_ack
      -- 
    final_index_ack_1566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_441_offset_inst_ack_0, ack => cp_elements(123)); -- 
    -- CP-element group 124 transition  output  bypass 
    -- predecessors 115 
    -- successors 125 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_base_plus_offset/sum_rename_req
      -- 
    cp_elements(124) <= cp_elements(115);
    sum_rename_req_1570_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(124), ack => array_obj_ref_441_root_address_inst_req_0); -- 
    -- CP-element group 125 transition  input  bypass 
    -- predecessors 124 
    -- successors 113 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_441_base_plus_offset/$exit
      -- 
    sum_rename_ack_1571_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_441_root_address_inst_ack_0, ack => cp_elements(125)); -- 
    -- CP-element group 126 transition  output  bypass 
    -- predecessors 111 
    -- successors 127 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_complete/final_reg_req
      -- 
    cp_elements(126) <= cp_elements(111);
    final_reg_req_1575_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(126), ack => addr_of_442_final_reg_req_0); -- 
    -- CP-element group 127 transition  input  bypass 
    -- predecessors 126 
    -- successors 112 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_442_complete/final_reg_ack
      -- 
    final_reg_ack_1576_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_442_final_reg_ack_0, ack => cp_elements(127)); -- 
    -- CP-element group 128 transition  bypass 
    -- predecessors 7 
    -- successors 129 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_trigger_
      -- 
    cp_elements(128) <= cp_elements(7);
    -- CP-element group 129 join  transition  bypass 
    -- predecessors 128 131 
    -- marked predecessors 817 
    -- successors 144 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_active_
      -- 
    cpelement_group_129 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(128);
      predecessors(1) <= cp_elements(131);
      marked_predecessors(0) <= cp_elements(817);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(129)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(129),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 130 fork  transition  bypass 
    -- predecessors 145 
    -- successors 822 
    -- marked successors 103 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_448_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_448_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_448_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_657_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_657_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_657_completed_
      -- 
    cp_elements(130) <= cp_elements(145);
    -- CP-element group 131 transition  bypass 
    -- predecessors 143 
    -- successors 129 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_root_address_calculated
      -- 
    cp_elements(131) <= cp_elements(143);
    -- CP-element group 132 transition  bypass 
    -- predecessors 139 
    -- successors 140 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_indices_scaled
      -- 
    cp_elements(132) <= cp_elements(139);
    -- CP-element group 133 transition  bypass 
    -- predecessors 141 
    -- successors 142 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_offset_calculated
      -- 
    cp_elements(133) <= cp_elements(141);
    -- CP-element group 134 transition  bypass 
    -- predecessors 137 
    -- successors 138 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_resized_0
      -- 
    cp_elements(134) <= cp_elements(137);
    -- CP-element group 135 transition  bypass 
    -- predecessors 100 
    -- successors 136 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_445_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_445_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_445_completed_
      -- 
    cp_elements(135) <= cp_elements(100);
    -- CP-element group 136 transition  output  bypass 
    -- predecessors 135 
    -- successors 137 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_resize_0/index_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_resize_0/$entry
      -- 
    cp_elements(136) <= cp_elements(135);
    index_resize_req_1594_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(136), ack => array_obj_ref_446_index_0_resize_req_0); -- 
    -- CP-element group 137 transition  input  bypass 
    -- predecessors 136 
    -- successors 134 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_resize_0/$exit
      -- 
    index_resize_ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_446_index_0_resize_ack_0, ack => cp_elements(137)); -- 
    -- CP-element group 138 transition  output  bypass 
    -- predecessors 134 
    -- successors 139 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_scale_0/$entry
      -- 
    cp_elements(138) <= cp_elements(134);
    scale_rename_req_1599_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(138), ack => array_obj_ref_446_index_0_rename_req_0); -- 
    -- CP-element group 139 transition  input  bypass 
    -- predecessors 138 
    -- successors 132 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_index_scale_0/$exit
      -- 
    scale_rename_ack_1600_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_446_index_0_rename_ack_0, ack => cp_elements(139)); -- 
    -- CP-element group 140 transition  output  bypass 
    -- predecessors 132 
    -- successors 141 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_add_indices/final_index_req
      -- 
    cp_elements(140) <= cp_elements(132);
    final_index_req_1604_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(140), ack => array_obj_ref_446_offset_inst_req_0); -- 
    -- CP-element group 141 transition  input  bypass 
    -- predecessors 140 
    -- successors 133 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_add_indices/final_index_ack
      -- 
    final_index_ack_1605_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_446_offset_inst_ack_0, ack => cp_elements(141)); -- 
    -- CP-element group 142 transition  output  bypass 
    -- predecessors 133 
    -- successors 143 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_base_plus_offset/$entry
      -- 
    cp_elements(142) <= cp_elements(133);
    sum_rename_req_1609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(142), ack => array_obj_ref_446_root_address_inst_req_0); -- 
    -- CP-element group 143 transition  input  bypass 
    -- predecessors 142 
    -- successors 131 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_446_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_446_root_address_inst_ack_0, ack => cp_elements(143)); -- 
    -- CP-element group 144 transition  output  bypass 
    -- predecessors 129 
    -- successors 145 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_complete/final_reg_req
      -- 
    cp_elements(144) <= cp_elements(129);
    final_reg_req_1614_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(144), ack => addr_of_447_final_reg_req_0); -- 
    -- CP-element group 145 transition  input  bypass 
    -- predecessors 144 
    -- successors 130 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_447_complete/final_reg_ack
      -- 
    final_reg_ack_1615_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_447_final_reg_ack_0, ack => cp_elements(145)); -- 
    -- CP-element group 146 transition  bypass 
    -- predecessors 7 
    -- successors 147 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_trigger_
      -- 
    cp_elements(146) <= cp_elements(7);
    -- CP-element group 147 join  transition  bypass 
    -- predecessors 146 149 
    -- marked predecessors 801 
    -- successors 162 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_active_
      -- 
    cpelement_group_147 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(146);
      predecessors(1) <= cp_elements(149);
      marked_predecessors(0) <= cp_elements(801);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(147)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 148 fork  transition  bypass 
    -- predecessors 163 
    -- successors 806 
    -- marked successors 103 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_453_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_453_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_453_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_653_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_653_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_653_completed_
      -- 
    cp_elements(148) <= cp_elements(163);
    -- CP-element group 149 transition  bypass 
    -- predecessors 161 
    -- successors 147 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_root_address_calculated
      -- 
    cp_elements(149) <= cp_elements(161);
    -- CP-element group 150 transition  bypass 
    -- predecessors 157 
    -- successors 158 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_indices_scaled
      -- 
    cp_elements(150) <= cp_elements(157);
    -- CP-element group 151 transition  bypass 
    -- predecessors 159 
    -- successors 160 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_offset_calculated
      -- 
    cp_elements(151) <= cp_elements(159);
    -- CP-element group 152 transition  bypass 
    -- predecessors 155 
    -- successors 156 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_resized_0
      -- 
    cp_elements(152) <= cp_elements(155);
    -- CP-element group 153 transition  bypass 
    -- predecessors 100 
    -- successors 154 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_450_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_450_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_450_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_computed_0
      -- 
    cp_elements(153) <= cp_elements(100);
    -- CP-element group 154 transition  output  bypass 
    -- predecessors 153 
    -- successors 155 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_resize_0/index_resize_req
      -- 
    cp_elements(154) <= cp_elements(153);
    index_resize_req_1633_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(154), ack => array_obj_ref_451_index_0_resize_req_0); -- 
    -- CP-element group 155 transition  input  bypass 
    -- predecessors 154 
    -- successors 152 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1634_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_index_0_resize_ack_0, ack => cp_elements(155)); -- 
    -- CP-element group 156 transition  output  bypass 
    -- predecessors 152 
    -- successors 157 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_scale_0/$entry
      -- 
    cp_elements(156) <= cp_elements(152);
    scale_rename_req_1638_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(156), ack => array_obj_ref_451_index_0_rename_req_0); -- 
    -- CP-element group 157 transition  input  bypass 
    -- predecessors 156 
    -- successors 150 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_index_scale_0/$exit
      -- 
    scale_rename_ack_1639_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_index_0_rename_ack_0, ack => cp_elements(157)); -- 
    -- CP-element group 158 transition  output  bypass 
    -- predecessors 150 
    -- successors 159 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_add_indices/final_index_req
      -- 
    cp_elements(158) <= cp_elements(150);
    final_index_req_1643_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(158), ack => array_obj_ref_451_offset_inst_req_0); -- 
    -- CP-element group 159 transition  input  bypass 
    -- predecessors 158 
    -- successors 151 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_add_indices/final_index_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_add_indices/$exit
      -- 
    final_index_ack_1644_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_offset_inst_ack_0, ack => cp_elements(159)); -- 
    -- CP-element group 160 transition  output  bypass 
    -- predecessors 151 
    -- successors 161 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_base_plus_offset/sum_rename_req
      -- 
    cp_elements(160) <= cp_elements(151);
    sum_rename_req_1648_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(160), ack => array_obj_ref_451_root_address_inst_req_0); -- 
    -- CP-element group 161 transition  input  bypass 
    -- predecessors 160 
    -- successors 149 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_451_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1649_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_451_root_address_inst_ack_0, ack => cp_elements(161)); -- 
    -- CP-element group 162 transition  output  bypass 
    -- predecessors 147 
    -- successors 163 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_complete/final_reg_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_complete/$entry
      -- 
    cp_elements(162) <= cp_elements(147);
    final_reg_req_1653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(162), ack => addr_of_452_final_reg_req_0); -- 
    -- CP-element group 163 transition  input  bypass 
    -- predecessors 162 
    -- successors 148 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_452_complete/final_reg_ack
      -- 
    final_reg_ack_1654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_452_final_reg_ack_0, ack => cp_elements(163)); -- 
    -- CP-element group 164 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_active_
      -- 
    cp_elements(164) <= cp_elements(7);
    -- CP-element group 165 join  fork  transition  bypass 
    -- predecessors 167 169 
    -- successors 182 200 218 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_459_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_459_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_459_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_completed_
      -- 
    cpelement_group_165 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(167);
      predecessors(1) <= cp_elements(169);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(165)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(165),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 166 join  transition  bypass 
    -- predecessors 170 
    -- marked predecessors 167 
    -- successors 171 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_sample_start_
      -- 
    cpelement_group_166 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(170);
      marked_predecessors(0) <= cp_elements(167);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(166)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 167 fork  transition  bypass 
    -- predecessors 172 
    -- successors 165 
    -- marked successors 166 27 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_sample_completed_
      -- 
    cp_elements(167) <= cp_elements(172);
    -- CP-element group 168 join  transition  bypass 
    -- predecessors 170 
    -- marked predecessors 177 195 213 
    -- successors 173 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_update_start_
      -- 
    cpelement_group_168 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(170);
      marked_predecessors(0) <= cp_elements(177);
      marked_predecessors(1) <= cp_elements(195);
      marked_predecessors(2) <= cp_elements(213);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(168)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 169 transition  bypass 
    -- predecessors 174 
    -- successors 165 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_update_completed_
      -- 
    cp_elements(169) <= cp_elements(174);
    -- CP-element group 170 fork  transition  bypass 
    -- predecessors 24 
    -- successors 166 168 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_455_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_455_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_455_trigger_
      -- 
    cp_elements(170) <= cp_elements(24);
    -- CP-element group 171 transition  output  bypass 
    -- predecessors 166 
    -- successors 172 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Sample/rr
      -- 
    cp_elements(171) <= cp_elements(166);
    rr_1671_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(171), ack => binary_458_inst_req_0); -- 
    -- CP-element group 172 transition  input  bypass 
    -- predecessors 171 
    -- successors 167 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Sample/ra
      -- 
    ra_1672_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_458_inst_ack_0, ack => cp_elements(172)); -- 
    -- CP-element group 173 transition  output  bypass 
    -- predecessors 168 
    -- successors 174 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Update/cr
      -- 
    cp_elements(173) <= cp_elements(168);
    cr_1676_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(173), ack => binary_458_inst_req_1); -- 
    -- CP-element group 174 transition  input  bypass 
    -- predecessors 173 
    -- successors 169 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_458_Update/ca
      -- 
    ca_1677_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_458_inst_ack_1, ack => cp_elements(174)); -- 
    -- CP-element group 175 transition  bypass 
    -- predecessors 7 
    -- successors 176 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_trigger_
      -- 
    cp_elements(175) <= cp_elements(7);
    -- CP-element group 176 join  transition  bypass 
    -- predecessors 175 178 
    -- marked predecessors 1047 
    -- successors 191 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_active_
      -- 
    cpelement_group_176 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(175);
      predecessors(1) <= cp_elements(178);
      marked_predecessors(0) <= cp_elements(1047);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(176)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(176),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 177 join  fork  transition  bypass 
    -- predecessors 192 
    -- marked predecessors 1050 
    -- successors 1048 
    -- marked successors 168 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_464_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_464_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_464_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_774_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_774_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_774_completed_
      -- 
    cpelement_group_177 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(192);
      marked_predecessors(0) <= cp_elements(1050);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(177)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(177),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 178 transition  bypass 
    -- predecessors 190 
    -- successors 176 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_root_address_calculated
      -- 
    cp_elements(178) <= cp_elements(190);
    -- CP-element group 179 transition  bypass 
    -- predecessors 186 
    -- successors 187 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_indices_scaled
      -- 
    cp_elements(179) <= cp_elements(186);
    -- CP-element group 180 transition  bypass 
    -- predecessors 188 
    -- successors 189 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_offset_calculated
      -- 
    cp_elements(180) <= cp_elements(188);
    -- CP-element group 181 transition  bypass 
    -- predecessors 184 
    -- successors 185 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_resized_0
      -- 
    cp_elements(181) <= cp_elements(184);
    -- CP-element group 182 transition  bypass 
    -- predecessors 165 
    -- successors 183 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_461_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_461_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_461_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_computed_0
      -- 
    cp_elements(182) <= cp_elements(165);
    -- CP-element group 183 transition  output  bypass 
    -- predecessors 182 
    -- successors 184 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_resize_0/index_resize_req
      -- 
    cp_elements(183) <= cp_elements(182);
    index_resize_req_1695_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(183), ack => array_obj_ref_462_index_0_resize_req_0); -- 
    -- CP-element group 184 transition  input  bypass 
    -- predecessors 183 
    -- successors 181 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_resize_0/$exit
      -- 
    index_resize_ack_1696_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_0_resize_ack_0, ack => cp_elements(184)); -- 
    -- CP-element group 185 transition  output  bypass 
    -- predecessors 181 
    -- successors 186 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_scale_0/$entry
      -- 
    cp_elements(185) <= cp_elements(181);
    scale_rename_req_1700_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(185), ack => array_obj_ref_462_index_0_rename_req_0); -- 
    -- CP-element group 186 transition  input  bypass 
    -- predecessors 185 
    -- successors 179 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1701_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_index_0_rename_ack_0, ack => cp_elements(186)); -- 
    -- CP-element group 187 transition  output  bypass 
    -- predecessors 179 
    -- successors 188 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_add_indices/final_index_req
      -- 
    cp_elements(187) <= cp_elements(179);
    final_index_req_1705_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(187), ack => array_obj_ref_462_offset_inst_req_0); -- 
    -- CP-element group 188 transition  input  bypass 
    -- predecessors 187 
    -- successors 180 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_add_indices/final_index_ack
      -- 
    final_index_ack_1706_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_offset_inst_ack_0, ack => cp_elements(188)); -- 
    -- CP-element group 189 transition  output  bypass 
    -- predecessors 180 
    -- successors 190 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_base_plus_offset/sum_rename_req
      -- 
    cp_elements(189) <= cp_elements(180);
    sum_rename_req_1710_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(189), ack => array_obj_ref_462_root_address_inst_req_0); -- 
    -- CP-element group 190 transition  input  bypass 
    -- predecessors 189 
    -- successors 178 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_462_base_plus_offset/$exit
      -- 
    sum_rename_ack_1711_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_462_root_address_inst_ack_0, ack => cp_elements(190)); -- 
    -- CP-element group 191 transition  output  bypass 
    -- predecessors 176 
    -- successors 192 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_complete/final_reg_req
      -- 
    cp_elements(191) <= cp_elements(176);
    final_reg_req_1715_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(191), ack => addr_of_463_final_reg_req_0); -- 
    -- CP-element group 192 transition  input  bypass 
    -- predecessors 191 
    -- successors 177 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_complete/final_reg_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_463_complete/$exit
      -- 
    final_reg_ack_1716_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_463_final_reg_ack_0, ack => cp_elements(192)); -- 
    -- CP-element group 193 transition  bypass 
    -- predecessors 7 
    -- successors 194 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_trigger_
      -- 
    cp_elements(193) <= cp_elements(7);
    -- CP-element group 194 join  transition  bypass 
    -- predecessors 193 196 
    -- marked predecessors 774 
    -- successors 209 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_active_
      -- 
    cpelement_group_194 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(193);
      predecessors(1) <= cp_elements(196);
      marked_predecessors(0) <= cp_elements(774);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(194)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(194),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 195 fork  transition  bypass 
    -- predecessors 210 
    -- successors 779 
    -- marked successors 168 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_469_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_469_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_469_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_644_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_644_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_644_completed_
      -- 
    cp_elements(195) <= cp_elements(210);
    -- CP-element group 196 transition  bypass 
    -- predecessors 208 
    -- successors 194 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_root_address_calculated
      -- 
    cp_elements(196) <= cp_elements(208);
    -- CP-element group 197 transition  bypass 
    -- predecessors 204 
    -- successors 205 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_indices_scaled
      -- 
    cp_elements(197) <= cp_elements(204);
    -- CP-element group 198 transition  bypass 
    -- predecessors 206 
    -- successors 207 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_offset_calculated
      -- 
    cp_elements(198) <= cp_elements(206);
    -- CP-element group 199 transition  bypass 
    -- predecessors 202 
    -- successors 203 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_resized_0
      -- 
    cp_elements(199) <= cp_elements(202);
    -- CP-element group 200 transition  bypass 
    -- predecessors 165 
    -- successors 201 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_466_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_466_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_466_trigger_
      -- 
    cp_elements(200) <= cp_elements(165);
    -- CP-element group 201 transition  output  bypass 
    -- predecessors 200 
    -- successors 202 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_resize_0/index_resize_req
      -- 
    cp_elements(201) <= cp_elements(200);
    index_resize_req_1734_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(201), ack => array_obj_ref_467_index_0_resize_req_0); -- 
    -- CP-element group 202 transition  input  bypass 
    -- predecessors 201 
    -- successors 199 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1735_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_467_index_0_resize_ack_0, ack => cp_elements(202)); -- 
    -- CP-element group 203 transition  output  bypass 
    -- predecessors 199 
    -- successors 204 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_scale_0/scale_rename_req
      -- 
    cp_elements(203) <= cp_elements(199);
    scale_rename_req_1739_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(203), ack => array_obj_ref_467_index_0_rename_req_0); -- 
    -- CP-element group 204 transition  input  bypass 
    -- predecessors 203 
    -- successors 197 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1740_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_467_index_0_rename_ack_0, ack => cp_elements(204)); -- 
    -- CP-element group 205 transition  output  bypass 
    -- predecessors 197 
    -- successors 206 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_add_indices/final_index_req
      -- 
    cp_elements(205) <= cp_elements(197);
    final_index_req_1744_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(205), ack => array_obj_ref_467_offset_inst_req_0); -- 
    -- CP-element group 206 transition  input  bypass 
    -- predecessors 205 
    -- successors 198 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_add_indices/final_index_ack
      -- 
    final_index_ack_1745_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_467_offset_inst_ack_0, ack => cp_elements(206)); -- 
    -- CP-element group 207 transition  output  bypass 
    -- predecessors 198 
    -- successors 208 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_base_plus_offset/sum_rename_req
      -- 
    cp_elements(207) <= cp_elements(198);
    sum_rename_req_1749_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(207), ack => array_obj_ref_467_root_address_inst_req_0); -- 
    -- CP-element group 208 transition  input  bypass 
    -- predecessors 207 
    -- successors 196 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_467_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1750_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_467_root_address_inst_ack_0, ack => cp_elements(208)); -- 
    -- CP-element group 209 transition  output  bypass 
    -- predecessors 194 
    -- successors 210 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_complete/final_reg_req
      -- 
    cp_elements(209) <= cp_elements(194);
    final_reg_req_1754_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(209), ack => addr_of_468_final_reg_req_0); -- 
    -- CP-element group 210 transition  input  bypass 
    -- predecessors 209 
    -- successors 195 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_468_complete/final_reg_ack
      -- 
    final_reg_ack_1755_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_468_final_reg_ack_0, ack => cp_elements(210)); -- 
    -- CP-element group 211 transition  bypass 
    -- predecessors 7 
    -- successors 212 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_trigger_
      -- 
    cp_elements(211) <= cp_elements(7);
    -- CP-element group 212 join  transition  bypass 
    -- predecessors 211 214 
    -- marked predecessors 758 
    -- successors 227 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_active_
      -- 
    cpelement_group_212 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(211);
      predecessors(1) <= cp_elements(214);
      marked_predecessors(0) <= cp_elements(758);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(212)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(212),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 213 fork  transition  bypass 
    -- predecessors 228 
    -- successors 763 
    -- marked successors 168 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_474_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_474_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_474_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_640_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_640_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_640_completed_
      -- 
    cp_elements(213) <= cp_elements(228);
    -- CP-element group 214 transition  bypass 
    -- predecessors 226 
    -- successors 212 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_root_address_calculated
      -- 
    cp_elements(214) <= cp_elements(226);
    -- CP-element group 215 transition  bypass 
    -- predecessors 222 
    -- successors 223 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_indices_scaled
      -- 
    cp_elements(215) <= cp_elements(222);
    -- CP-element group 216 transition  bypass 
    -- predecessors 224 
    -- successors 225 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_offset_calculated
      -- 
    cp_elements(216) <= cp_elements(224);
    -- CP-element group 217 transition  bypass 
    -- predecessors 220 
    -- successors 221 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_resized_0
      -- 
    cp_elements(217) <= cp_elements(220);
    -- CP-element group 218 transition  bypass 
    -- predecessors 165 
    -- successors 219 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_471_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_471_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_471_completed_
      -- 
    cp_elements(218) <= cp_elements(165);
    -- CP-element group 219 transition  output  bypass 
    -- predecessors 218 
    -- successors 220 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_resize_0/index_resize_req
      -- 
    cp_elements(219) <= cp_elements(218);
    index_resize_req_1773_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(219), ack => array_obj_ref_472_index_0_resize_req_0); -- 
    -- CP-element group 220 transition  input  bypass 
    -- predecessors 219 
    -- successors 217 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1774_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_472_index_0_resize_ack_0, ack => cp_elements(220)); -- 
    -- CP-element group 221 transition  output  bypass 
    -- predecessors 217 
    -- successors 222 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_scale_0/scale_rename_req
      -- 
    cp_elements(221) <= cp_elements(217);
    scale_rename_req_1778_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(221), ack => array_obj_ref_472_index_0_rename_req_0); -- 
    -- CP-element group 222 transition  input  bypass 
    -- predecessors 221 
    -- successors 215 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1779_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_472_index_0_rename_ack_0, ack => cp_elements(222)); -- 
    -- CP-element group 223 transition  output  bypass 
    -- predecessors 215 
    -- successors 224 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_add_indices/final_index_req
      -- 
    cp_elements(223) <= cp_elements(215);
    final_index_req_1783_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(223), ack => array_obj_ref_472_offset_inst_req_0); -- 
    -- CP-element group 224 transition  input  bypass 
    -- predecessors 223 
    -- successors 216 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_add_indices/final_index_ack
      -- 
    final_index_ack_1784_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_472_offset_inst_ack_0, ack => cp_elements(224)); -- 
    -- CP-element group 225 transition  output  bypass 
    -- predecessors 216 
    -- successors 226 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_base_plus_offset/sum_rename_req
      -- 
    cp_elements(225) <= cp_elements(216);
    sum_rename_req_1788_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(225), ack => array_obj_ref_472_root_address_inst_req_0); -- 
    -- CP-element group 226 transition  input  bypass 
    -- predecessors 225 
    -- successors 214 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_472_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1789_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_472_root_address_inst_ack_0, ack => cp_elements(226)); -- 
    -- CP-element group 227 transition  output  bypass 
    -- predecessors 212 
    -- successors 228 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_complete/final_reg_req
      -- 
    cp_elements(227) <= cp_elements(212);
    final_reg_req_1793_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(227), ack => addr_of_473_final_reg_req_0); -- 
    -- CP-element group 228 transition  input  bypass 
    -- predecessors 227 
    -- successors 213 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_473_complete/final_reg_ack
      -- 
    final_reg_ack_1794_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_473_final_reg_ack_0, ack => cp_elements(228)); -- 
    -- CP-element group 229 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_active_
      -- 
    cp_elements(229) <= cp_elements(7);
    -- CP-element group 230 join  fork  transition  bypass 
    -- predecessors 232 234 
    -- successors 247 265 283 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_480_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_480_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_480_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_completed_
      -- 
    cpelement_group_230 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(232);
      predecessors(1) <= cp_elements(234);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(230)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(230),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 231 join  transition  bypass 
    -- predecessors 235 
    -- marked predecessors 232 
    -- successors 236 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_sample_start_
      -- 
    cpelement_group_231 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(235);
      marked_predecessors(0) <= cp_elements(232);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(231)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(231),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 232 fork  transition  bypass 
    -- predecessors 237 
    -- successors 230 
    -- marked successors 27 231 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_sample_completed_
      -- 
    cp_elements(232) <= cp_elements(237);
    -- CP-element group 233 join  transition  bypass 
    -- predecessors 235 
    -- marked predecessors 242 260 278 
    -- successors 238 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_update_start_
      -- 
    cpelement_group_233 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(235);
      marked_predecessors(0) <= cp_elements(242);
      marked_predecessors(1) <= cp_elements(260);
      marked_predecessors(2) <= cp_elements(278);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(233)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(233),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 234 transition  bypass 
    -- predecessors 239 
    -- successors 230 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_update_completed_
      -- 
    cp_elements(234) <= cp_elements(239);
    -- CP-element group 235 fork  transition  bypass 
    -- predecessors 24 
    -- successors 231 233 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_476_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_476_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_476_completed_
      -- 
    cp_elements(235) <= cp_elements(24);
    -- CP-element group 236 transition  output  bypass 
    -- predecessors 231 
    -- successors 237 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Sample/rr
      -- 
    cp_elements(236) <= cp_elements(231);
    rr_1811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(236), ack => binary_479_inst_req_0); -- 
    -- CP-element group 237 transition  input  bypass 
    -- predecessors 236 
    -- successors 232 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Sample/ra
      -- 
    ra_1812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_479_inst_ack_0, ack => cp_elements(237)); -- 
    -- CP-element group 238 transition  output  bypass 
    -- predecessors 233 
    -- successors 239 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Update/cr
      -- 
    cp_elements(238) <= cp_elements(233);
    cr_1816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(238), ack => binary_479_inst_req_1); -- 
    -- CP-element group 239 transition  input  bypass 
    -- predecessors 238 
    -- successors 234 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_479_Update/ca
      -- 
    ca_1817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_479_inst_ack_1, ack => cp_elements(239)); -- 
    -- CP-element group 240 transition  bypass 
    -- predecessors 7 
    -- successors 241 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_trigger_
      -- 
    cp_elements(240) <= cp_elements(7);
    -- CP-element group 241 join  transition  bypass 
    -- predecessors 240 243 
    -- marked predecessors 1015 
    -- successors 256 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_active_
      -- 
    cpelement_group_241 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(240);
      predecessors(1) <= cp_elements(243);
      marked_predecessors(0) <= cp_elements(1015);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(241)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(241),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 242 join  fork  transition  bypass 
    -- predecessors 257 
    -- marked predecessors 1018 
    -- successors 1016 
    -- marked successors 233 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_485_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_485_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_485_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_755_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_755_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_755_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_trigger_
      -- 
    cpelement_group_242 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(257);
      marked_predecessors(0) <= cp_elements(1018);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(242)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(242),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 243 transition  bypass 
    -- predecessors 255 
    -- successors 241 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_root_address_calculated
      -- 
    cp_elements(243) <= cp_elements(255);
    -- CP-element group 244 transition  bypass 
    -- predecessors 251 
    -- successors 252 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_indices_scaled
      -- 
    cp_elements(244) <= cp_elements(251);
    -- CP-element group 245 transition  bypass 
    -- predecessors 253 
    -- successors 254 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_offset_calculated
      -- 
    cp_elements(245) <= cp_elements(253);
    -- CP-element group 246 transition  bypass 
    -- predecessors 249 
    -- successors 250 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_resized_0
      -- 
    cp_elements(246) <= cp_elements(249);
    -- CP-element group 247 transition  bypass 
    -- predecessors 230 
    -- successors 248 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_482_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_482_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_482_completed_
      -- 
    cp_elements(247) <= cp_elements(230);
    -- CP-element group 248 transition  output  bypass 
    -- predecessors 247 
    -- successors 249 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_resize_0/index_resize_req
      -- 
    cp_elements(248) <= cp_elements(247);
    index_resize_req_1835_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(248), ack => array_obj_ref_483_index_0_resize_req_0); -- 
    -- CP-element group 249 transition  input  bypass 
    -- predecessors 248 
    -- successors 246 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1836_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_index_0_resize_ack_0, ack => cp_elements(249)); -- 
    -- CP-element group 250 transition  output  bypass 
    -- predecessors 246 
    -- successors 251 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_scale_0/scale_rename_req
      -- 
    cp_elements(250) <= cp_elements(246);
    scale_rename_req_1840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(250), ack => array_obj_ref_483_index_0_rename_req_0); -- 
    -- CP-element group 251 transition  input  bypass 
    -- predecessors 250 
    -- successors 244 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_index_0_rename_ack_0, ack => cp_elements(251)); -- 
    -- CP-element group 252 transition  output  bypass 
    -- predecessors 244 
    -- successors 253 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_add_indices/final_index_req
      -- 
    cp_elements(252) <= cp_elements(244);
    final_index_req_1845_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(252), ack => array_obj_ref_483_offset_inst_req_0); -- 
    -- CP-element group 253 transition  input  bypass 
    -- predecessors 252 
    -- successors 245 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_add_indices/final_index_ack
      -- 
    final_index_ack_1846_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_offset_inst_ack_0, ack => cp_elements(253)); -- 
    -- CP-element group 254 transition  output  bypass 
    -- predecessors 245 
    -- successors 255 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_base_plus_offset/sum_rename_req
      -- 
    cp_elements(254) <= cp_elements(245);
    sum_rename_req_1850_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(254), ack => array_obj_ref_483_root_address_inst_req_0); -- 
    -- CP-element group 255 transition  input  bypass 
    -- predecessors 254 
    -- successors 243 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_483_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1851_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_483_root_address_inst_ack_0, ack => cp_elements(255)); -- 
    -- CP-element group 256 transition  output  bypass 
    -- predecessors 241 
    -- successors 257 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_complete/final_reg_req
      -- 
    cp_elements(256) <= cp_elements(241);
    final_reg_req_1855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(256), ack => addr_of_484_final_reg_req_0); -- 
    -- CP-element group 257 transition  input  bypass 
    -- predecessors 256 
    -- successors 242 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_484_complete/final_reg_ack
      -- 
    final_reg_ack_1856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_484_final_reg_ack_0, ack => cp_elements(257)); -- 
    -- CP-element group 258 transition  bypass 
    -- predecessors 7 
    -- successors 259 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_trigger_
      -- 
    cp_elements(258) <= cp_elements(7);
    -- CP-element group 259 join  transition  bypass 
    -- predecessors 258 261 
    -- marked predecessors 731 
    -- successors 274 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_active_
      -- 
    cpelement_group_259 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(258);
      predecessors(1) <= cp_elements(261);
      marked_predecessors(0) <= cp_elements(731);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(259)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(259),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 260 fork  transition  bypass 
    -- predecessors 275 
    -- successors 736 
    -- marked successors 233 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_490_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_490_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_490_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_631_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_631_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_631_completed_
      -- 
    cp_elements(260) <= cp_elements(275);
    -- CP-element group 261 transition  bypass 
    -- predecessors 273 
    -- successors 259 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_root_address_calculated
      -- 
    cp_elements(261) <= cp_elements(273);
    -- CP-element group 262 transition  bypass 
    -- predecessors 269 
    -- successors 270 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_indices_scaled
      -- 
    cp_elements(262) <= cp_elements(269);
    -- CP-element group 263 transition  bypass 
    -- predecessors 271 
    -- successors 272 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_offset_calculated
      -- 
    cp_elements(263) <= cp_elements(271);
    -- CP-element group 264 transition  bypass 
    -- predecessors 267 
    -- successors 268 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_resized_0
      -- 
    cp_elements(264) <= cp_elements(267);
    -- CP-element group 265 transition  bypass 
    -- predecessors 230 
    -- successors 266 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_487_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_487_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_487_completed_
      -- 
    cp_elements(265) <= cp_elements(230);
    -- CP-element group 266 transition  output  bypass 
    -- predecessors 265 
    -- successors 267 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_resize_0/index_resize_req
      -- 
    cp_elements(266) <= cp_elements(265);
    index_resize_req_1874_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(266), ack => array_obj_ref_488_index_0_resize_req_0); -- 
    -- CP-element group 267 transition  input  bypass 
    -- predecessors 266 
    -- successors 264 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1875_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_488_index_0_resize_ack_0, ack => cp_elements(267)); -- 
    -- CP-element group 268 transition  output  bypass 
    -- predecessors 264 
    -- successors 269 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_scale_0/scale_rename_req
      -- 
    cp_elements(268) <= cp_elements(264);
    scale_rename_req_1879_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(268), ack => array_obj_ref_488_index_0_rename_req_0); -- 
    -- CP-element group 269 transition  input  bypass 
    -- predecessors 268 
    -- successors 262 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1880_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_488_index_0_rename_ack_0, ack => cp_elements(269)); -- 
    -- CP-element group 270 transition  output  bypass 
    -- predecessors 262 
    -- successors 271 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_add_indices/final_index_req
      -- 
    cp_elements(270) <= cp_elements(262);
    final_index_req_1884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(270), ack => array_obj_ref_488_offset_inst_req_0); -- 
    -- CP-element group 271 transition  input  bypass 
    -- predecessors 270 
    -- successors 263 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_add_indices/final_index_ack
      -- 
    final_index_ack_1885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_488_offset_inst_ack_0, ack => cp_elements(271)); -- 
    -- CP-element group 272 transition  output  bypass 
    -- predecessors 263 
    -- successors 273 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_base_plus_offset/sum_rename_req
      -- 
    cp_elements(272) <= cp_elements(263);
    sum_rename_req_1889_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(272), ack => array_obj_ref_488_root_address_inst_req_0); -- 
    -- CP-element group 273 transition  input  bypass 
    -- predecessors 272 
    -- successors 261 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_488_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1890_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_488_root_address_inst_ack_0, ack => cp_elements(273)); -- 
    -- CP-element group 274 transition  output  bypass 
    -- predecessors 259 
    -- successors 275 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_complete/final_reg_req
      -- 
    cp_elements(274) <= cp_elements(259);
    final_reg_req_1894_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(274), ack => addr_of_489_final_reg_req_0); -- 
    -- CP-element group 275 transition  input  bypass 
    -- predecessors 274 
    -- successors 260 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_489_complete/final_reg_ack
      -- 
    final_reg_ack_1895_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_489_final_reg_ack_0, ack => cp_elements(275)); -- 
    -- CP-element group 276 transition  bypass 
    -- predecessors 7 
    -- successors 277 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_trigger_
      -- 
    cp_elements(276) <= cp_elements(7);
    -- CP-element group 277 join  transition  bypass 
    -- predecessors 276 279 
    -- marked predecessors 715 
    -- successors 292 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_active_
      -- 
    cpelement_group_277 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(276);
      predecessors(1) <= cp_elements(279);
      marked_predecessors(0) <= cp_elements(715);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(277)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(277),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 278 fork  transition  bypass 
    -- predecessors 293 
    -- successors 720 
    -- marked successors 233 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_495_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_495_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_495_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_627_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_627_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_627_completed_
      -- 
    cp_elements(278) <= cp_elements(293);
    -- CP-element group 279 transition  bypass 
    -- predecessors 291 
    -- successors 277 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_root_address_calculated
      -- 
    cp_elements(279) <= cp_elements(291);
    -- CP-element group 280 transition  bypass 
    -- predecessors 287 
    -- successors 288 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_indices_scaled
      -- 
    cp_elements(280) <= cp_elements(287);
    -- CP-element group 281 transition  bypass 
    -- predecessors 289 
    -- successors 290 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_offset_calculated
      -- 
    cp_elements(281) <= cp_elements(289);
    -- CP-element group 282 transition  bypass 
    -- predecessors 285 
    -- successors 286 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_resized_0
      -- 
    cp_elements(282) <= cp_elements(285);
    -- CP-element group 283 transition  bypass 
    -- predecessors 230 
    -- successors 284 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_492_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_492_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_492_completed_
      -- 
    cp_elements(283) <= cp_elements(230);
    -- CP-element group 284 transition  output  bypass 
    -- predecessors 283 
    -- successors 285 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_resize_0/index_resize_req
      -- 
    cp_elements(284) <= cp_elements(283);
    index_resize_req_1913_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(284), ack => array_obj_ref_493_index_0_resize_req_0); -- 
    -- CP-element group 285 transition  input  bypass 
    -- predecessors 284 
    -- successors 282 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1914_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_493_index_0_resize_ack_0, ack => cp_elements(285)); -- 
    -- CP-element group 286 transition  output  bypass 
    -- predecessors 282 
    -- successors 287 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_scale_0/scale_rename_req
      -- 
    cp_elements(286) <= cp_elements(282);
    scale_rename_req_1918_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(286), ack => array_obj_ref_493_index_0_rename_req_0); -- 
    -- CP-element group 287 transition  input  bypass 
    -- predecessors 286 
    -- successors 280 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1919_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_493_index_0_rename_ack_0, ack => cp_elements(287)); -- 
    -- CP-element group 288 transition  output  bypass 
    -- predecessors 280 
    -- successors 289 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_add_indices/final_index_req
      -- 
    cp_elements(288) <= cp_elements(280);
    final_index_req_1923_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(288), ack => array_obj_ref_493_offset_inst_req_0); -- 
    -- CP-element group 289 transition  input  bypass 
    -- predecessors 288 
    -- successors 281 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_add_indices/final_index_ack
      -- 
    final_index_ack_1924_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_493_offset_inst_ack_0, ack => cp_elements(289)); -- 
    -- CP-element group 290 transition  output  bypass 
    -- predecessors 281 
    -- successors 291 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_base_plus_offset/sum_rename_req
      -- 
    cp_elements(290) <= cp_elements(281);
    sum_rename_req_1928_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(290), ack => array_obj_ref_493_root_address_inst_req_0); -- 
    -- CP-element group 291 transition  input  bypass 
    -- predecessors 290 
    -- successors 279 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_493_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1929_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_493_root_address_inst_ack_0, ack => cp_elements(291)); -- 
    -- CP-element group 292 transition  output  bypass 
    -- predecessors 277 
    -- successors 293 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_complete/final_reg_req
      -- 
    cp_elements(292) <= cp_elements(277);
    final_reg_req_1933_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(292), ack => addr_of_494_final_reg_req_0); -- 
    -- CP-element group 293 transition  input  bypass 
    -- predecessors 292 
    -- successors 278 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_494_complete/final_reg_ack
      -- 
    final_reg_ack_1934_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_494_final_reg_ack_0, ack => cp_elements(293)); -- 
    -- CP-element group 294 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_active_
      -- 
    cp_elements(294) <= cp_elements(7);
    -- CP-element group 295 join  fork  transition  bypass 
    -- predecessors 297 299 
    -- successors 348 312 330 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_501_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_501_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_501_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_completed_
      -- 
    cpelement_group_295 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(297);
      predecessors(1) <= cp_elements(299);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(295)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(295),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 296 join  transition  bypass 
    -- predecessors 300 
    -- marked predecessors 297 
    -- successors 301 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_sample_start_
      -- 
    cpelement_group_296 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(300);
      marked_predecessors(0) <= cp_elements(297);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(296)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(296),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 297 fork  transition  bypass 
    -- predecessors 302 
    -- successors 295 
    -- marked successors 27 296 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_sample_completed_
      -- 
    cp_elements(297) <= cp_elements(302);
    -- CP-element group 298 join  transition  bypass 
    -- predecessors 300 
    -- marked predecessors 343 307 325 
    -- successors 303 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_update_start_
      -- 
    cpelement_group_298 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(300);
      marked_predecessors(0) <= cp_elements(343);
      marked_predecessors(1) <= cp_elements(307);
      marked_predecessors(2) <= cp_elements(325);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(298)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(298),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 299 transition  bypass 
    -- predecessors 304 
    -- successors 295 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_update_completed_
      -- 
    cp_elements(299) <= cp_elements(304);
    -- CP-element group 300 fork  transition  bypass 
    -- predecessors 24 
    -- successors 296 298 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_497_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_497_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_497_completed_
      -- 
    cp_elements(300) <= cp_elements(24);
    -- CP-element group 301 transition  output  bypass 
    -- predecessors 296 
    -- successors 302 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Sample/rr
      -- 
    cp_elements(301) <= cp_elements(296);
    rr_1951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(301), ack => binary_500_inst_req_0); -- 
    -- CP-element group 302 transition  input  bypass 
    -- predecessors 301 
    -- successors 297 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Sample/ra
      -- 
    ra_1952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_500_inst_ack_0, ack => cp_elements(302)); -- 
    -- CP-element group 303 transition  output  bypass 
    -- predecessors 298 
    -- successors 304 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Update/cr
      -- 
    cp_elements(303) <= cp_elements(298);
    cr_1956_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(303), ack => binary_500_inst_req_1); -- 
    -- CP-element group 304 transition  input  bypass 
    -- predecessors 303 
    -- successors 299 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_500_Update/ca
      -- 
    ca_1957_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_500_inst_ack_1, ack => cp_elements(304)); -- 
    -- CP-element group 305 transition  bypass 
    -- predecessors 7 
    -- successors 306 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_trigger_
      -- 
    cp_elements(305) <= cp_elements(7);
    -- CP-element group 306 join  transition  bypass 
    -- predecessors 308 305 
    -- marked predecessors 983 
    -- successors 321 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_active_
      -- 
    cpelement_group_306 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(308);
      predecessors(1) <= cp_elements(305);
      marked_predecessors(0) <= cp_elements(983);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(306)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(306),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 307 join  fork  transition  bypass 
    -- predecessors 322 
    -- marked predecessors 986 
    -- successors 984 
    -- marked successors 298 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_506_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_506_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_506_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_736_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_736_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_736_active_
      -- 
    cpelement_group_307 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(322);
      marked_predecessors(0) <= cp_elements(986);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(307)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(307),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 308 transition  bypass 
    -- predecessors 320 
    -- successors 306 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_root_address_calculated
      -- 
    cp_elements(308) <= cp_elements(320);
    -- CP-element group 309 transition  bypass 
    -- predecessors 316 
    -- successors 317 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_indices_scaled
      -- 
    cp_elements(309) <= cp_elements(316);
    -- CP-element group 310 transition  bypass 
    -- predecessors 318 
    -- successors 319 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_offset_calculated
      -- 
    cp_elements(310) <= cp_elements(318);
    -- CP-element group 311 transition  bypass 
    -- predecessors 314 
    -- successors 315 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_resized_0
      -- 
    cp_elements(311) <= cp_elements(314);
    -- CP-element group 312 transition  bypass 
    -- predecessors 295 
    -- successors 313 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_503_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_503_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_503_completed_
      -- 
    cp_elements(312) <= cp_elements(295);
    -- CP-element group 313 transition  output  bypass 
    -- predecessors 312 
    -- successors 314 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_resize_0/index_resize_req
      -- 
    cp_elements(313) <= cp_elements(312);
    index_resize_req_1975_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(313), ack => array_obj_ref_504_index_0_resize_req_0); -- 
    -- CP-element group 314 transition  input  bypass 
    -- predecessors 313 
    -- successors 311 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_1976_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_504_index_0_resize_ack_0, ack => cp_elements(314)); -- 
    -- CP-element group 315 transition  output  bypass 
    -- predecessors 311 
    -- successors 316 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_scale_0/scale_rename_req
      -- 
    cp_elements(315) <= cp_elements(311);
    scale_rename_req_1980_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(315), ack => array_obj_ref_504_index_0_rename_req_0); -- 
    -- CP-element group 316 transition  input  bypass 
    -- predecessors 315 
    -- successors 309 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_1981_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_504_index_0_rename_ack_0, ack => cp_elements(316)); -- 
    -- CP-element group 317 transition  output  bypass 
    -- predecessors 309 
    -- successors 318 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_add_indices/final_index_req
      -- 
    cp_elements(317) <= cp_elements(309);
    final_index_req_1985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(317), ack => array_obj_ref_504_offset_inst_req_0); -- 
    -- CP-element group 318 transition  input  bypass 
    -- predecessors 317 
    -- successors 310 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_add_indices/final_index_ack
      -- 
    final_index_ack_1986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_504_offset_inst_ack_0, ack => cp_elements(318)); -- 
    -- CP-element group 319 transition  output  bypass 
    -- predecessors 310 
    -- successors 320 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_base_plus_offset/sum_rename_req
      -- 
    cp_elements(319) <= cp_elements(310);
    sum_rename_req_1990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(319), ack => array_obj_ref_504_root_address_inst_req_0); -- 
    -- CP-element group 320 transition  input  bypass 
    -- predecessors 319 
    -- successors 308 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_504_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_1991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_504_root_address_inst_ack_0, ack => cp_elements(320)); -- 
    -- CP-element group 321 transition  output  bypass 
    -- predecessors 306 
    -- successors 322 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_complete/final_reg_req
      -- 
    cp_elements(321) <= cp_elements(306);
    final_reg_req_1995_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(321), ack => addr_of_505_final_reg_req_0); -- 
    -- CP-element group 322 transition  input  bypass 
    -- predecessors 321 
    -- successors 307 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_505_complete/final_reg_ack
      -- 
    final_reg_ack_1996_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_505_final_reg_ack_0, ack => cp_elements(322)); -- 
    -- CP-element group 323 transition  bypass 
    -- predecessors 7 
    -- successors 324 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_trigger_
      -- 
    cp_elements(323) <= cp_elements(7);
    -- CP-element group 324 join  transition  bypass 
    -- predecessors 323 326 
    -- marked predecessors 688 
    -- successors 339 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_active_
      -- 
    cpelement_group_324 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(323);
      predecessors(1) <= cp_elements(326);
      marked_predecessors(0) <= cp_elements(688);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(324)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(324),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 325 fork  transition  bypass 
    -- predecessors 340 
    -- successors 693 
    -- marked successors 298 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_511_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_511_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_511_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_618_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_618_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_618_completed_
      -- 
    cp_elements(325) <= cp_elements(340);
    -- CP-element group 326 transition  bypass 
    -- predecessors 338 
    -- successors 324 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_root_address_calculated
      -- 
    cp_elements(326) <= cp_elements(338);
    -- CP-element group 327 transition  bypass 
    -- predecessors 334 
    -- successors 335 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_indices_scaled
      -- 
    cp_elements(327) <= cp_elements(334);
    -- CP-element group 328 transition  bypass 
    -- predecessors 336 
    -- successors 337 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_offset_calculated
      -- 
    cp_elements(328) <= cp_elements(336);
    -- CP-element group 329 transition  bypass 
    -- predecessors 332 
    -- successors 333 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_resized_0
      -- 
    cp_elements(329) <= cp_elements(332);
    -- CP-element group 330 transition  bypass 
    -- predecessors 295 
    -- successors 331 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_508_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_508_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_508_completed_
      -- 
    cp_elements(330) <= cp_elements(295);
    -- CP-element group 331 transition  output  bypass 
    -- predecessors 330 
    -- successors 332 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_resize_0/index_resize_req
      -- 
    cp_elements(331) <= cp_elements(330);
    index_resize_req_2014_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(331), ack => array_obj_ref_509_index_0_resize_req_0); -- 
    -- CP-element group 332 transition  input  bypass 
    -- predecessors 331 
    -- successors 329 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2015_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_509_index_0_resize_ack_0, ack => cp_elements(332)); -- 
    -- CP-element group 333 transition  output  bypass 
    -- predecessors 329 
    -- successors 334 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_scale_0/scale_rename_req
      -- 
    cp_elements(333) <= cp_elements(329);
    scale_rename_req_2019_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(333), ack => array_obj_ref_509_index_0_rename_req_0); -- 
    -- CP-element group 334 transition  input  bypass 
    -- predecessors 333 
    -- successors 327 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2020_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_509_index_0_rename_ack_0, ack => cp_elements(334)); -- 
    -- CP-element group 335 transition  output  bypass 
    -- predecessors 327 
    -- successors 336 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_add_indices/final_index_req
      -- 
    cp_elements(335) <= cp_elements(327);
    final_index_req_2024_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(335), ack => array_obj_ref_509_offset_inst_req_0); -- 
    -- CP-element group 336 transition  input  bypass 
    -- predecessors 335 
    -- successors 328 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_add_indices/final_index_ack
      -- 
    final_index_ack_2025_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_509_offset_inst_ack_0, ack => cp_elements(336)); -- 
    -- CP-element group 337 transition  output  bypass 
    -- predecessors 328 
    -- successors 338 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_base_plus_offset/sum_rename_req
      -- 
    cp_elements(337) <= cp_elements(328);
    sum_rename_req_2029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(337), ack => array_obj_ref_509_root_address_inst_req_0); -- 
    -- CP-element group 338 transition  input  bypass 
    -- predecessors 337 
    -- successors 326 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_509_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_509_root_address_inst_ack_0, ack => cp_elements(338)); -- 
    -- CP-element group 339 transition  output  bypass 
    -- predecessors 324 
    -- successors 340 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_complete/final_reg_req
      -- 
    cp_elements(339) <= cp_elements(324);
    final_reg_req_2034_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(339), ack => addr_of_510_final_reg_req_0); -- 
    -- CP-element group 340 transition  input  bypass 
    -- predecessors 339 
    -- successors 325 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_510_complete/final_reg_ack
      -- 
    final_reg_ack_2035_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_510_final_reg_ack_0, ack => cp_elements(340)); -- 
    -- CP-element group 341 transition  bypass 
    -- predecessors 7 
    -- successors 342 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_trigger_
      -- 
    cp_elements(341) <= cp_elements(7);
    -- CP-element group 342 join  transition  bypass 
    -- predecessors 341 344 
    -- marked predecessors 672 
    -- successors 357 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_active_
      -- 
    cpelement_group_342 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(341);
      predecessors(1) <= cp_elements(344);
      marked_predecessors(0) <= cp_elements(672);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(342)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(342),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 343 fork  transition  bypass 
    -- predecessors 358 
    -- successors 677 
    -- marked successors 298 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_516_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_516_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_516_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_614_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_614_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_614_completed_
      -- 
    cp_elements(343) <= cp_elements(358);
    -- CP-element group 344 transition  bypass 
    -- predecessors 356 
    -- successors 342 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_root_address_calculated
      -- 
    cp_elements(344) <= cp_elements(356);
    -- CP-element group 345 transition  bypass 
    -- predecessors 352 
    -- successors 353 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_indices_scaled
      -- 
    cp_elements(345) <= cp_elements(352);
    -- CP-element group 346 transition  bypass 
    -- predecessors 354 
    -- successors 355 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_offset_calculated
      -- 
    cp_elements(346) <= cp_elements(354);
    -- CP-element group 347 transition  bypass 
    -- predecessors 350 
    -- successors 351 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_resized_0
      -- 
    cp_elements(347) <= cp_elements(350);
    -- CP-element group 348 transition  bypass 
    -- predecessors 295 
    -- successors 349 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_513_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_513_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_513_completed_
      -- 
    cp_elements(348) <= cp_elements(295);
    -- CP-element group 349 transition  output  bypass 
    -- predecessors 348 
    -- successors 350 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_resize_0/index_resize_req
      -- 
    cp_elements(349) <= cp_elements(348);
    index_resize_req_2053_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(349), ack => array_obj_ref_514_index_0_resize_req_0); -- 
    -- CP-element group 350 transition  input  bypass 
    -- predecessors 349 
    -- successors 347 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2054_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_index_0_resize_ack_0, ack => cp_elements(350)); -- 
    -- CP-element group 351 transition  output  bypass 
    -- predecessors 347 
    -- successors 352 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_scale_0/scale_rename_req
      -- 
    cp_elements(351) <= cp_elements(347);
    scale_rename_req_2058_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(351), ack => array_obj_ref_514_index_0_rename_req_0); -- 
    -- CP-element group 352 transition  input  bypass 
    -- predecessors 351 
    -- successors 345 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2059_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_index_0_rename_ack_0, ack => cp_elements(352)); -- 
    -- CP-element group 353 transition  output  bypass 
    -- predecessors 345 
    -- successors 354 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_add_indices/final_index_req
      -- 
    cp_elements(353) <= cp_elements(345);
    final_index_req_2063_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(353), ack => array_obj_ref_514_offset_inst_req_0); -- 
    -- CP-element group 354 transition  input  bypass 
    -- predecessors 353 
    -- successors 346 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_add_indices/final_index_ack
      -- 
    final_index_ack_2064_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_offset_inst_ack_0, ack => cp_elements(354)); -- 
    -- CP-element group 355 transition  output  bypass 
    -- predecessors 346 
    -- successors 356 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_base_plus_offset/sum_rename_req
      -- 
    cp_elements(355) <= cp_elements(346);
    sum_rename_req_2068_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(355), ack => array_obj_ref_514_root_address_inst_req_0); -- 
    -- CP-element group 356 transition  input  bypass 
    -- predecessors 355 
    -- successors 344 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_514_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2069_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_514_root_address_inst_ack_0, ack => cp_elements(356)); -- 
    -- CP-element group 357 transition  output  bypass 
    -- predecessors 342 
    -- successors 358 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_complete/final_reg_req
      -- 
    cp_elements(357) <= cp_elements(342);
    final_reg_req_2073_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(357), ack => addr_of_515_final_reg_req_0); -- 
    -- CP-element group 358 transition  input  bypass 
    -- predecessors 357 
    -- successors 343 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_515_complete/final_reg_ack
      -- 
    final_reg_ack_2074_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_515_final_reg_ack_0, ack => cp_elements(358)); -- 
    -- CP-element group 359 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_active_
      -- 
    cp_elements(359) <= cp_elements(7);
    -- CP-element group 360 join  fork  transition  bypass 
    -- predecessors 362 364 
    -- successors 377 395 413 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_522_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_522_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_522_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_completed_
      -- 
    cpelement_group_360 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(362);
      predecessors(1) <= cp_elements(364);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(360)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(360),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 361 join  transition  bypass 
    -- predecessors 365 
    -- marked predecessors 362 
    -- successors 366 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_sample_start_
      -- 
    cpelement_group_361 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(365);
      marked_predecessors(0) <= cp_elements(362);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(361)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(361),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 362 fork  transition  bypass 
    -- predecessors 367 
    -- successors 360 
    -- marked successors 361 27 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_sample_completed_
      -- 
    cp_elements(362) <= cp_elements(367);
    -- CP-element group 363 join  transition  bypass 
    -- predecessors 365 
    -- marked predecessors 372 390 408 
    -- successors 368 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_update_start_
      -- 
    cpelement_group_363 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(365);
      marked_predecessors(0) <= cp_elements(372);
      marked_predecessors(1) <= cp_elements(390);
      marked_predecessors(2) <= cp_elements(408);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(363)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(363),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 364 transition  bypass 
    -- predecessors 369 
    -- successors 360 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_update_completed_
      -- 
    cp_elements(364) <= cp_elements(369);
    -- CP-element group 365 fork  transition  bypass 
    -- predecessors 24 
    -- successors 361 363 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_518_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_518_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_518_completed_
      -- 
    cp_elements(365) <= cp_elements(24);
    -- CP-element group 366 transition  output  bypass 
    -- predecessors 361 
    -- successors 367 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Sample/rr
      -- 
    cp_elements(366) <= cp_elements(361);
    rr_2091_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(366), ack => binary_521_inst_req_0); -- 
    -- CP-element group 367 transition  input  bypass 
    -- predecessors 366 
    -- successors 362 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Sample/ra
      -- 
    ra_2092_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_521_inst_ack_0, ack => cp_elements(367)); -- 
    -- CP-element group 368 transition  output  bypass 
    -- predecessors 363 
    -- successors 369 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Update/cr
      -- 
    cp_elements(368) <= cp_elements(363);
    cr_2096_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(368), ack => binary_521_inst_req_1); -- 
    -- CP-element group 369 transition  input  bypass 
    -- predecessors 368 
    -- successors 364 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_521_Update/ca
      -- 
    ca_2097_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_521_inst_ack_1, ack => cp_elements(369)); -- 
    -- CP-element group 370 transition  bypass 
    -- predecessors 7 
    -- successors 371 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_trigger_
      -- 
    cp_elements(370) <= cp_elements(7);
    -- CP-element group 371 join  transition  bypass 
    -- predecessors 370 373 
    -- marked predecessors 951 
    -- successors 386 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_active_
      -- 
    cpelement_group_371 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(370);
      predecessors(1) <= cp_elements(373);
      marked_predecessors(0) <= cp_elements(951);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(371)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(371),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 372 join  fork  transition  bypass 
    -- predecessors 387 
    -- marked predecessors 954 
    -- successors 952 
    -- marked successors 363 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_527_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_527_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_527_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_717_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_717_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_717_completed_
      -- 
    cpelement_group_372 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(387);
      marked_predecessors(0) <= cp_elements(954);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(372)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(372),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 373 transition  bypass 
    -- predecessors 385 
    -- successors 371 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_root_address_calculated
      -- 
    cp_elements(373) <= cp_elements(385);
    -- CP-element group 374 transition  bypass 
    -- predecessors 381 
    -- successors 382 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_indices_scaled
      -- 
    cp_elements(374) <= cp_elements(381);
    -- CP-element group 375 transition  bypass 
    -- predecessors 383 
    -- successors 384 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_offset_calculated
      -- 
    cp_elements(375) <= cp_elements(383);
    -- CP-element group 376 transition  bypass 
    -- predecessors 379 
    -- successors 380 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_resized_0
      -- 
    cp_elements(376) <= cp_elements(379);
    -- CP-element group 377 transition  bypass 
    -- predecessors 360 
    -- successors 378 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_524_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_524_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_524_completed_
      -- 
    cp_elements(377) <= cp_elements(360);
    -- CP-element group 378 transition  output  bypass 
    -- predecessors 377 
    -- successors 379 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_resize_0/index_resize_req
      -- 
    cp_elements(378) <= cp_elements(377);
    index_resize_req_2115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(378), ack => array_obj_ref_525_index_0_resize_req_0); -- 
    -- CP-element group 379 transition  input  bypass 
    -- predecessors 378 
    -- successors 376 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_525_index_0_resize_ack_0, ack => cp_elements(379)); -- 
    -- CP-element group 380 transition  output  bypass 
    -- predecessors 376 
    -- successors 381 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_scale_0/scale_rename_req
      -- 
    cp_elements(380) <= cp_elements(376);
    scale_rename_req_2120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(380), ack => array_obj_ref_525_index_0_rename_req_0); -- 
    -- CP-element group 381 transition  input  bypass 
    -- predecessors 380 
    -- successors 374 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_525_index_0_rename_ack_0, ack => cp_elements(381)); -- 
    -- CP-element group 382 transition  output  bypass 
    -- predecessors 374 
    -- successors 383 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_add_indices/final_index_req
      -- 
    cp_elements(382) <= cp_elements(374);
    final_index_req_2125_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(382), ack => array_obj_ref_525_offset_inst_req_0); -- 
    -- CP-element group 383 transition  input  bypass 
    -- predecessors 382 
    -- successors 375 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_add_indices/final_index_ack
      -- 
    final_index_ack_2126_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_525_offset_inst_ack_0, ack => cp_elements(383)); -- 
    -- CP-element group 384 transition  output  bypass 
    -- predecessors 375 
    -- successors 385 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_base_plus_offset/sum_rename_req
      -- 
    cp_elements(384) <= cp_elements(375);
    sum_rename_req_2130_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(384), ack => array_obj_ref_525_root_address_inst_req_0); -- 
    -- CP-element group 385 transition  input  bypass 
    -- predecessors 384 
    -- successors 373 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_525_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2131_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_525_root_address_inst_ack_0, ack => cp_elements(385)); -- 
    -- CP-element group 386 transition  output  bypass 
    -- predecessors 371 
    -- successors 387 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_complete/final_reg_req
      -- 
    cp_elements(386) <= cp_elements(371);
    final_reg_req_2135_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(386), ack => addr_of_526_final_reg_req_0); -- 
    -- CP-element group 387 transition  input  bypass 
    -- predecessors 386 
    -- successors 372 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_526_complete/final_reg_ack
      -- 
    final_reg_ack_2136_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_526_final_reg_ack_0, ack => cp_elements(387)); -- 
    -- CP-element group 388 transition  bypass 
    -- predecessors 7 
    -- successors 389 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_trigger_
      -- 
    cp_elements(388) <= cp_elements(7);
    -- CP-element group 389 join  transition  bypass 
    -- predecessors 388 391 
    -- marked predecessors 645 
    -- successors 404 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_active_
      -- 
    cpelement_group_389 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(388);
      predecessors(1) <= cp_elements(391);
      marked_predecessors(0) <= cp_elements(645);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(389)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(389),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 390 fork  transition  bypass 
    -- predecessors 405 
    -- successors 650 
    -- marked successors 363 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_532_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_532_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_532_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_605_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_605_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_605_completed_
      -- 
    cp_elements(390) <= cp_elements(405);
    -- CP-element group 391 transition  bypass 
    -- predecessors 403 
    -- successors 389 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_root_address_calculated
      -- 
    cp_elements(391) <= cp_elements(403);
    -- CP-element group 392 transition  bypass 
    -- predecessors 399 
    -- successors 400 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_indices_scaled
      -- 
    cp_elements(392) <= cp_elements(399);
    -- CP-element group 393 transition  bypass 
    -- predecessors 401 
    -- successors 402 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_offset_calculated
      -- 
    cp_elements(393) <= cp_elements(401);
    -- CP-element group 394 transition  bypass 
    -- predecessors 397 
    -- successors 398 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_resized_0
      -- 
    cp_elements(394) <= cp_elements(397);
    -- CP-element group 395 transition  bypass 
    -- predecessors 360 
    -- successors 396 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_529_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_529_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_529_completed_
      -- 
    cp_elements(395) <= cp_elements(360);
    -- CP-element group 396 transition  output  bypass 
    -- predecessors 395 
    -- successors 397 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_resize_0/index_resize_req
      -- 
    cp_elements(396) <= cp_elements(395);
    index_resize_req_2154_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(396), ack => array_obj_ref_530_index_0_resize_req_0); -- 
    -- CP-element group 397 transition  input  bypass 
    -- predecessors 396 
    -- successors 394 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2155_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_530_index_0_resize_ack_0, ack => cp_elements(397)); -- 
    -- CP-element group 398 transition  output  bypass 
    -- predecessors 394 
    -- successors 399 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_scale_0/scale_rename_req
      -- 
    cp_elements(398) <= cp_elements(394);
    scale_rename_req_2159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(398), ack => array_obj_ref_530_index_0_rename_req_0); -- 
    -- CP-element group 399 transition  input  bypass 
    -- predecessors 398 
    -- successors 392 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_530_index_0_rename_ack_0, ack => cp_elements(399)); -- 
    -- CP-element group 400 transition  output  bypass 
    -- predecessors 392 
    -- successors 401 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_add_indices/final_index_req
      -- 
    cp_elements(400) <= cp_elements(392);
    final_index_req_2164_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(400), ack => array_obj_ref_530_offset_inst_req_0); -- 
    -- CP-element group 401 transition  input  bypass 
    -- predecessors 400 
    -- successors 393 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_add_indices/final_index_ack
      -- 
    final_index_ack_2165_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_530_offset_inst_ack_0, ack => cp_elements(401)); -- 
    -- CP-element group 402 transition  output  bypass 
    -- predecessors 393 
    -- successors 403 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_base_plus_offset/sum_rename_req
      -- 
    cp_elements(402) <= cp_elements(393);
    sum_rename_req_2169_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(402), ack => array_obj_ref_530_root_address_inst_req_0); -- 
    -- CP-element group 403 transition  input  bypass 
    -- predecessors 402 
    -- successors 391 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_530_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2170_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_530_root_address_inst_ack_0, ack => cp_elements(403)); -- 
    -- CP-element group 404 transition  output  bypass 
    -- predecessors 389 
    -- successors 405 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_complete/final_reg_req
      -- 
    cp_elements(404) <= cp_elements(389);
    final_reg_req_2174_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(404), ack => addr_of_531_final_reg_req_0); -- 
    -- CP-element group 405 transition  input  bypass 
    -- predecessors 404 
    -- successors 390 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_531_complete/final_reg_ack
      -- 
    final_reg_ack_2175_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_531_final_reg_ack_0, ack => cp_elements(405)); -- 
    -- CP-element group 406 transition  bypass 
    -- predecessors 7 
    -- successors 407 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_trigger_
      -- 
    cp_elements(406) <= cp_elements(7);
    -- CP-element group 407 join  transition  bypass 
    -- predecessors 406 409 
    -- marked predecessors 629 
    -- successors 422 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_active_
      -- 
    cpelement_group_407 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(406);
      predecessors(1) <= cp_elements(409);
      marked_predecessors(0) <= cp_elements(629);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(407)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(407),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 408 fork  transition  bypass 
    -- predecessors 423 
    -- successors 634 
    -- marked successors 363 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_537_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_537_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_537_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_601_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_601_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_601_completed_
      -- 
    cp_elements(408) <= cp_elements(423);
    -- CP-element group 409 transition  bypass 
    -- predecessors 421 
    -- successors 407 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_root_address_calculated
      -- 
    cp_elements(409) <= cp_elements(421);
    -- CP-element group 410 transition  bypass 
    -- predecessors 417 
    -- successors 418 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_indices_scaled
      -- 
    cp_elements(410) <= cp_elements(417);
    -- CP-element group 411 transition  bypass 
    -- predecessors 419 
    -- successors 420 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_offset_calculated
      -- 
    cp_elements(411) <= cp_elements(419);
    -- CP-element group 412 transition  bypass 
    -- predecessors 415 
    -- successors 416 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_resized_0
      -- 
    cp_elements(412) <= cp_elements(415);
    -- CP-element group 413 transition  bypass 
    -- predecessors 360 
    -- successors 414 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_534_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_534_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_534_completed_
      -- 
    cp_elements(413) <= cp_elements(360);
    -- CP-element group 414 transition  output  bypass 
    -- predecessors 413 
    -- successors 415 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_resize_0/index_resize_req
      -- 
    cp_elements(414) <= cp_elements(413);
    index_resize_req_2193_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(414), ack => array_obj_ref_535_index_0_resize_req_0); -- 
    -- CP-element group 415 transition  input  bypass 
    -- predecessors 414 
    -- successors 412 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_535_index_0_resize_ack_0, ack => cp_elements(415)); -- 
    -- CP-element group 416 transition  output  bypass 
    -- predecessors 412 
    -- successors 417 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_scale_0/scale_rename_req
      -- 
    cp_elements(416) <= cp_elements(412);
    scale_rename_req_2198_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(416), ack => array_obj_ref_535_index_0_rename_req_0); -- 
    -- CP-element group 417 transition  input  bypass 
    -- predecessors 416 
    -- successors 410 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2199_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_535_index_0_rename_ack_0, ack => cp_elements(417)); -- 
    -- CP-element group 418 transition  output  bypass 
    -- predecessors 410 
    -- successors 419 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_add_indices/final_index_req
      -- 
    cp_elements(418) <= cp_elements(410);
    final_index_req_2203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(418), ack => array_obj_ref_535_offset_inst_req_0); -- 
    -- CP-element group 419 transition  input  bypass 
    -- predecessors 418 
    -- successors 411 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_add_indices/final_index_ack
      -- 
    final_index_ack_2204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_535_offset_inst_ack_0, ack => cp_elements(419)); -- 
    -- CP-element group 420 transition  output  bypass 
    -- predecessors 411 
    -- successors 421 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_base_plus_offset/sum_rename_req
      -- 
    cp_elements(420) <= cp_elements(411);
    sum_rename_req_2208_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(420), ack => array_obj_ref_535_root_address_inst_req_0); -- 
    -- CP-element group 421 transition  input  bypass 
    -- predecessors 420 
    -- successors 409 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_535_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2209_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_535_root_address_inst_ack_0, ack => cp_elements(421)); -- 
    -- CP-element group 422 transition  output  bypass 
    -- predecessors 407 
    -- successors 423 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_complete/final_reg_req
      -- 
    cp_elements(422) <= cp_elements(407);
    final_reg_req_2213_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(422), ack => addr_of_536_final_reg_req_0); -- 
    -- CP-element group 423 transition  input  bypass 
    -- predecessors 422 
    -- successors 408 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_536_complete/final_reg_ack
      -- 
    final_reg_ack_2214_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_536_final_reg_ack_0, ack => cp_elements(423)); -- 
    -- CP-element group 424 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_active_
      -- 
    cp_elements(424) <= cp_elements(7);
    -- CP-element group 425 join  fork  transition  bypass 
    -- predecessors 427 429 
    -- successors 442 460 478 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_543_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_543_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_543_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_completed_
      -- 
    cpelement_group_425 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(427);
      predecessors(1) <= cp_elements(429);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(425)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(425),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 426 join  transition  bypass 
    -- predecessors 430 
    -- marked predecessors 427 
    -- successors 431 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_sample_start_
      -- 
    cpelement_group_426 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(430);
      marked_predecessors(0) <= cp_elements(427);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(426)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(426),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 427 fork  transition  bypass 
    -- predecessors 432 
    -- successors 425 
    -- marked successors 27 426 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_sample_completed_
      -- 
    cp_elements(427) <= cp_elements(432);
    -- CP-element group 428 join  transition  bypass 
    -- predecessors 430 
    -- marked predecessors 437 455 473 
    -- successors 433 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_update_start_
      -- 
    cpelement_group_428 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(2 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(430);
      marked_predecessors(0) <= cp_elements(437);
      marked_predecessors(1) <= cp_elements(455);
      marked_predecessors(2) <= cp_elements(473);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(428)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(428),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 429 transition  bypass 
    -- predecessors 434 
    -- successors 425 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_update_completed_
      -- 
    cp_elements(429) <= cp_elements(434);
    -- CP-element group 430 fork  transition  bypass 
    -- predecessors 24 
    -- successors 426 428 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_539_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_539_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_539_completed_
      -- 
    cp_elements(430) <= cp_elements(24);
    -- CP-element group 431 transition  output  bypass 
    -- predecessors 426 
    -- successors 432 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Sample/rr
      -- 
    cp_elements(431) <= cp_elements(426);
    rr_2231_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(431), ack => binary_542_inst_req_0); -- 
    -- CP-element group 432 transition  input  bypass 
    -- predecessors 431 
    -- successors 427 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Sample/ra
      -- 
    ra_2232_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_542_inst_ack_0, ack => cp_elements(432)); -- 
    -- CP-element group 433 transition  output  bypass 
    -- predecessors 428 
    -- successors 434 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Update/cr
      -- 
    cp_elements(433) <= cp_elements(428);
    cr_2236_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(433), ack => binary_542_inst_req_1); -- 
    -- CP-element group 434 transition  input  bypass 
    -- predecessors 433 
    -- successors 429 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_542_Update/ca
      -- 
    ca_2237_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_542_inst_ack_1, ack => cp_elements(434)); -- 
    -- CP-element group 435 transition  bypass 
    -- predecessors 7 
    -- successors 436 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_trigger_
      -- 
    cp_elements(435) <= cp_elements(7);
    -- CP-element group 436 join  transition  bypass 
    -- predecessors 435 438 
    -- marked predecessors 919 
    -- successors 451 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_active_
      -- 
    cpelement_group_436 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(435);
      predecessors(1) <= cp_elements(438);
      marked_predecessors(0) <= cp_elements(919);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(436)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(436),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 437 join  fork  transition  bypass 
    -- predecessors 452 
    -- marked predecessors 922 
    -- successors 920 
    -- marked successors 428 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_548_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_548_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_548_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_698_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_698_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_698_completed_
      -- 
    cpelement_group_437 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(452);
      marked_predecessors(0) <= cp_elements(922);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(437)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(437),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 438 transition  bypass 
    -- predecessors 450 
    -- successors 436 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_root_address_calculated
      -- 
    cp_elements(438) <= cp_elements(450);
    -- CP-element group 439 transition  bypass 
    -- predecessors 446 
    -- successors 447 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_indices_scaled
      -- 
    cp_elements(439) <= cp_elements(446);
    -- CP-element group 440 transition  bypass 
    -- predecessors 448 
    -- successors 449 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_offset_calculated
      -- 
    cp_elements(440) <= cp_elements(448);
    -- CP-element group 441 transition  bypass 
    -- predecessors 444 
    -- successors 445 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_resized_0
      -- 
    cp_elements(441) <= cp_elements(444);
    -- CP-element group 442 transition  bypass 
    -- predecessors 425 
    -- successors 443 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_545_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_545_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_545_completed_
      -- 
    cp_elements(442) <= cp_elements(425);
    -- CP-element group 443 transition  output  bypass 
    -- predecessors 442 
    -- successors 444 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_resize_0/index_resize_req
      -- 
    cp_elements(443) <= cp_elements(442);
    index_resize_req_2255_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(443), ack => array_obj_ref_546_index_0_resize_req_0); -- 
    -- CP-element group 444 transition  input  bypass 
    -- predecessors 443 
    -- successors 441 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2256_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_546_index_0_resize_ack_0, ack => cp_elements(444)); -- 
    -- CP-element group 445 transition  output  bypass 
    -- predecessors 441 
    -- successors 446 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_scale_0/scale_rename_req
      -- 
    cp_elements(445) <= cp_elements(441);
    scale_rename_req_2260_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(445), ack => array_obj_ref_546_index_0_rename_req_0); -- 
    -- CP-element group 446 transition  input  bypass 
    -- predecessors 445 
    -- successors 439 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2261_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_546_index_0_rename_ack_0, ack => cp_elements(446)); -- 
    -- CP-element group 447 transition  output  bypass 
    -- predecessors 439 
    -- successors 448 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_add_indices/final_index_req
      -- 
    cp_elements(447) <= cp_elements(439);
    final_index_req_2265_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(447), ack => array_obj_ref_546_offset_inst_req_0); -- 
    -- CP-element group 448 transition  input  bypass 
    -- predecessors 447 
    -- successors 440 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_add_indices/final_index_ack
      -- 
    final_index_ack_2266_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_546_offset_inst_ack_0, ack => cp_elements(448)); -- 
    -- CP-element group 449 transition  output  bypass 
    -- predecessors 440 
    -- successors 450 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_base_plus_offset/sum_rename_req
      -- 
    cp_elements(449) <= cp_elements(440);
    sum_rename_req_2270_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(449), ack => array_obj_ref_546_root_address_inst_req_0); -- 
    -- CP-element group 450 transition  input  bypass 
    -- predecessors 449 
    -- successors 438 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_546_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2271_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_546_root_address_inst_ack_0, ack => cp_elements(450)); -- 
    -- CP-element group 451 transition  output  bypass 
    -- predecessors 436 
    -- successors 452 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_complete/final_reg_req
      -- 
    cp_elements(451) <= cp_elements(436);
    final_reg_req_2275_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(451), ack => addr_of_547_final_reg_req_0); -- 
    -- CP-element group 452 transition  input  bypass 
    -- predecessors 451 
    -- successors 437 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_547_complete/final_reg_ack
      -- 
    final_reg_ack_2276_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_547_final_reg_ack_0, ack => cp_elements(452)); -- 
    -- CP-element group 453 transition  bypass 
    -- predecessors 7 
    -- successors 454 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_trigger_
      -- 
    cp_elements(453) <= cp_elements(7);
    -- CP-element group 454 join  transition  bypass 
    -- predecessors 453 456 
    -- marked predecessors 602 
    -- successors 469 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_active_
      -- 
    cpelement_group_454 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(453);
      predecessors(1) <= cp_elements(456);
      marked_predecessors(0) <= cp_elements(602);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(454)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(454),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 455 fork  transition  bypass 
    -- predecessors 470 
    -- successors 607 
    -- marked successors 428 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_553_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_553_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_553_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_592_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_592_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_592_completed_
      -- 
    cp_elements(455) <= cp_elements(470);
    -- CP-element group 456 transition  bypass 
    -- predecessors 468 
    -- successors 454 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_root_address_calculated
      -- 
    cp_elements(456) <= cp_elements(468);
    -- CP-element group 457 transition  bypass 
    -- predecessors 464 
    -- successors 465 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_indices_scaled
      -- 
    cp_elements(457) <= cp_elements(464);
    -- CP-element group 458 transition  bypass 
    -- predecessors 466 
    -- successors 467 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_offset_calculated
      -- 
    cp_elements(458) <= cp_elements(466);
    -- CP-element group 459 transition  bypass 
    -- predecessors 462 
    -- successors 463 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_resized_0
      -- 
    cp_elements(459) <= cp_elements(462);
    -- CP-element group 460 transition  bypass 
    -- predecessors 425 
    -- successors 461 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_550_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_550_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_550_completed_
      -- 
    cp_elements(460) <= cp_elements(425);
    -- CP-element group 461 transition  output  bypass 
    -- predecessors 460 
    -- successors 462 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_resize_0/index_resize_req
      -- 
    cp_elements(461) <= cp_elements(460);
    index_resize_req_2294_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(461), ack => array_obj_ref_551_index_0_resize_req_0); -- 
    -- CP-element group 462 transition  input  bypass 
    -- predecessors 461 
    -- successors 459 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2295_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_551_index_0_resize_ack_0, ack => cp_elements(462)); -- 
    -- CP-element group 463 transition  output  bypass 
    -- predecessors 459 
    -- successors 464 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_scale_0/scale_rename_req
      -- 
    cp_elements(463) <= cp_elements(459);
    scale_rename_req_2299_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(463), ack => array_obj_ref_551_index_0_rename_req_0); -- 
    -- CP-element group 464 transition  input  bypass 
    -- predecessors 463 
    -- successors 457 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2300_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_551_index_0_rename_ack_0, ack => cp_elements(464)); -- 
    -- CP-element group 465 transition  output  bypass 
    -- predecessors 457 
    -- successors 466 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_add_indices/$entry
      -- 
    cp_elements(465) <= cp_elements(457);
    final_index_req_2304_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(465), ack => array_obj_ref_551_offset_inst_req_0); -- 
    -- CP-element group 466 transition  input  bypass 
    -- predecessors 465 
    -- successors 458 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_add_indices/final_index_ack
      -- 
    final_index_ack_2305_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_551_offset_inst_ack_0, ack => cp_elements(466)); -- 
    -- CP-element group 467 transition  output  bypass 
    -- predecessors 458 
    -- successors 468 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_base_plus_offset/sum_rename_req
      -- 
    cp_elements(467) <= cp_elements(458);
    sum_rename_req_2309_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(467), ack => array_obj_ref_551_root_address_inst_req_0); -- 
    -- CP-element group 468 transition  input  bypass 
    -- predecessors 467 
    -- successors 456 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_551_base_plus_offset/$exit
      -- 
    sum_rename_ack_2310_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_551_root_address_inst_ack_0, ack => cp_elements(468)); -- 
    -- CP-element group 469 transition  output  bypass 
    -- predecessors 454 
    -- successors 470 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_complete/final_reg_req
      -- 
    cp_elements(469) <= cp_elements(454);
    final_reg_req_2314_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(469), ack => addr_of_552_final_reg_req_0); -- 
    -- CP-element group 470 transition  input  bypass 
    -- predecessors 469 
    -- successors 455 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_552_complete/final_reg_ack
      -- 
    final_reg_ack_2315_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_552_final_reg_ack_0, ack => cp_elements(470)); -- 
    -- CP-element group 471 transition  bypass 
    -- predecessors 7 
    -- successors 472 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_trigger_
      -- 
    cp_elements(471) <= cp_elements(7);
    -- CP-element group 472 join  transition  bypass 
    -- predecessors 471 474 
    -- marked predecessors 586 
    -- successors 487 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_active_
      -- 
    cpelement_group_472 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(471);
      predecessors(1) <= cp_elements(474);
      marked_predecessors(0) <= cp_elements(586);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(472)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(472),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 473 fork  transition  bypass 
    -- predecessors 488 
    -- successors 591 
    -- marked successors 428 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_558_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_558_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_558_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_588_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_588_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_588_completed_
      -- 
    cp_elements(473) <= cp_elements(488);
    -- CP-element group 474 transition  bypass 
    -- predecessors 486 
    -- successors 472 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_root_address_calculated
      -- 
    cp_elements(474) <= cp_elements(486);
    -- CP-element group 475 transition  bypass 
    -- predecessors 482 
    -- successors 483 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_indices_scaled
      -- 
    cp_elements(475) <= cp_elements(482);
    -- CP-element group 476 transition  bypass 
    -- predecessors 484 
    -- successors 485 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_offset_calculated
      -- 
    cp_elements(476) <= cp_elements(484);
    -- CP-element group 477 transition  bypass 
    -- predecessors 480 
    -- successors 481 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_resized_0
      -- 
    cp_elements(477) <= cp_elements(480);
    -- CP-element group 478 transition  bypass 
    -- predecessors 425 
    -- successors 479 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_555_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_555_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_555_active_
      -- 
    cp_elements(478) <= cp_elements(425);
    -- CP-element group 479 transition  output  bypass 
    -- predecessors 478 
    -- successors 480 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_resize_0/index_resize_req
      -- 
    cp_elements(479) <= cp_elements(478);
    index_resize_req_2333_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(479), ack => array_obj_ref_556_index_0_resize_req_0); -- 
    -- CP-element group 480 transition  input  bypass 
    -- predecessors 479 
    -- successors 477 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2334_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_556_index_0_resize_ack_0, ack => cp_elements(480)); -- 
    -- CP-element group 481 transition  output  bypass 
    -- predecessors 477 
    -- successors 482 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_scale_0/scale_rename_req
      -- 
    cp_elements(481) <= cp_elements(477);
    scale_rename_req_2338_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(481), ack => array_obj_ref_556_index_0_rename_req_0); -- 
    -- CP-element group 482 transition  input  bypass 
    -- predecessors 481 
    -- successors 475 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_index_scale_0/$exit
      -- 
    scale_rename_ack_2339_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_556_index_0_rename_ack_0, ack => cp_elements(482)); -- 
    -- CP-element group 483 transition  output  bypass 
    -- predecessors 475 
    -- successors 484 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_add_indices/$entry
      -- 
    cp_elements(483) <= cp_elements(475);
    final_index_req_2343_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(483), ack => array_obj_ref_556_offset_inst_req_0); -- 
    -- CP-element group 484 transition  input  bypass 
    -- predecessors 483 
    -- successors 476 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_add_indices/final_index_ack
      -- 
    final_index_ack_2344_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_556_offset_inst_ack_0, ack => cp_elements(484)); -- 
    -- CP-element group 485 transition  output  bypass 
    -- predecessors 476 
    -- successors 486 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_base_plus_offset/sum_rename_req
      -- 
    cp_elements(485) <= cp_elements(476);
    sum_rename_req_2348_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(485), ack => array_obj_ref_556_root_address_inst_req_0); -- 
    -- CP-element group 486 transition  input  bypass 
    -- predecessors 485 
    -- successors 474 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_556_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2349_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_556_root_address_inst_ack_0, ack => cp_elements(486)); -- 
    -- CP-element group 487 transition  output  bypass 
    -- predecessors 472 
    -- successors 488 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_complete/final_reg_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_complete/$entry
      -- 
    cp_elements(487) <= cp_elements(472);
    final_reg_req_2353_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(487), ack => addr_of_557_final_reg_req_0); -- 
    -- CP-element group 488 transition  input  bypass 
    -- predecessors 487 
    -- successors 473 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_complete/final_reg_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_557_complete/$exit
      -- 
    final_reg_ack_2354_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_557_final_reg_ack_0, ack => cp_elements(488)); -- 
    -- CP-element group 489 transition  bypass 
    -- predecessors 7 
    -- successors 490 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_trigger_
      -- 
    cp_elements(489) <= cp_elements(7);
    -- CP-element group 490 join  transition  bypass 
    -- predecessors 489 492 
    -- marked predecessors 887 
    -- successors 505 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_active_
      -- 
    cpelement_group_490 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(489);
      predecessors(1) <= cp_elements(492);
      marked_predecessors(0) <= cp_elements(887);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(490)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(490),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 491 join  fork  transition  bypass 
    -- predecessors 506 
    -- marked predecessors 890 
    -- successors 888 
    -- marked successors 27 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_563_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_563_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_563_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_679_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_679_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_679_completed_
      -- 
    cpelement_group_491 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(506);
      marked_predecessors(0) <= cp_elements(890);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(491)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(491),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 492 transition  bypass 
    -- predecessors 504 
    -- successors 490 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_root_address_calculated
      -- 
    cp_elements(492) <= cp_elements(504);
    -- CP-element group 493 transition  bypass 
    -- predecessors 500 
    -- successors 501 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_indices_scaled
      -- 
    cp_elements(493) <= cp_elements(500);
    -- CP-element group 494 transition  bypass 
    -- predecessors 502 
    -- successors 503 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_offset_calculated
      -- 
    cp_elements(494) <= cp_elements(502);
    -- CP-element group 495 transition  bypass 
    -- predecessors 498 
    -- successors 499 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_resized_0
      -- 
    cp_elements(495) <= cp_elements(498);
    -- CP-element group 496 transition  bypass 
    -- predecessors 24 
    -- successors 497 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_560_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_560_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_560_completed_
      -- 
    cp_elements(496) <= cp_elements(24);
    -- CP-element group 497 transition  output  bypass 
    -- predecessors 496 
    -- successors 498 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_resize_0/index_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_resize_0/$entry
      -- 
    cp_elements(497) <= cp_elements(496);
    index_resize_req_2372_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(497), ack => array_obj_ref_561_index_0_resize_req_0); -- 
    -- CP-element group 498 transition  input  bypass 
    -- predecessors 497 
    -- successors 495 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_resize_0/$exit
      -- 
    index_resize_ack_2373_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_index_0_resize_ack_0, ack => cp_elements(498)); -- 
    -- CP-element group 499 transition  output  bypass 
    -- predecessors 495 
    -- successors 500 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_scale_0/scale_rename_req
      -- 
    cp_elements(499) <= cp_elements(495);
    scale_rename_req_2377_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(499), ack => array_obj_ref_561_index_0_rename_req_0); -- 
    -- CP-element group 500 transition  input  bypass 
    -- predecessors 499 
    -- successors 493 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_scale_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_index_scale_0/scale_rename_ack
      -- 
    scale_rename_ack_2378_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_index_0_rename_ack_0, ack => cp_elements(500)); -- 
    -- CP-element group 501 transition  output  bypass 
    -- predecessors 493 
    -- successors 502 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_add_indices/$entry
      -- 
    cp_elements(501) <= cp_elements(493);
    final_index_req_2382_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(501), ack => array_obj_ref_561_offset_inst_req_0); -- 
    -- CP-element group 502 transition  input  bypass 
    -- predecessors 501 
    -- successors 494 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_add_indices/final_index_ack
      -- 
    final_index_ack_2383_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_offset_inst_ack_0, ack => cp_elements(502)); -- 
    -- CP-element group 503 transition  output  bypass 
    -- predecessors 494 
    -- successors 504 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_base_plus_offset/sum_rename_req
      -- 
    cp_elements(503) <= cp_elements(494);
    sum_rename_req_2387_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(503), ack => array_obj_ref_561_root_address_inst_req_0); -- 
    -- CP-element group 504 transition  input  bypass 
    -- predecessors 503 
    -- successors 492 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_561_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2388_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_561_root_address_inst_ack_0, ack => cp_elements(504)); -- 
    -- CP-element group 505 transition  output  bypass 
    -- predecessors 490 
    -- successors 506 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_complete/final_reg_req
      -- 
    cp_elements(505) <= cp_elements(490);
    final_reg_req_2392_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(505), ack => addr_of_562_final_reg_req_0); -- 
    -- CP-element group 506 transition  input  bypass 
    -- predecessors 505 
    -- successors 491 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_562_complete/final_reg_ack
      -- 
    final_reg_ack_2393_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_562_final_reg_ack_0, ack => cp_elements(506)); -- 
    -- CP-element group 507 transition  bypass 
    -- predecessors 7 
    -- successors 508 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_trigger_
      -- 
    cp_elements(507) <= cp_elements(7);
    -- CP-element group 508 join  transition  bypass 
    -- predecessors 507 510 
    -- marked predecessors 559 
    -- successors 523 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_active_
      -- 
    cpelement_group_508 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(507);
      predecessors(1) <= cp_elements(510);
      marked_predecessors(0) <= cp_elements(559);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(508)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(508),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 509 fork  transition  bypass 
    -- predecessors 524 
    -- successors 564 
    -- marked successors 27 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_568_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_568_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_568_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_579_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_579_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_579_completed_
      -- 
    cp_elements(509) <= cp_elements(524);
    -- CP-element group 510 transition  bypass 
    -- predecessors 522 
    -- successors 508 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_root_address_calculated
      -- 
    cp_elements(510) <= cp_elements(522);
    -- CP-element group 511 transition  bypass 
    -- predecessors 518 
    -- successors 519 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_indices_scaled
      -- 
    cp_elements(511) <= cp_elements(518);
    -- CP-element group 512 transition  bypass 
    -- predecessors 520 
    -- successors 521 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_offset_calculated
      -- 
    cp_elements(512) <= cp_elements(520);
    -- CP-element group 513 transition  bypass 
    -- predecessors 516 
    -- successors 517 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_resized_0
      -- 
    cp_elements(513) <= cp_elements(516);
    -- CP-element group 514 transition  bypass 
    -- predecessors 24 
    -- successors 515 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_565_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_565_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_565_active_
      -- 
    cp_elements(514) <= cp_elements(24);
    -- CP-element group 515 transition  output  bypass 
    -- predecessors 514 
    -- successors 516 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_resize_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_resize_0/index_resize_req
      -- 
    cp_elements(515) <= cp_elements(514);
    index_resize_req_2411_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(515), ack => array_obj_ref_566_index_0_resize_req_0); -- 
    -- CP-element group 516 transition  input  bypass 
    -- predecessors 515 
    -- successors 513 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_resize_0/index_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_resize_0/$exit
      -- 
    index_resize_ack_2412_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_566_index_0_resize_ack_0, ack => cp_elements(516)); -- 
    -- CP-element group 517 transition  output  bypass 
    -- predecessors 513 
    -- successors 518 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_scale_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_scale_0/scale_rename_req
      -- 
    cp_elements(517) <= cp_elements(513);
    scale_rename_req_2416_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(517), ack => array_obj_ref_566_index_0_rename_req_0); -- 
    -- CP-element group 518 transition  input  bypass 
    -- predecessors 517 
    -- successors 511 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_index_scale_0/$exit
      -- 
    scale_rename_ack_2417_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_566_index_0_rename_ack_0, ack => cp_elements(518)); -- 
    -- CP-element group 519 transition  output  bypass 
    -- predecessors 511 
    -- successors 520 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_add_indices/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_add_indices/final_index_req
      -- 
    cp_elements(519) <= cp_elements(511);
    final_index_req_2421_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(519), ack => array_obj_ref_566_offset_inst_req_0); -- 
    -- CP-element group 520 transition  input  bypass 
    -- predecessors 519 
    -- successors 512 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_add_indices/final_index_ack
      -- 
    final_index_ack_2422_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_566_offset_inst_ack_0, ack => cp_elements(520)); -- 
    -- CP-element group 521 transition  output  bypass 
    -- predecessors 512 
    -- successors 522 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_base_plus_offset/$entry
      -- 
    cp_elements(521) <= cp_elements(512);
    sum_rename_req_2426_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(521), ack => array_obj_ref_566_root_address_inst_req_0); -- 
    -- CP-element group 522 transition  input  bypass 
    -- predecessors 521 
    -- successors 510 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_566_base_plus_offset/$exit
      -- 
    sum_rename_ack_2427_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_566_root_address_inst_ack_0, ack => cp_elements(522)); -- 
    -- CP-element group 523 transition  output  bypass 
    -- predecessors 508 
    -- successors 524 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_complete/final_reg_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_complete/$entry
      -- 
    cp_elements(523) <= cp_elements(508);
    final_reg_req_2431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(523), ack => addr_of_567_final_reg_req_0); -- 
    -- CP-element group 524 transition  input  bypass 
    -- predecessors 523 
    -- successors 509 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_complete/final_reg_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_567_complete/$exit
      -- 
    final_reg_ack_2432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_567_final_reg_ack_0, ack => cp_elements(524)); -- 
    -- CP-element group 525 transition  bypass 
    -- predecessors 7 
    -- successors 526 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_trigger_
      -- 
    cp_elements(525) <= cp_elements(7);
    -- CP-element group 526 join  transition  bypass 
    -- predecessors 525 528 
    -- marked predecessors 543 
    -- successors 541 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_active_
      -- 
    cpelement_group_526 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(525);
      predecessors(1) <= cp_elements(528);
      marked_predecessors(0) <= cp_elements(543);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(526)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(526),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 527 fork  transition  bypass 
    -- predecessors 542 
    -- successors 548 
    -- marked successors 27 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_573_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_573_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_573_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_575_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_575_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_575_completed_
      -- 
    cp_elements(527) <= cp_elements(542);
    -- CP-element group 528 transition  bypass 
    -- predecessors 540 
    -- successors 526 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_root_address_calculated
      -- 
    cp_elements(528) <= cp_elements(540);
    -- CP-element group 529 transition  bypass 
    -- predecessors 536 
    -- successors 537 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_indices_scaled
      -- 
    cp_elements(529) <= cp_elements(536);
    -- CP-element group 530 transition  bypass 
    -- predecessors 538 
    -- successors 539 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_offset_calculated
      -- 
    cp_elements(530) <= cp_elements(538);
    -- CP-element group 531 transition  bypass 
    -- predecessors 534 
    -- successors 535 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_resized_0
      -- 
    cp_elements(531) <= cp_elements(534);
    -- CP-element group 532 transition  bypass 
    -- predecessors 24 
    -- successors 533 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_570_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_570_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_computed_0
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_570_completed_
      -- 
    cp_elements(532) <= cp_elements(24);
    -- CP-element group 533 transition  output  bypass 
    -- predecessors 532 
    -- successors 534 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_resize_0/index_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_resize_0/$entry
      -- 
    cp_elements(533) <= cp_elements(532);
    index_resize_req_2450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(533), ack => array_obj_ref_571_index_0_resize_req_0); -- 
    -- CP-element group 534 transition  input  bypass 
    -- predecessors 533 
    -- successors 531 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_resize_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_resize_0/index_resize_ack
      -- 
    index_resize_ack_2451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_index_0_resize_ack_0, ack => cp_elements(534)); -- 
    -- CP-element group 535 transition  output  bypass 
    -- predecessors 531 
    -- successors 536 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_scale_0/scale_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_scale_0/$entry
      -- 
    cp_elements(535) <= cp_elements(531);
    scale_rename_req_2455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(535), ack => array_obj_ref_571_index_0_rename_req_0); -- 
    -- CP-element group 536 transition  input  bypass 
    -- predecessors 535 
    -- successors 529 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_scale_0/scale_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_index_scale_0/$exit
      -- 
    scale_rename_ack_2456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_index_0_rename_ack_0, ack => cp_elements(536)); -- 
    -- CP-element group 537 transition  output  bypass 
    -- predecessors 529 
    -- successors 538 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_add_indices/final_index_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_add_indices/$entry
      -- 
    cp_elements(537) <= cp_elements(529);
    final_index_req_2460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(537), ack => array_obj_ref_571_offset_inst_req_0); -- 
    -- CP-element group 538 transition  input  bypass 
    -- predecessors 537 
    -- successors 530 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_add_indices/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_add_indices/final_index_ack
      -- 
    final_index_ack_2461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_offset_inst_ack_0, ack => cp_elements(538)); -- 
    -- CP-element group 539 transition  output  bypass 
    -- predecessors 530 
    -- successors 540 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_base_plus_offset/sum_rename_req
      -- 
    cp_elements(539) <= cp_elements(530);
    sum_rename_req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(539), ack => array_obj_ref_571_root_address_inst_req_0); -- 
    -- CP-element group 540 transition  input  bypass 
    -- predecessors 539 
    -- successors 528 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/array_obj_ref_571_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_571_root_address_inst_ack_0, ack => cp_elements(540)); -- 
    -- CP-element group 541 transition  output  bypass 
    -- predecessors 526 
    -- successors 542 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_complete/final_reg_req
      -- 
    cp_elements(541) <= cp_elements(526);
    final_reg_req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(541), ack => addr_of_572_final_reg_req_0); -- 
    -- CP-element group 542 transition  input  bypass 
    -- predecessors 541 
    -- successors 527 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/addr_of_572_complete/final_reg_ack
      -- 
    final_reg_ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => addr_of_572_final_reg_ack_0, ack => cp_elements(542)); -- 
    -- CP-element group 543 join  fork  transition  bypass 
    -- predecessors 555 
    -- marked predecessors 579 
    -- successors 556 
    -- marked successors 526 545 546 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_active_
      -- 
    cpelement_group_543 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(555);
      marked_predecessors(0) <= cp_elements(579);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(543)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(543),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 544 transition  bypass 
    -- predecessors 558 
    -- successors 575 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_577_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_577_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_577_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_583_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_583_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_583_completed_
      -- 
    cp_elements(544) <= cp_elements(558);
    -- CP-element group 545 join  transition  bypass 
    -- predecessors 553 
    -- marked predecessors 543 
    -- successors 554 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_word_address_calculated
      -- 
    cpelement_group_545 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(553);
      marked_predecessors(0) <= cp_elements(543);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(545)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(545),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 546 join  transition  bypass 
    -- predecessors 551 
    -- marked predecessors 543 
    -- successors 552 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_root_address_calculated
      -- 
    cpelement_group_546 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(551);
      marked_predecessors(0) <= cp_elements(543);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(546)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(546),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 547 transition  bypass 
    -- predecessors 549 
    -- successors 550 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_address_resized
      -- 
    cp_elements(547) <= cp_elements(549);
    -- CP-element group 548 transition  output  bypass 
    -- predecessors 527 
    -- successors 549 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_addr_resize/base_resize_req
      -- 
    cp_elements(548) <= cp_elements(527);
    base_resize_req_2488_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(548), ack => ptr_deref_576_base_resize_req_0); -- 
    -- CP-element group 549 transition  input  bypass 
    -- predecessors 548 
    -- successors 547 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2489_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_base_resize_ack_0, ack => cp_elements(549)); -- 
    -- CP-element group 550 transition  output  bypass 
    -- predecessors 547 
    -- successors 551 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_plus_offset/sum_rename_req
      -- 
    cp_elements(550) <= cp_elements(547);
    sum_rename_req_2493_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(550), ack => ptr_deref_576_root_address_inst_req_0); -- 
    -- CP-element group 551 transition  input  bypass 
    -- predecessors 550 
    -- successors 546 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2494_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_root_address_inst_ack_0, ack => cp_elements(551)); -- 
    -- CP-element group 552 transition  output  bypass 
    -- predecessors 546 
    -- successors 553 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_word_addrgen/root_register_req
      -- 
    cp_elements(552) <= cp_elements(546);
    root_register_req_2498_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(552), ack => ptr_deref_576_addr_0_req_0); -- 
    -- CP-element group 553 transition  input  bypass 
    -- predecessors 552 
    -- successors 545 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_word_addrgen/root_register_ack
      -- 
    root_register_ack_2499_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_addr_0_ack_0, ack => cp_elements(553)); -- 
    -- CP-element group 554 transition  output  bypass 
    -- predecessors 545 
    -- successors 555 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/word_access_0/rr
      -- 
    cp_elements(554) <= cp_elements(545);
    rr_2509_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(554), ack => ptr_deref_576_load_0_req_0); -- 
    -- CP-element group 555 transition  input  bypass 
    -- predecessors 554 
    -- successors 543 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_request/word_access/word_access_0/ra
      -- 
    ra_2510_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_load_0_ack_0, ack => cp_elements(555)); -- 
    -- CP-element group 556 transition  output  bypass 
    -- predecessors 543 
    -- successors 557 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/word_access_0/cr
      -- 
    cp_elements(556) <= cp_elements(543);
    cr_2520_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(556), ack => ptr_deref_576_load_0_req_1); -- 
    -- CP-element group 557 transition  input  output  bypass 
    -- predecessors 556 
    -- successors 558 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/merge_req
      -- 
    ca_2521_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_load_0_ack_1, ack => cp_elements(557)); -- 
    merge_req_2522_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(557), ack => ptr_deref_576_gather_scatter_req_0); -- 
    -- CP-element group 558 transition  input  bypass 
    -- predecessors 557 
    -- successors 544 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_576_complete/merge_ack
      -- 
    merge_ack_2523_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_576_gather_scatter_ack_0, ack => cp_elements(558)); -- 
    -- CP-element group 559 join  fork  transition  bypass 
    -- predecessors 571 
    -- marked predecessors 579 
    -- successors 572 
    -- marked successors 508 561 562 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_active_
      -- 
    cpelement_group_559 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(571);
      marked_predecessors(0) <= cp_elements(579);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(559)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(559),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 560 transition  bypass 
    -- predecessors 574 
    -- successors 575 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_581_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_581_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_581_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_584_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_584_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_584_completed_
      -- 
    cp_elements(560) <= cp_elements(574);
    -- CP-element group 561 join  transition  bypass 
    -- predecessors 569 
    -- marked predecessors 559 
    -- successors 570 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_word_address_calculated
      -- 
    cpelement_group_561 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(569);
      marked_predecessors(0) <= cp_elements(559);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(561)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(561),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 562 join  transition  bypass 
    -- predecessors 567 
    -- marked predecessors 559 
    -- successors 568 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_root_address_calculated
      -- 
    cpelement_group_562 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(567);
      marked_predecessors(0) <= cp_elements(559);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(562)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(562),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 563 transition  bypass 
    -- predecessors 565 
    -- successors 566 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_address_resized
      -- 
    cp_elements(563) <= cp_elements(565);
    -- CP-element group 564 transition  output  bypass 
    -- predecessors 509 
    -- successors 565 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_addr_resize/base_resize_req
      -- 
    cp_elements(564) <= cp_elements(509);
    base_resize_req_2540_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(564), ack => ptr_deref_580_base_resize_req_0); -- 
    -- CP-element group 565 transition  input  bypass 
    -- predecessors 564 
    -- successors 563 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2541_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_base_resize_ack_0, ack => cp_elements(565)); -- 
    -- CP-element group 566 transition  output  bypass 
    -- predecessors 563 
    -- successors 567 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_plus_offset/sum_rename_req
      -- 
    cp_elements(566) <= cp_elements(563);
    sum_rename_req_2545_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(566), ack => ptr_deref_580_root_address_inst_req_0); -- 
    -- CP-element group 567 transition  input  bypass 
    -- predecessors 566 
    -- successors 562 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2546_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_root_address_inst_ack_0, ack => cp_elements(567)); -- 
    -- CP-element group 568 transition  output  bypass 
    -- predecessors 562 
    -- successors 569 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_word_addrgen/root_register_req
      -- 
    cp_elements(568) <= cp_elements(562);
    root_register_req_2550_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(568), ack => ptr_deref_580_addr_0_req_0); -- 
    -- CP-element group 569 transition  input  bypass 
    -- predecessors 568 
    -- successors 561 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_word_addrgen/root_register_ack
      -- 
    root_register_ack_2551_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_addr_0_ack_0, ack => cp_elements(569)); -- 
    -- CP-element group 570 transition  output  bypass 
    -- predecessors 561 
    -- successors 571 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/word_access_0/rr
      -- 
    cp_elements(570) <= cp_elements(561);
    rr_2561_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(570), ack => ptr_deref_580_load_0_req_0); -- 
    -- CP-element group 571 transition  input  bypass 
    -- predecessors 570 
    -- successors 559 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_request/word_access/word_access_0/ra
      -- 
    ra_2562_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_load_0_ack_0, ack => cp_elements(571)); -- 
    -- CP-element group 572 transition  output  bypass 
    -- predecessors 559 
    -- successors 573 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/word_access_0/cr
      -- 
    cp_elements(572) <= cp_elements(559);
    cr_2572_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(572), ack => ptr_deref_580_load_0_req_1); -- 
    -- CP-element group 573 transition  input  output  bypass 
    -- predecessors 572 
    -- successors 574 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/merge_req
      -- 
    ca_2573_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_load_0_ack_1, ack => cp_elements(573)); -- 
    merge_req_2574_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(573), ack => ptr_deref_580_gather_scatter_req_0); -- 
    -- CP-element group 574 transition  input  bypass 
    -- predecessors 573 
    -- successors 560 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_580_complete/merge_ack
      -- 
    merge_ack_2575_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_580_gather_scatter_ack_0, ack => cp_elements(574)); -- 
    -- CP-element group 575 join  fork  transition  bypass 
    -- predecessors 544 560 
    -- successors 578 580 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_trigger_
      -- 
    cpelement_group_575 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(544);
      predecessors(1) <= cp_elements(560);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(575)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(575),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 576 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_active_
      -- 
    cp_elements(576) <= cp_elements(7);
    -- CP-element group 577 join  transition  bypass 
    -- predecessors 579 581 
    -- successors 902 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_586_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_586_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_586_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_696_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_696_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_695_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_695_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_695_completed_
      -- 
    cpelement_group_577 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(579);
      predecessors(1) <= cp_elements(581);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(577)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(577),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 578 join  transition  bypass 
    -- predecessors 575 
    -- marked predecessors 579 
    -- successors 582 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_sample_start_
      -- 
    cpelement_group_578 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(575);
      marked_predecessors(0) <= cp_elements(579);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(578)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(578),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 579 fork  transition  bypass 
    -- predecessors 583 
    -- successors 577 
    -- marked successors 543 559 578 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_sample_completed_
      -- 
    cp_elements(579) <= cp_elements(583);
    -- CP-element group 580 join  transition  bypass 
    -- predecessors 575 
    -- marked predecessors 904 
    -- successors 584 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_update_start_
      -- 
    cpelement_group_580 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(575);
      marked_predecessors(0) <= cp_elements(904);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(580)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(580),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 581 transition  bypass 
    -- predecessors 585 
    -- successors 577 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_update_completed_
      -- 
    cp_elements(581) <= cp_elements(585);
    -- CP-element group 582 transition  output  bypass 
    -- predecessors 578 
    -- successors 583 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Sample/rr
      -- 
    cp_elements(582) <= cp_elements(578);
    rr_2595_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(582), ack => binary_585_inst_req_0); -- 
    -- CP-element group 583 transition  input  bypass 
    -- predecessors 582 
    -- successors 579 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Sample/ra
      -- 
    ra_2596_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_585_inst_ack_0, ack => cp_elements(583)); -- 
    -- CP-element group 584 transition  output  bypass 
    -- predecessors 580 
    -- successors 585 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Update/cr
      -- 
    cp_elements(584) <= cp_elements(580);
    cr_2600_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(584), ack => binary_585_inst_req_1); -- 
    -- CP-element group 585 transition  input  bypass 
    -- predecessors 584 
    -- successors 581 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_585_Update/ca
      -- 
    ca_2601_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_585_inst_ack_1, ack => cp_elements(585)); -- 
    -- CP-element group 586 join  fork  transition  bypass 
    -- predecessors 598 
    -- marked predecessors 622 
    -- successors 599 
    -- marked successors 588 589 472 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_active_
      -- 
    cpelement_group_586 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(598);
      marked_predecessors(0) <= cp_elements(622);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(586)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(586),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 587 transition  bypass 
    -- predecessors 601 
    -- successors 618 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_590_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_590_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_590_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_596_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_596_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_596_completed_
      -- 
    cp_elements(587) <= cp_elements(601);
    -- CP-element group 588 join  transition  bypass 
    -- predecessors 596 
    -- marked predecessors 586 
    -- successors 597 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_word_address_calculated
      -- 
    cpelement_group_588 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(596);
      marked_predecessors(0) <= cp_elements(586);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(588)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(588),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 589 join  transition  bypass 
    -- predecessors 594 
    -- marked predecessors 586 
    -- successors 595 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_root_address_calculated
      -- 
    cpelement_group_589 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(594);
      marked_predecessors(0) <= cp_elements(586);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(589)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(589),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 590 transition  bypass 
    -- predecessors 592 
    -- successors 593 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_address_resized
      -- 
    cp_elements(590) <= cp_elements(592);
    -- CP-element group 591 transition  output  bypass 
    -- predecessors 473 
    -- successors 592 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_addr_resize/base_resize_req
      -- 
    cp_elements(591) <= cp_elements(473);
    base_resize_req_2618_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(591), ack => ptr_deref_589_base_resize_req_0); -- 
    -- CP-element group 592 transition  input  bypass 
    -- predecessors 591 
    -- successors 590 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2619_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_base_resize_ack_0, ack => cp_elements(592)); -- 
    -- CP-element group 593 transition  output  bypass 
    -- predecessors 590 
    -- successors 594 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_plus_offset/sum_rename_req
      -- 
    cp_elements(593) <= cp_elements(590);
    sum_rename_req_2623_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(593), ack => ptr_deref_589_root_address_inst_req_0); -- 
    -- CP-element group 594 transition  input  bypass 
    -- predecessors 593 
    -- successors 589 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2624_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_root_address_inst_ack_0, ack => cp_elements(594)); -- 
    -- CP-element group 595 transition  output  bypass 
    -- predecessors 589 
    -- successors 596 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_word_addrgen/root_register_req
      -- 
    cp_elements(595) <= cp_elements(589);
    root_register_req_2628_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(595), ack => ptr_deref_589_addr_0_req_0); -- 
    -- CP-element group 596 transition  input  bypass 
    -- predecessors 595 
    -- successors 588 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_word_addrgen/root_register_ack
      -- 
    root_register_ack_2629_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_addr_0_ack_0, ack => cp_elements(596)); -- 
    -- CP-element group 597 transition  output  bypass 
    -- predecessors 588 
    -- successors 598 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/word_access_0/rr
      -- 
    cp_elements(597) <= cp_elements(588);
    rr_2639_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(597), ack => ptr_deref_589_load_0_req_0); -- 
    -- CP-element group 598 transition  input  bypass 
    -- predecessors 597 
    -- successors 586 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_request/word_access/word_access_0/ra
      -- 
    ra_2640_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_load_0_ack_0, ack => cp_elements(598)); -- 
    -- CP-element group 599 transition  output  bypass 
    -- predecessors 586 
    -- successors 600 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/word_access_0/cr
      -- 
    cp_elements(599) <= cp_elements(586);
    cr_2650_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(599), ack => ptr_deref_589_load_0_req_1); -- 
    -- CP-element group 600 transition  input  output  bypass 
    -- predecessors 599 
    -- successors 601 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/merge_req
      -- 
    ca_2651_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_load_0_ack_1, ack => cp_elements(600)); -- 
    merge_req_2652_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(600), ack => ptr_deref_589_gather_scatter_req_0); -- 
    -- CP-element group 601 transition  input  bypass 
    -- predecessors 600 
    -- successors 587 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_589_complete/merge_ack
      -- 
    merge_ack_2653_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_589_gather_scatter_ack_0, ack => cp_elements(601)); -- 
    -- CP-element group 602 join  fork  transition  bypass 
    -- predecessors 614 
    -- marked predecessors 622 
    -- successors 615 
    -- marked successors 604 605 454 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_active_
      -- 
    cpelement_group_602 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(614);
      marked_predecessors(0) <= cp_elements(622);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(602)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(602),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 603 transition  bypass 
    -- predecessors 617 
    -- successors 618 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_594_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_594_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_594_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_597_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_597_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_597_completed_
      -- 
    cp_elements(603) <= cp_elements(617);
    -- CP-element group 604 join  transition  bypass 
    -- predecessors 612 
    -- marked predecessors 602 
    -- successors 613 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_word_address_calculated
      -- 
    cpelement_group_604 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(612);
      marked_predecessors(0) <= cp_elements(602);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(604)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(604),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 605 join  transition  bypass 
    -- predecessors 610 
    -- marked predecessors 602 
    -- successors 611 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_root_address_calculated
      -- 
    cpelement_group_605 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(610);
      marked_predecessors(0) <= cp_elements(602);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(605)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(605),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 606 transition  bypass 
    -- predecessors 608 
    -- successors 609 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_address_resized
      -- 
    cp_elements(606) <= cp_elements(608);
    -- CP-element group 607 transition  output  bypass 
    -- predecessors 455 
    -- successors 608 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_addr_resize/base_resize_req
      -- 
    cp_elements(607) <= cp_elements(455);
    base_resize_req_2670_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(607), ack => ptr_deref_593_base_resize_req_0); -- 
    -- CP-element group 608 transition  input  bypass 
    -- predecessors 607 
    -- successors 606 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2671_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_base_resize_ack_0, ack => cp_elements(608)); -- 
    -- CP-element group 609 transition  output  bypass 
    -- predecessors 606 
    -- successors 610 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_plus_offset/sum_rename_req
      -- 
    cp_elements(609) <= cp_elements(606);
    sum_rename_req_2675_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(609), ack => ptr_deref_593_root_address_inst_req_0); -- 
    -- CP-element group 610 transition  input  bypass 
    -- predecessors 609 
    -- successors 605 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2676_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_root_address_inst_ack_0, ack => cp_elements(610)); -- 
    -- CP-element group 611 transition  output  bypass 
    -- predecessors 605 
    -- successors 612 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_word_addrgen/root_register_req
      -- 
    cp_elements(611) <= cp_elements(605);
    root_register_req_2680_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(611), ack => ptr_deref_593_addr_0_req_0); -- 
    -- CP-element group 612 transition  input  bypass 
    -- predecessors 611 
    -- successors 604 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_word_addrgen/root_register_ack
      -- 
    root_register_ack_2681_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_addr_0_ack_0, ack => cp_elements(612)); -- 
    -- CP-element group 613 transition  output  bypass 
    -- predecessors 604 
    -- successors 614 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/word_access_0/rr
      -- 
    cp_elements(613) <= cp_elements(604);
    rr_2691_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(613), ack => ptr_deref_593_load_0_req_0); -- 
    -- CP-element group 614 transition  input  bypass 
    -- predecessors 613 
    -- successors 602 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_request/word_access/word_access_0/ra
      -- 
    ra_2692_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_load_0_ack_0, ack => cp_elements(614)); -- 
    -- CP-element group 615 transition  output  bypass 
    -- predecessors 602 
    -- successors 616 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/word_access_0/cr
      -- 
    cp_elements(615) <= cp_elements(602);
    cr_2702_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(615), ack => ptr_deref_593_load_0_req_1); -- 
    -- CP-element group 616 transition  input  output  bypass 
    -- predecessors 615 
    -- successors 617 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/merge_req
      -- 
    ca_2703_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_load_0_ack_1, ack => cp_elements(616)); -- 
    merge_req_2704_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(616), ack => ptr_deref_593_gather_scatter_req_0); -- 
    -- CP-element group 617 transition  input  bypass 
    -- predecessors 616 
    -- successors 603 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_593_complete/merge_ack
      -- 
    merge_ack_2705_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_593_gather_scatter_ack_0, ack => cp_elements(617)); -- 
    -- CP-element group 618 join  fork  transition  bypass 
    -- predecessors 587 603 
    -- successors 621 623 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_trigger_
      -- 
    cpelement_group_618 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(587);
      predecessors(1) <= cp_elements(603);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(618)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(618),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 619 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_active_
      -- 
    cp_elements(619) <= cp_elements(7);
    -- CP-element group 620 join  transition  bypass 
    -- predecessors 622 624 
    -- successors 934 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_599_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_599_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_599_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_714_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_714_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_714_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_715_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_715_trigger_
      -- 
    cpelement_group_620 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(622);
      predecessors(1) <= cp_elements(624);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(620)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(620),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 621 join  transition  bypass 
    -- predecessors 618 
    -- marked predecessors 622 
    -- successors 625 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_sample_start_
      -- 
    cpelement_group_621 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(618);
      marked_predecessors(0) <= cp_elements(622);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(621)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(621),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 622 fork  transition  bypass 
    -- predecessors 626 
    -- successors 620 
    -- marked successors 586 602 621 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_sample_completed_
      -- 
    cp_elements(622) <= cp_elements(626);
    -- CP-element group 623 join  transition  bypass 
    -- predecessors 618 
    -- marked predecessors 936 
    -- successors 627 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_update_start_
      -- 
    cpelement_group_623 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(618);
      marked_predecessors(0) <= cp_elements(936);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(623)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(623),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 624 transition  bypass 
    -- predecessors 628 
    -- successors 620 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_update_completed_
      -- 
    cp_elements(624) <= cp_elements(628);
    -- CP-element group 625 transition  output  bypass 
    -- predecessors 621 
    -- successors 626 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Sample/rr
      -- 
    cp_elements(625) <= cp_elements(621);
    rr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(625), ack => binary_598_inst_req_0); -- 
    -- CP-element group 626 transition  input  bypass 
    -- predecessors 625 
    -- successors 622 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Sample/ra
      -- 
    ra_2726_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_598_inst_ack_0, ack => cp_elements(626)); -- 
    -- CP-element group 627 transition  output  bypass 
    -- predecessors 623 
    -- successors 628 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Update/cr
      -- 
    cp_elements(627) <= cp_elements(623);
    cr_2730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(627), ack => binary_598_inst_req_1); -- 
    -- CP-element group 628 transition  input  bypass 
    -- predecessors 627 
    -- successors 624 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_598_Update/ca
      -- 
    ca_2731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_598_inst_ack_1, ack => cp_elements(628)); -- 
    -- CP-element group 629 join  fork  transition  bypass 
    -- predecessors 641 
    -- marked predecessors 665 
    -- successors 642 
    -- marked successors 631 632 407 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_active_
      -- 
    cpelement_group_629 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(641);
      marked_predecessors(0) <= cp_elements(665);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(629)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(629),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 630 transition  bypass 
    -- predecessors 644 
    -- successors 661 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_603_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_603_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_603_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_609_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_609_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_609_completed_
      -- 
    cp_elements(630) <= cp_elements(644);
    -- CP-element group 631 join  transition  bypass 
    -- predecessors 639 
    -- marked predecessors 629 
    -- successors 640 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_word_address_calculated
      -- 
    cpelement_group_631 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(639);
      marked_predecessors(0) <= cp_elements(629);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(631)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(631),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 632 join  transition  bypass 
    -- predecessors 637 
    -- marked predecessors 629 
    -- successors 638 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_root_address_calculated
      -- 
    cpelement_group_632 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(637);
      marked_predecessors(0) <= cp_elements(629);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(632)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(632),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 633 transition  bypass 
    -- predecessors 635 
    -- successors 636 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_address_resized
      -- 
    cp_elements(633) <= cp_elements(635);
    -- CP-element group 634 transition  output  bypass 
    -- predecessors 408 
    -- successors 635 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_addr_resize/base_resize_req
      -- 
    cp_elements(634) <= cp_elements(408);
    base_resize_req_2748_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(634), ack => ptr_deref_602_base_resize_req_0); -- 
    -- CP-element group 635 transition  input  bypass 
    -- predecessors 634 
    -- successors 633 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2749_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_base_resize_ack_0, ack => cp_elements(635)); -- 
    -- CP-element group 636 transition  output  bypass 
    -- predecessors 633 
    -- successors 637 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_plus_offset/sum_rename_req
      -- 
    cp_elements(636) <= cp_elements(633);
    sum_rename_req_2753_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(636), ack => ptr_deref_602_root_address_inst_req_0); -- 
    -- CP-element group 637 transition  input  bypass 
    -- predecessors 636 
    -- successors 632 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2754_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_root_address_inst_ack_0, ack => cp_elements(637)); -- 
    -- CP-element group 638 transition  output  bypass 
    -- predecessors 632 
    -- successors 639 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_word_addrgen/root_register_req
      -- 
    cp_elements(638) <= cp_elements(632);
    root_register_req_2758_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(638), ack => ptr_deref_602_addr_0_req_0); -- 
    -- CP-element group 639 transition  input  bypass 
    -- predecessors 638 
    -- successors 631 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_word_addrgen/root_register_ack
      -- 
    root_register_ack_2759_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_addr_0_ack_0, ack => cp_elements(639)); -- 
    -- CP-element group 640 transition  output  bypass 
    -- predecessors 631 
    -- successors 641 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/word_access_0/rr
      -- 
    cp_elements(640) <= cp_elements(631);
    rr_2769_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(640), ack => ptr_deref_602_load_0_req_0); -- 
    -- CP-element group 641 transition  input  bypass 
    -- predecessors 640 
    -- successors 629 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_request/word_access/word_access_0/ra
      -- 
    ra_2770_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_load_0_ack_0, ack => cp_elements(641)); -- 
    -- CP-element group 642 transition  output  bypass 
    -- predecessors 629 
    -- successors 643 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/word_access_0/cr
      -- 
    cp_elements(642) <= cp_elements(629);
    cr_2780_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(642), ack => ptr_deref_602_load_0_req_1); -- 
    -- CP-element group 643 transition  input  output  bypass 
    -- predecessors 642 
    -- successors 644 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/merge_req
      -- 
    ca_2781_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_load_0_ack_1, ack => cp_elements(643)); -- 
    merge_req_2782_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(643), ack => ptr_deref_602_gather_scatter_req_0); -- 
    -- CP-element group 644 transition  input  bypass 
    -- predecessors 643 
    -- successors 630 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_602_complete/merge_ack
      -- 
    merge_ack_2783_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_602_gather_scatter_ack_0, ack => cp_elements(644)); -- 
    -- CP-element group 645 join  fork  transition  bypass 
    -- predecessors 657 
    -- marked predecessors 665 
    -- successors 658 
    -- marked successors 389 647 648 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_active_
      -- 
    cpelement_group_645 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(657);
      marked_predecessors(0) <= cp_elements(665);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(645)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(645),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 646 transition  bypass 
    -- predecessors 660 
    -- successors 661 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_607_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_607_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_607_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_610_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_610_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_610_completed_
      -- 
    cp_elements(646) <= cp_elements(660);
    -- CP-element group 647 join  transition  bypass 
    -- predecessors 655 
    -- marked predecessors 645 
    -- successors 656 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_word_address_calculated
      -- 
    cpelement_group_647 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(655);
      marked_predecessors(0) <= cp_elements(645);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(647)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(647),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 648 join  transition  bypass 
    -- predecessors 653 
    -- marked predecessors 645 
    -- successors 654 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_root_address_calculated
      -- 
    cpelement_group_648 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(653);
      marked_predecessors(0) <= cp_elements(645);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(648)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(648),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 649 transition  bypass 
    -- predecessors 651 
    -- successors 652 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_address_resized
      -- 
    cp_elements(649) <= cp_elements(651);
    -- CP-element group 650 transition  output  bypass 
    -- predecessors 390 
    -- successors 651 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_addr_resize/base_resize_req
      -- 
    cp_elements(650) <= cp_elements(390);
    base_resize_req_2800_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(650), ack => ptr_deref_606_base_resize_req_0); -- 
    -- CP-element group 651 transition  input  bypass 
    -- predecessors 650 
    -- successors 649 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2801_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_base_resize_ack_0, ack => cp_elements(651)); -- 
    -- CP-element group 652 transition  output  bypass 
    -- predecessors 649 
    -- successors 653 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_plus_offset/sum_rename_req
      -- 
    cp_elements(652) <= cp_elements(649);
    sum_rename_req_2805_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(652), ack => ptr_deref_606_root_address_inst_req_0); -- 
    -- CP-element group 653 transition  input  bypass 
    -- predecessors 652 
    -- successors 648 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2806_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_root_address_inst_ack_0, ack => cp_elements(653)); -- 
    -- CP-element group 654 transition  output  bypass 
    -- predecessors 648 
    -- successors 655 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_word_addrgen/root_register_req
      -- 
    cp_elements(654) <= cp_elements(648);
    root_register_req_2810_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(654), ack => ptr_deref_606_addr_0_req_0); -- 
    -- CP-element group 655 transition  input  bypass 
    -- predecessors 654 
    -- successors 647 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_word_addrgen/root_register_ack
      -- 
    root_register_ack_2811_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_addr_0_ack_0, ack => cp_elements(655)); -- 
    -- CP-element group 656 transition  output  bypass 
    -- predecessors 647 
    -- successors 657 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/word_access_0/rr
      -- 
    cp_elements(656) <= cp_elements(647);
    rr_2821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(656), ack => ptr_deref_606_load_0_req_0); -- 
    -- CP-element group 657 transition  input  bypass 
    -- predecessors 656 
    -- successors 645 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_request/word_access/word_access_0/ra
      -- 
    ra_2822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_load_0_ack_0, ack => cp_elements(657)); -- 
    -- CP-element group 658 transition  output  bypass 
    -- predecessors 645 
    -- successors 659 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/word_access_0/cr
      -- 
    cp_elements(658) <= cp_elements(645);
    cr_2832_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(658), ack => ptr_deref_606_load_0_req_1); -- 
    -- CP-element group 659 transition  input  output  bypass 
    -- predecessors 658 
    -- successors 660 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/merge_req
      -- 
    ca_2833_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_load_0_ack_1, ack => cp_elements(659)); -- 
    merge_req_2834_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(659), ack => ptr_deref_606_gather_scatter_req_0); -- 
    -- CP-element group 660 transition  input  bypass 
    -- predecessors 659 
    -- successors 646 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_606_complete/merge_ack
      -- 
    merge_ack_2835_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_606_gather_scatter_ack_0, ack => cp_elements(660)); -- 
    -- CP-element group 661 join  fork  transition  bypass 
    -- predecessors 630 646 
    -- successors 664 666 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_trigger_
      -- 
    cpelement_group_661 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(630);
      predecessors(1) <= cp_elements(646);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(661)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(661),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 662 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_active_
      -- 
    cp_elements(662) <= cp_elements(7);
    -- CP-element group 663 join  transition  bypass 
    -- predecessors 665 667 
    -- successors 966 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_733_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_733_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_733_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_734_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_734_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_612_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_612_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_612_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_completed_
      -- 
    cpelement_group_663 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(665);
      predecessors(1) <= cp_elements(667);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(663)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(663),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 664 join  transition  bypass 
    -- predecessors 661 
    -- marked predecessors 665 
    -- successors 668 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_sample_start_
      -- 
    cpelement_group_664 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(661);
      marked_predecessors(0) <= cp_elements(665);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(664)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(664),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 665 fork  transition  bypass 
    -- predecessors 669 
    -- successors 663 
    -- marked successors 629 645 664 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_sample_completed_
      -- 
    cp_elements(665) <= cp_elements(669);
    -- CP-element group 666 join  transition  bypass 
    -- predecessors 661 
    -- marked predecessors 968 
    -- successors 670 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_update_start_
      -- 
    cpelement_group_666 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(661);
      marked_predecessors(0) <= cp_elements(968);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(666)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(666),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 667 transition  bypass 
    -- predecessors 671 
    -- successors 663 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_update_completed_
      -- 
    cp_elements(667) <= cp_elements(671);
    -- CP-element group 668 transition  output  bypass 
    -- predecessors 664 
    -- successors 669 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Sample/rr
      -- 
    cp_elements(668) <= cp_elements(664);
    rr_2855_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(668), ack => binary_611_inst_req_0); -- 
    -- CP-element group 669 transition  input  bypass 
    -- predecessors 668 
    -- successors 665 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Sample/ra
      -- 
    ra_2856_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_611_inst_ack_0, ack => cp_elements(669)); -- 
    -- CP-element group 670 transition  output  bypass 
    -- predecessors 666 
    -- successors 671 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Update/cr
      -- 
    cp_elements(670) <= cp_elements(666);
    cr_2860_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(670), ack => binary_611_inst_req_1); -- 
    -- CP-element group 671 transition  input  bypass 
    -- predecessors 670 
    -- successors 667 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_611_Update/ca
      -- 
    ca_2861_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_611_inst_ack_1, ack => cp_elements(671)); -- 
    -- CP-element group 672 join  fork  transition  bypass 
    -- predecessors 684 
    -- marked predecessors 708 
    -- successors 685 
    -- marked successors 342 674 675 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_active_
      -- 
    cpelement_group_672 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(684);
      marked_predecessors(0) <= cp_elements(708);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(672)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(672),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 673 transition  bypass 
    -- predecessors 687 
    -- successors 704 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_616_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_616_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_616_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_622_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_622_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_622_completed_
      -- 
    cp_elements(673) <= cp_elements(687);
    -- CP-element group 674 join  transition  bypass 
    -- predecessors 682 
    -- marked predecessors 672 
    -- successors 683 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_word_address_calculated
      -- 
    cpelement_group_674 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(682);
      marked_predecessors(0) <= cp_elements(672);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(674)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(674),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 675 join  transition  bypass 
    -- predecessors 680 
    -- marked predecessors 672 
    -- successors 681 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_root_address_calculated
      -- 
    cpelement_group_675 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(680);
      marked_predecessors(0) <= cp_elements(672);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(675)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(675),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 676 transition  bypass 
    -- predecessors 678 
    -- successors 679 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_address_resized
      -- 
    cp_elements(676) <= cp_elements(678);
    -- CP-element group 677 transition  output  bypass 
    -- predecessors 343 
    -- successors 678 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_addr_resize/base_resize_req
      -- 
    cp_elements(677) <= cp_elements(343);
    base_resize_req_2878_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(677), ack => ptr_deref_615_base_resize_req_0); -- 
    -- CP-element group 678 transition  input  bypass 
    -- predecessors 677 
    -- successors 676 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2879_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_base_resize_ack_0, ack => cp_elements(678)); -- 
    -- CP-element group 679 transition  output  bypass 
    -- predecessors 676 
    -- successors 680 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_plus_offset/sum_rename_req
      -- 
    cp_elements(679) <= cp_elements(676);
    sum_rename_req_2883_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(679), ack => ptr_deref_615_root_address_inst_req_0); -- 
    -- CP-element group 680 transition  input  bypass 
    -- predecessors 679 
    -- successors 675 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2884_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_root_address_inst_ack_0, ack => cp_elements(680)); -- 
    -- CP-element group 681 transition  output  bypass 
    -- predecessors 675 
    -- successors 682 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_word_addrgen/root_register_req
      -- 
    cp_elements(681) <= cp_elements(675);
    root_register_req_2888_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(681), ack => ptr_deref_615_addr_0_req_0); -- 
    -- CP-element group 682 transition  input  bypass 
    -- predecessors 681 
    -- successors 674 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_word_addrgen/root_register_ack
      -- 
    root_register_ack_2889_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_addr_0_ack_0, ack => cp_elements(682)); -- 
    -- CP-element group 683 transition  output  bypass 
    -- predecessors 674 
    -- successors 684 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/word_access_0/rr
      -- 
    cp_elements(683) <= cp_elements(674);
    rr_2899_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(683), ack => ptr_deref_615_load_0_req_0); -- 
    -- CP-element group 684 transition  input  bypass 
    -- predecessors 683 
    -- successors 672 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_request/word_access/word_access_0/ra
      -- 
    ra_2900_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_load_0_ack_0, ack => cp_elements(684)); -- 
    -- CP-element group 685 transition  output  bypass 
    -- predecessors 672 
    -- successors 686 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/word_access_0/cr
      -- 
    cp_elements(685) <= cp_elements(672);
    cr_2910_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(685), ack => ptr_deref_615_load_0_req_1); -- 
    -- CP-element group 686 transition  input  output  bypass 
    -- predecessors 685 
    -- successors 687 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/merge_req
      -- 
    ca_2911_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_load_0_ack_1, ack => cp_elements(686)); -- 
    merge_req_2912_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(686), ack => ptr_deref_615_gather_scatter_req_0); -- 
    -- CP-element group 687 transition  input  bypass 
    -- predecessors 686 
    -- successors 673 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_615_complete/merge_ack
      -- 
    merge_ack_2913_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_615_gather_scatter_ack_0, ack => cp_elements(687)); -- 
    -- CP-element group 688 join  fork  transition  bypass 
    -- predecessors 700 
    -- marked predecessors 708 
    -- successors 701 
    -- marked successors 690 691 324 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_active_
      -- 
    cpelement_group_688 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(700);
      marked_predecessors(0) <= cp_elements(708);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(688)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(688),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 689 transition  bypass 
    -- predecessors 703 
    -- successors 704 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_620_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_620_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_620_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_623_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_623_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_623_completed_
      -- 
    cp_elements(689) <= cp_elements(703);
    -- CP-element group 690 join  transition  bypass 
    -- predecessors 698 
    -- marked predecessors 688 
    -- successors 699 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_word_address_calculated
      -- 
    cpelement_group_690 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(698);
      marked_predecessors(0) <= cp_elements(688);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(690)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(690),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 691 join  transition  bypass 
    -- predecessors 696 
    -- marked predecessors 688 
    -- successors 697 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_root_address_calculated
      -- 
    cpelement_group_691 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(696);
      marked_predecessors(0) <= cp_elements(688);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(691)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(691),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 692 transition  bypass 
    -- predecessors 694 
    -- successors 695 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_address_resized
      -- 
    cp_elements(692) <= cp_elements(694);
    -- CP-element group 693 transition  output  bypass 
    -- predecessors 325 
    -- successors 694 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_addr_resize/base_resize_req
      -- 
    cp_elements(693) <= cp_elements(325);
    base_resize_req_2930_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(693), ack => ptr_deref_619_base_resize_req_0); -- 
    -- CP-element group 694 transition  input  bypass 
    -- predecessors 693 
    -- successors 692 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_2931_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_base_resize_ack_0, ack => cp_elements(694)); -- 
    -- CP-element group 695 transition  output  bypass 
    -- predecessors 692 
    -- successors 696 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_plus_offset/sum_rename_req
      -- 
    cp_elements(695) <= cp_elements(692);
    sum_rename_req_2935_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(695), ack => ptr_deref_619_root_address_inst_req_0); -- 
    -- CP-element group 696 transition  input  bypass 
    -- predecessors 695 
    -- successors 691 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_2936_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_root_address_inst_ack_0, ack => cp_elements(696)); -- 
    -- CP-element group 697 transition  output  bypass 
    -- predecessors 691 
    -- successors 698 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_word_addrgen/root_register_req
      -- 
    cp_elements(697) <= cp_elements(691);
    root_register_req_2940_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(697), ack => ptr_deref_619_addr_0_req_0); -- 
    -- CP-element group 698 transition  input  bypass 
    -- predecessors 697 
    -- successors 690 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_word_addrgen/root_register_ack
      -- 
    root_register_ack_2941_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_addr_0_ack_0, ack => cp_elements(698)); -- 
    -- CP-element group 699 transition  output  bypass 
    -- predecessors 690 
    -- successors 700 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/word_access_0/rr
      -- 
    cp_elements(699) <= cp_elements(690);
    rr_2951_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(699), ack => ptr_deref_619_load_0_req_0); -- 
    -- CP-element group 700 transition  input  bypass 
    -- predecessors 699 
    -- successors 688 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_request/word_access/word_access_0/ra
      -- 
    ra_2952_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_load_0_ack_0, ack => cp_elements(700)); -- 
    -- CP-element group 701 transition  output  bypass 
    -- predecessors 688 
    -- successors 702 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/word_access_0/cr
      -- 
    cp_elements(701) <= cp_elements(688);
    cr_2962_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(701), ack => ptr_deref_619_load_0_req_1); -- 
    -- CP-element group 702 transition  input  output  bypass 
    -- predecessors 701 
    -- successors 703 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/merge_req
      -- 
    ca_2963_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_load_0_ack_1, ack => cp_elements(702)); -- 
    merge_req_2964_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(702), ack => ptr_deref_619_gather_scatter_req_0); -- 
    -- CP-element group 703 transition  input  bypass 
    -- predecessors 702 
    -- successors 689 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_619_complete/merge_ack
      -- 
    merge_ack_2965_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_619_gather_scatter_ack_0, ack => cp_elements(703)); -- 
    -- CP-element group 704 join  fork  transition  bypass 
    -- predecessors 689 673 
    -- successors 707 709 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_trigger_
      -- 
    cpelement_group_704 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(689);
      predecessors(1) <= cp_elements(673);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(704)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(704),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 705 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_active_
      -- 
    cp_elements(705) <= cp_elements(7);
    -- CP-element group 706 join  transition  bypass 
    -- predecessors 708 710 
    -- successors 998 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_752_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_752_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_752_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_753_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_753_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_625_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_625_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_625_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_completed_
      -- 
    cpelement_group_706 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(708);
      predecessors(1) <= cp_elements(710);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(706)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(706),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 707 join  transition  bypass 
    -- predecessors 704 
    -- marked predecessors 708 
    -- successors 711 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_sample_start_
      -- 
    cpelement_group_707 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(704);
      marked_predecessors(0) <= cp_elements(708);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(707)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(707),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 708 fork  transition  bypass 
    -- predecessors 712 
    -- successors 706 
    -- marked successors 688 707 672 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_sample_completed_
      -- 
    cp_elements(708) <= cp_elements(712);
    -- CP-element group 709 join  transition  bypass 
    -- predecessors 704 
    -- marked predecessors 1000 
    -- successors 713 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_update_start_
      -- 
    cpelement_group_709 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(704);
      marked_predecessors(0) <= cp_elements(1000);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(709)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(709),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 710 transition  bypass 
    -- predecessors 714 
    -- successors 706 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_update_completed_
      -- 
    cp_elements(710) <= cp_elements(714);
    -- CP-element group 711 transition  output  bypass 
    -- predecessors 707 
    -- successors 712 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Sample/rr
      -- 
    cp_elements(711) <= cp_elements(707);
    rr_2985_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(711), ack => binary_624_inst_req_0); -- 
    -- CP-element group 712 transition  input  bypass 
    -- predecessors 711 
    -- successors 708 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Sample/ra
      -- 
    ra_2986_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_624_inst_ack_0, ack => cp_elements(712)); -- 
    -- CP-element group 713 transition  output  bypass 
    -- predecessors 709 
    -- successors 714 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Update/cr
      -- 
    cp_elements(713) <= cp_elements(709);
    cr_2990_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(713), ack => binary_624_inst_req_1); -- 
    -- CP-element group 714 transition  input  bypass 
    -- predecessors 713 
    -- successors 710 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_624_Update/ca
      -- 
    ca_2991_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_624_inst_ack_1, ack => cp_elements(714)); -- 
    -- CP-element group 715 join  fork  transition  bypass 
    -- predecessors 727 
    -- marked predecessors 751 
    -- successors 728 
    -- marked successors 717 718 277 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_active_
      -- 
    cpelement_group_715 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(727);
      marked_predecessors(0) <= cp_elements(751);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(715)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(715),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 716 transition  bypass 
    -- predecessors 730 
    -- successors 747 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_629_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_629_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_629_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_635_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_635_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_635_completed_
      -- 
    cp_elements(716) <= cp_elements(730);
    -- CP-element group 717 join  transition  bypass 
    -- predecessors 725 
    -- marked predecessors 715 
    -- successors 726 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_word_address_calculated
      -- 
    cpelement_group_717 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(725);
      marked_predecessors(0) <= cp_elements(715);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(717)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(717),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 718 join  transition  bypass 
    -- predecessors 723 
    -- marked predecessors 715 
    -- successors 724 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_root_address_calculated
      -- 
    cpelement_group_718 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(723);
      marked_predecessors(0) <= cp_elements(715);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(718)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(718),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 719 transition  bypass 
    -- predecessors 721 
    -- successors 722 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_address_resized
      -- 
    cp_elements(719) <= cp_elements(721);
    -- CP-element group 720 transition  output  bypass 
    -- predecessors 278 
    -- successors 721 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_addr_resize/base_resize_req
      -- 
    cp_elements(720) <= cp_elements(278);
    base_resize_req_3008_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(720), ack => ptr_deref_628_base_resize_req_0); -- 
    -- CP-element group 721 transition  input  bypass 
    -- predecessors 720 
    -- successors 719 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3009_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_base_resize_ack_0, ack => cp_elements(721)); -- 
    -- CP-element group 722 transition  output  bypass 
    -- predecessors 719 
    -- successors 723 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_plus_offset/sum_rename_req
      -- 
    cp_elements(722) <= cp_elements(719);
    sum_rename_req_3013_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(722), ack => ptr_deref_628_root_address_inst_req_0); -- 
    -- CP-element group 723 transition  input  bypass 
    -- predecessors 722 
    -- successors 718 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3014_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_root_address_inst_ack_0, ack => cp_elements(723)); -- 
    -- CP-element group 724 transition  output  bypass 
    -- predecessors 718 
    -- successors 725 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_word_addrgen/root_register_req
      -- 
    cp_elements(724) <= cp_elements(718);
    root_register_req_3018_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(724), ack => ptr_deref_628_addr_0_req_0); -- 
    -- CP-element group 725 transition  input  bypass 
    -- predecessors 724 
    -- successors 717 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_word_addrgen/root_register_ack
      -- 
    root_register_ack_3019_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_addr_0_ack_0, ack => cp_elements(725)); -- 
    -- CP-element group 726 transition  output  bypass 
    -- predecessors 717 
    -- successors 727 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/word_access_0/rr
      -- 
    cp_elements(726) <= cp_elements(717);
    rr_3029_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(726), ack => ptr_deref_628_load_0_req_0); -- 
    -- CP-element group 727 transition  input  bypass 
    -- predecessors 726 
    -- successors 715 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_request/word_access/word_access_0/ra
      -- 
    ra_3030_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_load_0_ack_0, ack => cp_elements(727)); -- 
    -- CP-element group 728 transition  output  bypass 
    -- predecessors 715 
    -- successors 729 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/word_access_0/cr
      -- 
    cp_elements(728) <= cp_elements(715);
    cr_3040_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(728), ack => ptr_deref_628_load_0_req_1); -- 
    -- CP-element group 729 transition  input  output  bypass 
    -- predecessors 728 
    -- successors 730 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/merge_req
      -- 
    ca_3041_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_load_0_ack_1, ack => cp_elements(729)); -- 
    merge_req_3042_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(729), ack => ptr_deref_628_gather_scatter_req_0); -- 
    -- CP-element group 730 transition  input  bypass 
    -- predecessors 729 
    -- successors 716 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_628_complete/merge_ack
      -- 
    merge_ack_3043_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_628_gather_scatter_ack_0, ack => cp_elements(730)); -- 
    -- CP-element group 731 join  fork  transition  bypass 
    -- predecessors 743 
    -- marked predecessors 751 
    -- successors 744 
    -- marked successors 733 734 259 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_active_
      -- 
    cpelement_group_731 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(743);
      marked_predecessors(0) <= cp_elements(751);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(731)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(731),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 732 transition  bypass 
    -- predecessors 746 
    -- successors 747 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_633_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_633_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_633_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_636_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_636_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_636_completed_
      -- 
    cp_elements(732) <= cp_elements(746);
    -- CP-element group 733 join  transition  bypass 
    -- predecessors 741 
    -- marked predecessors 731 
    -- successors 742 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_word_address_calculated
      -- 
    cpelement_group_733 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(741);
      marked_predecessors(0) <= cp_elements(731);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(733)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(733),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 734 join  transition  bypass 
    -- predecessors 739 
    -- marked predecessors 731 
    -- successors 740 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_root_address_calculated
      -- 
    cpelement_group_734 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(739);
      marked_predecessors(0) <= cp_elements(731);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(734)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(734),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 735 transition  bypass 
    -- predecessors 737 
    -- successors 738 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_address_resized
      -- 
    cp_elements(735) <= cp_elements(737);
    -- CP-element group 736 transition  output  bypass 
    -- predecessors 260 
    -- successors 737 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_addr_resize/base_resize_req
      -- 
    cp_elements(736) <= cp_elements(260);
    base_resize_req_3060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(736), ack => ptr_deref_632_base_resize_req_0); -- 
    -- CP-element group 737 transition  input  bypass 
    -- predecessors 736 
    -- successors 735 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_base_resize_ack_0, ack => cp_elements(737)); -- 
    -- CP-element group 738 transition  output  bypass 
    -- predecessors 735 
    -- successors 739 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_plus_offset/sum_rename_req
      -- 
    cp_elements(738) <= cp_elements(735);
    sum_rename_req_3065_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(738), ack => ptr_deref_632_root_address_inst_req_0); -- 
    -- CP-element group 739 transition  input  bypass 
    -- predecessors 738 
    -- successors 734 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3066_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_root_address_inst_ack_0, ack => cp_elements(739)); -- 
    -- CP-element group 740 transition  output  bypass 
    -- predecessors 734 
    -- successors 741 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_word_addrgen/root_register_req
      -- 
    cp_elements(740) <= cp_elements(734);
    root_register_req_3070_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(740), ack => ptr_deref_632_addr_0_req_0); -- 
    -- CP-element group 741 transition  input  bypass 
    -- predecessors 740 
    -- successors 733 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_word_addrgen/root_register_ack
      -- 
    root_register_ack_3071_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_addr_0_ack_0, ack => cp_elements(741)); -- 
    -- CP-element group 742 transition  output  bypass 
    -- predecessors 733 
    -- successors 743 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/word_access_0/rr
      -- 
    cp_elements(742) <= cp_elements(733);
    rr_3081_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(742), ack => ptr_deref_632_load_0_req_0); -- 
    -- CP-element group 743 transition  input  bypass 
    -- predecessors 742 
    -- successors 731 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_request/word_access/word_access_0/ra
      -- 
    ra_3082_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_load_0_ack_0, ack => cp_elements(743)); -- 
    -- CP-element group 744 transition  output  bypass 
    -- predecessors 731 
    -- successors 745 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/word_access_0/cr
      -- 
    cp_elements(744) <= cp_elements(731);
    cr_3092_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(744), ack => ptr_deref_632_load_0_req_1); -- 
    -- CP-element group 745 transition  input  output  bypass 
    -- predecessors 744 
    -- successors 746 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/merge_req
      -- 
    ca_3093_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_load_0_ack_1, ack => cp_elements(745)); -- 
    merge_req_3094_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(745), ack => ptr_deref_632_gather_scatter_req_0); -- 
    -- CP-element group 746 transition  input  bypass 
    -- predecessors 745 
    -- successors 732 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_632_complete/merge_ack
      -- 
    merge_ack_3095_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_632_gather_scatter_ack_0, ack => cp_elements(746)); -- 
    -- CP-element group 747 join  fork  transition  bypass 
    -- predecessors 716 732 
    -- successors 752 750 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_trigger_
      -- 
    cpelement_group_747 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(716);
      predecessors(1) <= cp_elements(732);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(747)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(747),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 748 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_active_
      -- 
    cp_elements(748) <= cp_elements(7);
    -- CP-element group 749 join  transition  bypass 
    -- predecessors 751 753 
    -- successors 1030 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_638_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_638_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_638_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_772_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_771_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_772_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_771_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_771_active_
      -- 
    cpelement_group_749 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(751);
      predecessors(1) <= cp_elements(753);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(749)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(749),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 750 join  transition  bypass 
    -- predecessors 747 
    -- marked predecessors 751 
    -- successors 754 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_sample_start_
      -- 
    cpelement_group_750 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(747);
      marked_predecessors(0) <= cp_elements(751);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(750)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(750),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 751 fork  transition  bypass 
    -- predecessors 755 
    -- successors 749 
    -- marked successors 715 731 750 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_sample_completed_
      -- 
    cp_elements(751) <= cp_elements(755);
    -- CP-element group 752 join  transition  bypass 
    -- predecessors 747 
    -- marked predecessors 1032 
    -- successors 756 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_update_start_
      -- 
    cpelement_group_752 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(747);
      marked_predecessors(0) <= cp_elements(1032);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(752)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(752),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 753 transition  bypass 
    -- predecessors 757 
    -- successors 749 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_update_completed_
      -- 
    cp_elements(753) <= cp_elements(757);
    -- CP-element group 754 transition  output  bypass 
    -- predecessors 750 
    -- successors 755 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Sample/rr
      -- 
    cp_elements(754) <= cp_elements(750);
    rr_3115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(754), ack => binary_637_inst_req_0); -- 
    -- CP-element group 755 transition  input  bypass 
    -- predecessors 754 
    -- successors 751 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Sample/ra
      -- 
    ra_3116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_637_inst_ack_0, ack => cp_elements(755)); -- 
    -- CP-element group 756 transition  output  bypass 
    -- predecessors 752 
    -- successors 757 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Update/cr
      -- 
    cp_elements(756) <= cp_elements(752);
    cr_3120_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(756), ack => binary_637_inst_req_1); -- 
    -- CP-element group 757 transition  input  bypass 
    -- predecessors 756 
    -- successors 753 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_637_Update/ca
      -- 
    ca_3121_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_637_inst_ack_1, ack => cp_elements(757)); -- 
    -- CP-element group 758 join  fork  transition  bypass 
    -- predecessors 770 
    -- marked predecessors 794 
    -- successors 771 
    -- marked successors 760 761 212 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_active_
      -- 
    cpelement_group_758 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(770);
      marked_predecessors(0) <= cp_elements(794);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(758)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(758),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 759 transition  bypass 
    -- predecessors 773 
    -- successors 790 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_642_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_642_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_642_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_648_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_648_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_648_completed_
      -- 
    cp_elements(759) <= cp_elements(773);
    -- CP-element group 760 join  transition  bypass 
    -- predecessors 768 
    -- marked predecessors 758 
    -- successors 769 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_word_address_calculated
      -- 
    cpelement_group_760 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(768);
      marked_predecessors(0) <= cp_elements(758);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(760)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(760),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 761 join  transition  bypass 
    -- predecessors 766 
    -- marked predecessors 758 
    -- successors 767 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_root_address_calculated
      -- 
    cpelement_group_761 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(766);
      marked_predecessors(0) <= cp_elements(758);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(761)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(761),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 762 transition  bypass 
    -- predecessors 764 
    -- successors 765 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_address_resized
      -- 
    cp_elements(762) <= cp_elements(764);
    -- CP-element group 763 transition  output  bypass 
    -- predecessors 213 
    -- successors 764 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_addr_resize/base_resize_req
      -- 
    cp_elements(763) <= cp_elements(213);
    base_resize_req_3138_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(763), ack => ptr_deref_641_base_resize_req_0); -- 
    -- CP-element group 764 transition  input  bypass 
    -- predecessors 763 
    -- successors 762 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3139_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_base_resize_ack_0, ack => cp_elements(764)); -- 
    -- CP-element group 765 transition  output  bypass 
    -- predecessors 762 
    -- successors 766 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_plus_offset/sum_rename_req
      -- 
    cp_elements(765) <= cp_elements(762);
    sum_rename_req_3143_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(765), ack => ptr_deref_641_root_address_inst_req_0); -- 
    -- CP-element group 766 transition  input  bypass 
    -- predecessors 765 
    -- successors 761 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3144_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_root_address_inst_ack_0, ack => cp_elements(766)); -- 
    -- CP-element group 767 transition  output  bypass 
    -- predecessors 761 
    -- successors 768 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_word_addrgen/root_register_req
      -- 
    cp_elements(767) <= cp_elements(761);
    root_register_req_3148_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(767), ack => ptr_deref_641_addr_0_req_0); -- 
    -- CP-element group 768 transition  input  bypass 
    -- predecessors 767 
    -- successors 760 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_word_addrgen/root_register_ack
      -- 
    root_register_ack_3149_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_addr_0_ack_0, ack => cp_elements(768)); -- 
    -- CP-element group 769 transition  output  bypass 
    -- predecessors 760 
    -- successors 770 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/word_access_0/rr
      -- 
    cp_elements(769) <= cp_elements(760);
    rr_3159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(769), ack => ptr_deref_641_load_0_req_0); -- 
    -- CP-element group 770 transition  input  bypass 
    -- predecessors 769 
    -- successors 758 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_request/word_access/word_access_0/ra
      -- 
    ra_3160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_load_0_ack_0, ack => cp_elements(770)); -- 
    -- CP-element group 771 transition  output  bypass 
    -- predecessors 758 
    -- successors 772 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/word_access_0/cr
      -- 
    cp_elements(771) <= cp_elements(758);
    cr_3170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(771), ack => ptr_deref_641_load_0_req_1); -- 
    -- CP-element group 772 transition  input  output  bypass 
    -- predecessors 771 
    -- successors 773 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/merge_req
      -- 
    ca_3171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_load_0_ack_1, ack => cp_elements(772)); -- 
    merge_req_3172_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(772), ack => ptr_deref_641_gather_scatter_req_0); -- 
    -- CP-element group 773 transition  input  bypass 
    -- predecessors 772 
    -- successors 759 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_641_complete/merge_ack
      -- 
    merge_ack_3173_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_641_gather_scatter_ack_0, ack => cp_elements(773)); -- 
    -- CP-element group 774 join  fork  transition  bypass 
    -- predecessors 786 
    -- marked predecessors 794 
    -- successors 787 
    -- marked successors 776 777 194 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_active_
      -- 
    cpelement_group_774 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(786);
      marked_predecessors(0) <= cp_elements(794);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(774)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(774),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 775 transition  bypass 
    -- predecessors 789 
    -- successors 790 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_646_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_646_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_646_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_649_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_649_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_649_completed_
      -- 
    cp_elements(775) <= cp_elements(789);
    -- CP-element group 776 join  transition  bypass 
    -- predecessors 784 
    -- marked predecessors 774 
    -- successors 785 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_word_address_calculated
      -- 
    cpelement_group_776 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(784);
      marked_predecessors(0) <= cp_elements(774);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(776)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(776),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 777 join  transition  bypass 
    -- predecessors 782 
    -- marked predecessors 774 
    -- successors 783 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_root_address_calculated
      -- 
    cpelement_group_777 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(782);
      marked_predecessors(0) <= cp_elements(774);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(777)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(777),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 778 transition  bypass 
    -- predecessors 780 
    -- successors 781 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_address_resized
      -- 
    cp_elements(778) <= cp_elements(780);
    -- CP-element group 779 transition  output  bypass 
    -- predecessors 195 
    -- successors 780 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_addr_resize/base_resize_req
      -- 
    cp_elements(779) <= cp_elements(195);
    base_resize_req_3190_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(779), ack => ptr_deref_645_base_resize_req_0); -- 
    -- CP-element group 780 transition  input  bypass 
    -- predecessors 779 
    -- successors 778 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3191_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_base_resize_ack_0, ack => cp_elements(780)); -- 
    -- CP-element group 781 transition  output  bypass 
    -- predecessors 778 
    -- successors 782 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_plus_offset/sum_rename_req
      -- 
    cp_elements(781) <= cp_elements(778);
    sum_rename_req_3195_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(781), ack => ptr_deref_645_root_address_inst_req_0); -- 
    -- CP-element group 782 transition  input  bypass 
    -- predecessors 781 
    -- successors 777 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3196_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_root_address_inst_ack_0, ack => cp_elements(782)); -- 
    -- CP-element group 783 transition  output  bypass 
    -- predecessors 777 
    -- successors 784 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_word_addrgen/root_register_req
      -- 
    cp_elements(783) <= cp_elements(777);
    root_register_req_3200_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(783), ack => ptr_deref_645_addr_0_req_0); -- 
    -- CP-element group 784 transition  input  bypass 
    -- predecessors 783 
    -- successors 776 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_word_addrgen/root_register_ack
      -- 
    root_register_ack_3201_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_addr_0_ack_0, ack => cp_elements(784)); -- 
    -- CP-element group 785 transition  output  bypass 
    -- predecessors 776 
    -- successors 786 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/word_access_0/rr
      -- 
    cp_elements(785) <= cp_elements(776);
    rr_3211_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(785), ack => ptr_deref_645_load_0_req_0); -- 
    -- CP-element group 786 transition  input  bypass 
    -- predecessors 785 
    -- successors 774 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_request/word_access/word_access_0/ra
      -- 
    ra_3212_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_load_0_ack_0, ack => cp_elements(786)); -- 
    -- CP-element group 787 transition  output  bypass 
    -- predecessors 774 
    -- successors 788 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/word_access_0/cr
      -- 
    cp_elements(787) <= cp_elements(774);
    cr_3222_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(787), ack => ptr_deref_645_load_0_req_1); -- 
    -- CP-element group 788 transition  input  output  bypass 
    -- predecessors 787 
    -- successors 789 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/merge_req
      -- 
    ca_3223_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_load_0_ack_1, ack => cp_elements(788)); -- 
    merge_req_3224_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(788), ack => ptr_deref_645_gather_scatter_req_0); -- 
    -- CP-element group 789 transition  input  bypass 
    -- predecessors 788 
    -- successors 775 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_645_complete/merge_ack
      -- 
    merge_ack_3225_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_645_gather_scatter_ack_0, ack => cp_elements(789)); -- 
    -- CP-element group 790 join  fork  transition  bypass 
    -- predecessors 759 775 
    -- successors 793 795 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_trigger_
      -- 
    cpelement_group_790 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(759);
      predecessors(1) <= cp_elements(775);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(790)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(790),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 791 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_active_
      -- 
    cp_elements(791) <= cp_elements(7);
    -- CP-element group 792 join  transition  bypass 
    -- predecessors 794 796 
    -- successors 1062 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_651_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_651_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_651_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_791_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_791_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_790_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_790_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_790_completed_
      -- 
    cpelement_group_792 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(794);
      predecessors(1) <= cp_elements(796);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(792)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(792),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 793 join  transition  bypass 
    -- predecessors 790 
    -- marked predecessors 794 
    -- successors 797 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_sample_start_
      -- 
    cpelement_group_793 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(790);
      marked_predecessors(0) <= cp_elements(794);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(793)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(793),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 794 fork  transition  bypass 
    -- predecessors 798 
    -- successors 792 
    -- marked successors 758 774 793 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_sample_completed_
      -- 
    cp_elements(794) <= cp_elements(798);
    -- CP-element group 795 join  transition  bypass 
    -- predecessors 790 
    -- marked predecessors 1064 
    -- successors 799 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_update_start_
      -- 
    cpelement_group_795 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(790);
      marked_predecessors(0) <= cp_elements(1064);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(795)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(795),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 796 transition  bypass 
    -- predecessors 800 
    -- successors 792 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_update_completed_
      -- 
    cp_elements(796) <= cp_elements(800);
    -- CP-element group 797 transition  output  bypass 
    -- predecessors 793 
    -- successors 798 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Sample/rr
      -- 
    cp_elements(797) <= cp_elements(793);
    rr_3245_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(797), ack => binary_650_inst_req_0); -- 
    -- CP-element group 798 transition  input  bypass 
    -- predecessors 797 
    -- successors 794 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Sample/ra
      -- 
    ra_3246_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_650_inst_ack_0, ack => cp_elements(798)); -- 
    -- CP-element group 799 transition  output  bypass 
    -- predecessors 795 
    -- successors 800 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Update/cr
      -- 
    cp_elements(799) <= cp_elements(795);
    cr_3250_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(799), ack => binary_650_inst_req_1); -- 
    -- CP-element group 800 transition  input  bypass 
    -- predecessors 799 
    -- successors 796 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_650_Update/ca
      -- 
    ca_3251_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_650_inst_ack_1, ack => cp_elements(800)); -- 
    -- CP-element group 801 join  fork  transition  bypass 
    -- predecessors 813 
    -- marked predecessors 837 
    -- successors 814 
    -- marked successors 147 803 804 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_active_
      -- 
    cpelement_group_801 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(813);
      marked_predecessors(0) <= cp_elements(837);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(801)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(801),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 802 transition  bypass 
    -- predecessors 816 
    -- successors 833 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_655_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_655_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_655_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_661_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_661_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_661_completed_
      -- 
    cp_elements(802) <= cp_elements(816);
    -- CP-element group 803 join  transition  bypass 
    -- predecessors 811 
    -- marked predecessors 801 
    -- successors 812 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_word_address_calculated
      -- 
    cpelement_group_803 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(811);
      marked_predecessors(0) <= cp_elements(801);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(803)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(803),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 804 join  transition  bypass 
    -- predecessors 809 
    -- marked predecessors 801 
    -- successors 810 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_root_address_calculated
      -- 
    cpelement_group_804 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(809);
      marked_predecessors(0) <= cp_elements(801);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(804)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(804),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 805 transition  bypass 
    -- predecessors 807 
    -- successors 808 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_address_resized
      -- 
    cp_elements(805) <= cp_elements(807);
    -- CP-element group 806 transition  output  bypass 
    -- predecessors 148 
    -- successors 807 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_addr_resize/base_resize_req
      -- 
    cp_elements(806) <= cp_elements(148);
    base_resize_req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(806), ack => ptr_deref_654_base_resize_req_0); -- 
    -- CP-element group 807 transition  input  bypass 
    -- predecessors 806 
    -- successors 805 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_base_resize_ack_0, ack => cp_elements(807)); -- 
    -- CP-element group 808 transition  output  bypass 
    -- predecessors 805 
    -- successors 809 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_plus_offset/sum_rename_req
      -- 
    cp_elements(808) <= cp_elements(805);
    sum_rename_req_3273_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(808), ack => ptr_deref_654_root_address_inst_req_0); -- 
    -- CP-element group 809 transition  input  bypass 
    -- predecessors 808 
    -- successors 804 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3274_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_root_address_inst_ack_0, ack => cp_elements(809)); -- 
    -- CP-element group 810 transition  output  bypass 
    -- predecessors 804 
    -- successors 811 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_word_addrgen/root_register_req
      -- 
    cp_elements(810) <= cp_elements(804);
    root_register_req_3278_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(810), ack => ptr_deref_654_addr_0_req_0); -- 
    -- CP-element group 811 transition  input  bypass 
    -- predecessors 810 
    -- successors 803 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_word_addrgen/root_register_ack
      -- 
    root_register_ack_3279_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_addr_0_ack_0, ack => cp_elements(811)); -- 
    -- CP-element group 812 transition  output  bypass 
    -- predecessors 803 
    -- successors 813 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/word_access_0/rr
      -- 
    cp_elements(812) <= cp_elements(803);
    rr_3289_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(812), ack => ptr_deref_654_load_0_req_0); -- 
    -- CP-element group 813 transition  input  bypass 
    -- predecessors 812 
    -- successors 801 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_request/word_access/word_access_0/ra
      -- 
    ra_3290_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_load_0_ack_0, ack => cp_elements(813)); -- 
    -- CP-element group 814 transition  output  bypass 
    -- predecessors 801 
    -- successors 815 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/word_access_0/cr
      -- 
    cp_elements(814) <= cp_elements(801);
    cr_3300_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(814), ack => ptr_deref_654_load_0_req_1); -- 
    -- CP-element group 815 transition  input  output  bypass 
    -- predecessors 814 
    -- successors 816 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/merge_req
      -- 
    ca_3301_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_load_0_ack_1, ack => cp_elements(815)); -- 
    merge_req_3302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(815), ack => ptr_deref_654_gather_scatter_req_0); -- 
    -- CP-element group 816 transition  input  bypass 
    -- predecessors 815 
    -- successors 802 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_654_complete/merge_ack
      -- 
    merge_ack_3303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_654_gather_scatter_ack_0, ack => cp_elements(816)); -- 
    -- CP-element group 817 join  fork  transition  bypass 
    -- predecessors 829 
    -- marked predecessors 837 
    -- successors 830 
    -- marked successors 129 819 820 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_active_
      -- 
    cpelement_group_817 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(829);
      marked_predecessors(0) <= cp_elements(837);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(817)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(817),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 818 transition  bypass 
    -- predecessors 832 
    -- successors 833 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_659_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_659_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_659_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_662_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_662_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_662_completed_
      -- 
    cp_elements(818) <= cp_elements(832);
    -- CP-element group 819 join  transition  bypass 
    -- predecessors 827 
    -- marked predecessors 817 
    -- successors 828 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_word_address_calculated
      -- 
    cpelement_group_819 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(827);
      marked_predecessors(0) <= cp_elements(817);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(819)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(819),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 820 join  transition  bypass 
    -- predecessors 825 
    -- marked predecessors 817 
    -- successors 826 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_root_address_calculated
      -- 
    cpelement_group_820 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(825);
      marked_predecessors(0) <= cp_elements(817);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(820)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(820),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 821 transition  bypass 
    -- predecessors 823 
    -- successors 824 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_address_resized
      -- 
    cp_elements(821) <= cp_elements(823);
    -- CP-element group 822 transition  output  bypass 
    -- predecessors 130 
    -- successors 823 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_addr_resize/base_resize_req
      -- 
    cp_elements(822) <= cp_elements(130);
    base_resize_req_3320_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(822), ack => ptr_deref_658_base_resize_req_0); -- 
    -- CP-element group 823 transition  input  bypass 
    -- predecessors 822 
    -- successors 821 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3321_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_base_resize_ack_0, ack => cp_elements(823)); -- 
    -- CP-element group 824 transition  output  bypass 
    -- predecessors 821 
    -- successors 825 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_plus_offset/sum_rename_req
      -- 
    cp_elements(824) <= cp_elements(821);
    sum_rename_req_3325_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(824), ack => ptr_deref_658_root_address_inst_req_0); -- 
    -- CP-element group 825 transition  input  bypass 
    -- predecessors 824 
    -- successors 820 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3326_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_root_address_inst_ack_0, ack => cp_elements(825)); -- 
    -- CP-element group 826 transition  output  bypass 
    -- predecessors 820 
    -- successors 827 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_word_addrgen/root_register_req
      -- 
    cp_elements(826) <= cp_elements(820);
    root_register_req_3330_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(826), ack => ptr_deref_658_addr_0_req_0); -- 
    -- CP-element group 827 transition  input  bypass 
    -- predecessors 826 
    -- successors 819 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_word_addrgen/root_register_ack
      -- 
    root_register_ack_3331_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_addr_0_ack_0, ack => cp_elements(827)); -- 
    -- CP-element group 828 transition  output  bypass 
    -- predecessors 819 
    -- successors 829 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/word_access_0/rr
      -- 
    cp_elements(828) <= cp_elements(819);
    rr_3341_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(828), ack => ptr_deref_658_load_0_req_0); -- 
    -- CP-element group 829 transition  input  bypass 
    -- predecessors 828 
    -- successors 817 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_request/word_access/word_access_0/ra
      -- 
    ra_3342_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_load_0_ack_0, ack => cp_elements(829)); -- 
    -- CP-element group 830 transition  output  bypass 
    -- predecessors 817 
    -- successors 831 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/word_access_0/cr
      -- 
    cp_elements(830) <= cp_elements(817);
    cr_3352_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(830), ack => ptr_deref_658_load_0_req_1); -- 
    -- CP-element group 831 transition  input  output  bypass 
    -- predecessors 830 
    -- successors 832 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/merge_req
      -- 
    ca_3353_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_load_0_ack_1, ack => cp_elements(831)); -- 
    merge_req_3354_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(831), ack => ptr_deref_658_gather_scatter_req_0); -- 
    -- CP-element group 832 transition  input  bypass 
    -- predecessors 831 
    -- successors 818 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_658_complete/merge_ack
      -- 
    merge_ack_3355_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_658_gather_scatter_ack_0, ack => cp_elements(832)); -- 
    -- CP-element group 833 join  fork  transition  bypass 
    -- predecessors 802 818 
    -- successors 836 838 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_trigger_
      -- 
    cpelement_group_833 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(802);
      predecessors(1) <= cp_elements(818);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(833)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(833),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 834 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_active_
      -- 
    cp_elements(834) <= cp_elements(7);
    -- CP-element group 835 join  transition  bypass 
    -- predecessors 837 839 
    -- successors 1094 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_664_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_664_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_664_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_810_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_810_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_809_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_809_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_809_completed_
      -- 
    cpelement_group_835 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(837);
      predecessors(1) <= cp_elements(839);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(835)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(835),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 836 join  transition  bypass 
    -- predecessors 833 
    -- marked predecessors 837 
    -- successors 840 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_sample_start_
      -- 
    cpelement_group_836 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(833);
      marked_predecessors(0) <= cp_elements(837);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(836)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(836),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 837 fork  transition  bypass 
    -- predecessors 841 
    -- successors 835 
    -- marked successors 801 817 836 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_sample_completed_
      -- 
    cp_elements(837) <= cp_elements(841);
    -- CP-element group 838 join  transition  bypass 
    -- predecessors 833 
    -- marked predecessors 1096 
    -- successors 842 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_update_start_
      -- 
    cpelement_group_838 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(833);
      marked_predecessors(0) <= cp_elements(1096);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(838)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(838),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 839 transition  bypass 
    -- predecessors 843 
    -- successors 835 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_update_completed_
      -- 
    cp_elements(839) <= cp_elements(843);
    -- CP-element group 840 transition  output  bypass 
    -- predecessors 836 
    -- successors 841 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Sample/rr
      -- 
    cp_elements(840) <= cp_elements(836);
    rr_3375_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(840), ack => binary_663_inst_req_0); -- 
    -- CP-element group 841 transition  input  bypass 
    -- predecessors 840 
    -- successors 837 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Sample/ra
      -- 
    ra_3376_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_663_inst_ack_0, ack => cp_elements(841)); -- 
    -- CP-element group 842 transition  output  bypass 
    -- predecessors 838 
    -- successors 843 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Update/cr
      -- 
    cp_elements(842) <= cp_elements(838);
    cr_3380_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(842), ack => binary_663_inst_req_1); -- 
    -- CP-element group 843 transition  input  bypass 
    -- predecessors 842 
    -- successors 839 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_663_Update/ca
      -- 
    ca_3381_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_663_inst_ack_1, ack => cp_elements(843)); -- 
    -- CP-element group 844 join  fork  transition  bypass 
    -- predecessors 856 
    -- marked predecessors 880 
    -- successors 857 
    -- marked successors 82 846 847 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_active_
      -- 
    cpelement_group_844 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(856);
      marked_predecessors(0) <= cp_elements(880);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(844)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(844),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 845 transition  bypass 
    -- predecessors 859 
    -- successors 876 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_674_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_674_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_674_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_668_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_668_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_668_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_completed_
      -- 
    cp_elements(845) <= cp_elements(859);
    -- CP-element group 846 join  transition  bypass 
    -- predecessors 854 
    -- marked predecessors 844 
    -- successors 855 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_word_address_calculated
      -- 
    cpelement_group_846 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(854);
      marked_predecessors(0) <= cp_elements(844);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(846)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(846),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 847 join  transition  bypass 
    -- predecessors 852 
    -- marked predecessors 844 
    -- successors 853 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_root_address_calculated
      -- 
    cpelement_group_847 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(852);
      marked_predecessors(0) <= cp_elements(844);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(847)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(847),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 848 transition  bypass 
    -- predecessors 850 
    -- successors 851 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_address_resized
      -- 
    cp_elements(848) <= cp_elements(850);
    -- CP-element group 849 transition  output  bypass 
    -- predecessors 83 
    -- successors 850 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_addr_resize/base_resize_req
      -- 
    cp_elements(849) <= cp_elements(83);
    base_resize_req_3398_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(849), ack => ptr_deref_667_base_resize_req_0); -- 
    -- CP-element group 850 transition  input  bypass 
    -- predecessors 849 
    -- successors 848 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3399_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_base_resize_ack_0, ack => cp_elements(850)); -- 
    -- CP-element group 851 transition  output  bypass 
    -- predecessors 848 
    -- successors 852 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_plus_offset/sum_rename_req
      -- 
    cp_elements(851) <= cp_elements(848);
    sum_rename_req_3403_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(851), ack => ptr_deref_667_root_address_inst_req_0); -- 
    -- CP-element group 852 transition  input  bypass 
    -- predecessors 851 
    -- successors 847 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3404_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_root_address_inst_ack_0, ack => cp_elements(852)); -- 
    -- CP-element group 853 transition  output  bypass 
    -- predecessors 847 
    -- successors 854 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_word_addrgen/root_register_req
      -- 
    cp_elements(853) <= cp_elements(847);
    root_register_req_3408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(853), ack => ptr_deref_667_addr_0_req_0); -- 
    -- CP-element group 854 transition  input  bypass 
    -- predecessors 853 
    -- successors 846 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_word_addrgen/root_register_ack
      -- 
    root_register_ack_3409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_addr_0_ack_0, ack => cp_elements(854)); -- 
    -- CP-element group 855 transition  output  bypass 
    -- predecessors 846 
    -- successors 856 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/word_access_0/rr
      -- 
    cp_elements(855) <= cp_elements(846);
    rr_3419_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(855), ack => ptr_deref_667_load_0_req_0); -- 
    -- CP-element group 856 transition  input  bypass 
    -- predecessors 855 
    -- successors 844 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_request/word_access/word_access_0/ra
      -- 
    ra_3420_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_load_0_ack_0, ack => cp_elements(856)); -- 
    -- CP-element group 857 transition  output  bypass 
    -- predecessors 844 
    -- successors 858 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/word_access_0/cr
      -- 
    cp_elements(857) <= cp_elements(844);
    cr_3430_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(857), ack => ptr_deref_667_load_0_req_1); -- 
    -- CP-element group 858 transition  input  output  bypass 
    -- predecessors 857 
    -- successors 859 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/merge_req
      -- 
    ca_3431_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_load_0_ack_1, ack => cp_elements(858)); -- 
    merge_req_3432_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(858), ack => ptr_deref_667_gather_scatter_req_0); -- 
    -- CP-element group 859 transition  input  bypass 
    -- predecessors 858 
    -- successors 845 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_667_complete/merge_ack
      -- 
    merge_ack_3433_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_667_gather_scatter_ack_0, ack => cp_elements(859)); -- 
    -- CP-element group 860 join  fork  transition  bypass 
    -- predecessors 872 
    -- marked predecessors 880 
    -- successors 873 
    -- marked successors 64 862 863 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_active_
      -- 
    cpelement_group_860 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(872);
      marked_predecessors(0) <= cp_elements(880);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(860)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(860),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 861 transition  bypass 
    -- predecessors 875 
    -- successors 876 
    -- members (7) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_672_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_672_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_672_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_675_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_675_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_675_completed_
      -- 
    cp_elements(861) <= cp_elements(875);
    -- CP-element group 862 join  transition  bypass 
    -- predecessors 870 
    -- marked predecessors 860 
    -- successors 871 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_word_address_calculated
      -- 
    cpelement_group_862 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(870);
      marked_predecessors(0) <= cp_elements(860);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(862)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(862),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 863 join  transition  bypass 
    -- predecessors 868 
    -- marked predecessors 860 
    -- successors 869 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_root_address_calculated
      -- 
    cpelement_group_863 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(868);
      marked_predecessors(0) <= cp_elements(860);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(863)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(863),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 864 transition  bypass 
    -- predecessors 866 
    -- successors 867 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_address_resized
      -- 
    cp_elements(864) <= cp_elements(866);
    -- CP-element group 865 transition  output  bypass 
    -- predecessors 65 
    -- successors 866 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_addr_resize/base_resize_req
      -- 
    cp_elements(865) <= cp_elements(65);
    base_resize_req_3450_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(865), ack => ptr_deref_671_base_resize_req_0); -- 
    -- CP-element group 866 transition  input  bypass 
    -- predecessors 865 
    -- successors 864 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3451_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_base_resize_ack_0, ack => cp_elements(866)); -- 
    -- CP-element group 867 transition  output  bypass 
    -- predecessors 864 
    -- successors 868 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_plus_offset/sum_rename_req
      -- 
    cp_elements(867) <= cp_elements(864);
    sum_rename_req_3455_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(867), ack => ptr_deref_671_root_address_inst_req_0); -- 
    -- CP-element group 868 transition  input  bypass 
    -- predecessors 867 
    -- successors 863 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3456_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_root_address_inst_ack_0, ack => cp_elements(868)); -- 
    -- CP-element group 869 transition  output  bypass 
    -- predecessors 863 
    -- successors 870 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_word_addrgen/root_register_req
      -- 
    cp_elements(869) <= cp_elements(863);
    root_register_req_3460_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(869), ack => ptr_deref_671_addr_0_req_0); -- 
    -- CP-element group 870 transition  input  bypass 
    -- predecessors 869 
    -- successors 862 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_word_addrgen/root_register_ack
      -- 
    root_register_ack_3461_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_addr_0_ack_0, ack => cp_elements(870)); -- 
    -- CP-element group 871 transition  output  bypass 
    -- predecessors 862 
    -- successors 872 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/word_access_0/rr
      -- 
    cp_elements(871) <= cp_elements(862);
    rr_3471_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(871), ack => ptr_deref_671_load_0_req_0); -- 
    -- CP-element group 872 transition  input  bypass 
    -- predecessors 871 
    -- successors 860 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_request/word_access/word_access_0/ra
      -- 
    ra_3472_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_load_0_ack_0, ack => cp_elements(872)); -- 
    -- CP-element group 873 transition  output  bypass 
    -- predecessors 860 
    -- successors 874 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/word_access_0/cr
      -- 
    cp_elements(873) <= cp_elements(860);
    cr_3482_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(873), ack => ptr_deref_671_load_0_req_1); -- 
    -- CP-element group 874 transition  input  output  bypass 
    -- predecessors 873 
    -- successors 875 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/merge_req
      -- 
    ca_3483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_load_0_ack_1, ack => cp_elements(874)); -- 
    merge_req_3484_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(874), ack => ptr_deref_671_gather_scatter_req_0); -- 
    -- CP-element group 875 transition  input  bypass 
    -- predecessors 874 
    -- successors 861 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_671_complete/merge_ack
      -- 
    merge_ack_3485_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_671_gather_scatter_ack_0, ack => cp_elements(875)); -- 
    -- CP-element group 876 join  fork  transition  bypass 
    -- predecessors 845 861 
    -- successors 879 881 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_trigger_
      -- 
    cpelement_group_876 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(845);
      predecessors(1) <= cp_elements(861);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(876)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(876),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 877 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_active_
      -- 
    cp_elements(877) <= cp_elements(7);
    -- CP-element group 878 join  transition  bypass 
    -- predecessors 880 882 
    -- successors 1126 
    -- members (9) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_677_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_677_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_677_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_829_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_829_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_828_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_828_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_828_completed_
      -- 
    cpelement_group_878 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(880);
      predecessors(1) <= cp_elements(882);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(878)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(878),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 879 join  transition  bypass 
    -- predecessors 876 
    -- marked predecessors 880 
    -- successors 883 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_sample_start_
      -- 
    cpelement_group_879 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(876);
      marked_predecessors(0) <= cp_elements(880);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(879)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(879),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 880 fork  transition  bypass 
    -- predecessors 884 
    -- successors 878 
    -- marked successors 879 844 860 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_sample_completed_
      -- 
    cp_elements(880) <= cp_elements(884);
    -- CP-element group 881 join  transition  bypass 
    -- predecessors 876 
    -- marked predecessors 1128 
    -- successors 885 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_update_start_
      -- 
    cpelement_group_881 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(876);
      marked_predecessors(0) <= cp_elements(1128);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(881)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(881),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 882 transition  bypass 
    -- predecessors 886 
    -- successors 878 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_update_completed_
      -- 
    cp_elements(882) <= cp_elements(886);
    -- CP-element group 883 transition  output  bypass 
    -- predecessors 879 
    -- successors 884 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Sample/rr
      -- 
    cp_elements(883) <= cp_elements(879);
    rr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(883), ack => binary_676_inst_req_0); -- 
    -- CP-element group 884 transition  input  bypass 
    -- predecessors 883 
    -- successors 880 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Sample/ra
      -- 
    ra_3506_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_676_inst_ack_0, ack => cp_elements(884)); -- 
    -- CP-element group 885 transition  output  bypass 
    -- predecessors 881 
    -- successors 886 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Update/cr
      -- 
    cp_elements(885) <= cp_elements(881);
    cr_3510_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(885), ack => binary_676_inst_req_1); -- 
    -- CP-element group 886 transition  input  bypass 
    -- predecessors 885 
    -- successors 882 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_676_Update/ca
      -- 
    ca_3511_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_676_inst_ack_1, ack => cp_elements(886)); -- 
    -- CP-element group 887 join  fork  transition  bypass 
    -- predecessors 889 
    -- marked predecessors 893 
    -- successors 891 
    -- marked successors 490 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_682_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_682_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_682_completed_
      -- 
    cpelement_group_887 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(889);
      marked_predecessors(0) <= cp_elements(893);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(887)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(887),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 888 transition  output  bypass 
    -- predecessors 491 
    -- successors 889 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_register/req
      -- 
    cp_elements(888) <= cp_elements(491);
    req_3521_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(888), ack => simple_obj_ref_678_inst_req_0); -- 
    -- CP-element group 889 transition  input  bypass 
    -- predecessors 888 
    -- successors 887 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_680_register/ack
      -- 
    ack_3522_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_678_inst_ack_0, ack => cp_elements(889)); -- 
    -- CP-element group 890 join  fork  transition  bypass 
    -- predecessors 892 
    -- marked predecessors 896 
    -- successors 894 
    -- marked successors 491 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_685_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_685_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_685_completed_
      -- 
    cpelement_group_890 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(892);
      marked_predecessors(0) <= cp_elements(896);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(890)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(890),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 891 transition  output  bypass 
    -- predecessors 887 
    -- successors 892 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_register/req
      -- 
    cp_elements(891) <= cp_elements(887);
    req_3532_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(891), ack => simple_obj_ref_681_inst_req_0); -- 
    -- CP-element group 892 transition  input  bypass 
    -- predecessors 891 
    -- successors 890 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_683_register/ack
      -- 
    ack_3533_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_681_inst_ack_0, ack => cp_elements(892)); -- 
    -- CP-element group 893 join  fork  transition  bypass 
    -- predecessors 895 
    -- marked predecessors 899 
    -- successors 897 
    -- marked successors 887 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_688_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_688_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_688_completed_
      -- 
    cpelement_group_893 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(895);
      marked_predecessors(0) <= cp_elements(899);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(893)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(893),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 894 transition  output  bypass 
    -- predecessors 890 
    -- successors 895 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_register/req
      -- 
    cp_elements(894) <= cp_elements(890);
    req_3543_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(894), ack => simple_obj_ref_684_inst_req_0); -- 
    -- CP-element group 895 transition  input  bypass 
    -- predecessors 894 
    -- successors 893 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_686_register/ack
      -- 
    ack_3544_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_684_inst_ack_0, ack => cp_elements(895)); -- 
    -- CP-element group 896 join  fork  transition  bypass 
    -- predecessors 898 
    -- marked predecessors 903 
    -- successors 900 
    -- marked successors 890 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_691_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_691_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_691_completed_
      -- 
    cpelement_group_896 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(898);
      marked_predecessors(0) <= cp_elements(903);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(896)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(896),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 897 transition  output  bypass 
    -- predecessors 893 
    -- successors 898 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_register/req
      -- 
    cp_elements(897) <= cp_elements(893);
    req_3554_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(897), ack => simple_obj_ref_687_inst_req_0); -- 
    -- CP-element group 898 transition  input  bypass 
    -- predecessors 897 
    -- successors 896 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_689_register/ack
      -- 
    ack_3555_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_687_inst_ack_0, ack => cp_elements(898)); -- 
    -- CP-element group 899 fork  transition  bypass 
    -- predecessors 901 
    -- successors 908 
    -- marked successors 893 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_693_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_693_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_693_completed_
      -- 
    cp_elements(899) <= cp_elements(901);
    -- CP-element group 900 transition  output  bypass 
    -- predecessors 896 
    -- successors 901 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_register/req
      -- 
    cp_elements(900) <= cp_elements(896);
    req_3565_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(900), ack => simple_obj_ref_690_inst_req_0); -- 
    -- CP-element group 901 transition  input  bypass 
    -- predecessors 900 
    -- successors 899 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_692_register/ack
      -- 
    ack_3566_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_690_inst_ack_0, ack => cp_elements(901)); -- 
    -- CP-element group 902 join  transition  bypass 
    -- predecessors 905 577 
    -- marked predecessors 1174 
    -- successors 914 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_trigger_
      -- 
    cpelement_group_902 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(905);
      predecessors(1) <= cp_elements(577);
      marked_predecessors(0) <= cp_elements(1174);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(902)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(902),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 903 join  fork  transition  bypass 
    -- predecessors 916 
    -- marked predecessors 904 
    -- successors 917 934 
    -- marked successors 896 906 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_active_
      -- 
    cpelement_group_903 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(916);
      marked_predecessors(0) <= cp_elements(904);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(903)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(903),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 904 fork  transition  bypass 
    -- predecessors 918 
    -- successors 1175 
    -- marked successors 903 580 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_696_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_completed_
      -- 
    cp_elements(904) <= cp_elements(918);
    -- CP-element group 905 transition  bypass 
    -- predecessors 913 
    -- successors 902 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_word_address_calculated
      -- 
    cp_elements(905) <= cp_elements(913);
    -- CP-element group 906 join  transition  bypass 
    -- predecessors 911 
    -- marked predecessors 903 
    -- successors 912 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_root_address_calculated
      -- 
    cpelement_group_906 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(911);
      marked_predecessors(0) <= cp_elements(903);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(906)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(906),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 907 transition  bypass 
    -- predecessors 909 
    -- successors 910 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_address_resized
      -- 
    cp_elements(907) <= cp_elements(909);
    -- CP-element group 908 transition  output  bypass 
    -- predecessors 899 
    -- successors 909 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_addr_resize/base_resize_req
      -- 
    cp_elements(908) <= cp_elements(899);
    base_resize_req_3586_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(908), ack => ptr_deref_694_base_resize_req_0); -- 
    -- CP-element group 909 transition  input  bypass 
    -- predecessors 908 
    -- successors 907 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3587_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_base_resize_ack_0, ack => cp_elements(909)); -- 
    -- CP-element group 910 transition  output  bypass 
    -- predecessors 907 
    -- successors 911 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_plus_offset/sum_rename_req
      -- 
    cp_elements(910) <= cp_elements(907);
    sum_rename_req_3591_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(910), ack => ptr_deref_694_root_address_inst_req_0); -- 
    -- CP-element group 911 transition  input  bypass 
    -- predecessors 910 
    -- successors 906 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3592_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_root_address_inst_ack_0, ack => cp_elements(911)); -- 
    -- CP-element group 912 transition  output  bypass 
    -- predecessors 906 
    -- successors 913 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_word_addrgen/root_register_req
      -- 
    cp_elements(912) <= cp_elements(906);
    root_register_req_3596_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(912), ack => ptr_deref_694_addr_0_req_0); -- 
    -- CP-element group 913 transition  input  bypass 
    -- predecessors 912 
    -- successors 905 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_word_addrgen/root_register_ack
      -- 
    root_register_ack_3597_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_addr_0_ack_0, ack => cp_elements(913)); -- 
    -- CP-element group 914 transition  output  bypass 
    -- predecessors 902 
    -- successors 915 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/split_req
      -- 
    cp_elements(914) <= cp_elements(902);
    split_req_3601_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(914), ack => ptr_deref_694_gather_scatter_req_0); -- 
    -- CP-element group 915 transition  input  output  bypass 
    -- predecessors 914 
    -- successors 916 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/word_access_0/rr
      -- 
    split_ack_3602_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_gather_scatter_ack_0, ack => cp_elements(915)); -- 
    rr_3609_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(915), ack => ptr_deref_694_store_0_req_0); -- 
    -- CP-element group 916 transition  input  bypass 
    -- predecessors 915 
    -- successors 903 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_request/word_access/word_access_0/ra
      -- 
    ra_3610_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_store_0_ack_0, ack => cp_elements(916)); -- 
    -- CP-element group 917 transition  output  bypass 
    -- predecessors 903 
    -- successors 918 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/word_access_0/cr
      -- 
    cp_elements(917) <= cp_elements(903);
    cr_3620_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(917), ack => ptr_deref_694_store_0_req_1); -- 
    -- CP-element group 918 transition  input  bypass 
    -- predecessors 917 
    -- successors 904 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_694_complete/word_access/word_access_0/ca
      -- 
    ca_3621_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_694_store_0_ack_1, ack => cp_elements(918)); -- 
    -- CP-element group 919 join  fork  transition  bypass 
    -- predecessors 921 
    -- marked predecessors 925 
    -- successors 923 
    -- marked successors 436 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_701_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_701_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_701_completed_
      -- 
    cpelement_group_919 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(921);
      marked_predecessors(0) <= cp_elements(925);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(919)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(919),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 920 transition  output  bypass 
    -- predecessors 437 
    -- successors 921 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_register/req
      -- 
    cp_elements(920) <= cp_elements(437);
    req_3631_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(920), ack => simple_obj_ref_697_inst_req_0); -- 
    -- CP-element group 921 transition  input  bypass 
    -- predecessors 920 
    -- successors 919 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_699_register/ack
      -- 
    ack_3632_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_697_inst_ack_0, ack => cp_elements(921)); -- 
    -- CP-element group 922 join  fork  transition  bypass 
    -- predecessors 924 
    -- marked predecessors 928 
    -- successors 926 
    -- marked successors 437 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_704_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_704_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_704_completed_
      -- 
    cpelement_group_922 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(924);
      marked_predecessors(0) <= cp_elements(928);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(922)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(922),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 923 transition  output  bypass 
    -- predecessors 919 
    -- successors 924 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_register/req
      -- 
    cp_elements(923) <= cp_elements(919);
    req_3642_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(923), ack => simple_obj_ref_700_inst_req_0); -- 
    -- CP-element group 924 transition  input  bypass 
    -- predecessors 923 
    -- successors 922 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_702_register/ack
      -- 
    ack_3643_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_700_inst_ack_0, ack => cp_elements(924)); -- 
    -- CP-element group 925 join  fork  transition  bypass 
    -- predecessors 927 
    -- marked predecessors 931 
    -- successors 929 
    -- marked successors 919 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_707_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_707_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_707_completed_
      -- 
    cpelement_group_925 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(927);
      marked_predecessors(0) <= cp_elements(931);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(925)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(925),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 926 transition  output  bypass 
    -- predecessors 922 
    -- successors 927 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_register/req
      -- 
    cp_elements(926) <= cp_elements(922);
    req_3653_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(926), ack => simple_obj_ref_703_inst_req_0); -- 
    -- CP-element group 927 transition  input  bypass 
    -- predecessors 926 
    -- successors 925 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_705_register/ack
      -- 
    ack_3654_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_703_inst_ack_0, ack => cp_elements(927)); -- 
    -- CP-element group 928 join  fork  transition  bypass 
    -- predecessors 930 
    -- marked predecessors 935 
    -- successors 932 
    -- marked successors 922 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_710_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_710_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_710_completed_
      -- 
    cpelement_group_928 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(930);
      marked_predecessors(0) <= cp_elements(935);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(928)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(928),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 929 transition  output  bypass 
    -- predecessors 925 
    -- successors 930 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_register/req
      -- 
    cp_elements(929) <= cp_elements(925);
    req_3664_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(929), ack => simple_obj_ref_706_inst_req_0); -- 
    -- CP-element group 930 transition  input  bypass 
    -- predecessors 929 
    -- successors 928 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_708_register/ack
      -- 
    ack_3665_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_706_inst_ack_0, ack => cp_elements(930)); -- 
    -- CP-element group 931 fork  transition  bypass 
    -- predecessors 933 
    -- successors 940 
    -- marked successors 925 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_712_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_712_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_712_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_completed_
      -- 
    cp_elements(931) <= cp_elements(933);
    -- CP-element group 932 transition  output  bypass 
    -- predecessors 928 
    -- successors 933 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_register/req
      -- 
    cp_elements(932) <= cp_elements(928);
    req_3675_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(932), ack => simple_obj_ref_709_inst_req_0); -- 
    -- CP-element group 933 transition  input  bypass 
    -- predecessors 932 
    -- successors 931 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_711_register/ack
      -- 
    ack_3676_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_709_inst_ack_0, ack => cp_elements(933)); -- 
    -- CP-element group 934 join  transition  bypass 
    -- predecessors 903 937 620 
    -- marked predecessors 935 
    -- successors 946 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_trigger_
      -- 
    cpelement_group_934 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(903);
      predecessors(1) <= cp_elements(937);
      predecessors(2) <= cp_elements(620);
      marked_predecessors(0) <= cp_elements(935);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(934)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(934),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 935 join  fork  transition  bypass 
    -- predecessors 948 
    -- marked predecessors 936 
    -- successors 949 966 
    -- marked successors 928 934 938 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_active_
      -- 
    cpelement_group_935 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(948);
      marked_predecessors(0) <= cp_elements(936);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(935)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(935),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 936 fork  transition  bypass 
    -- predecessors 950 
    -- successors 1175 
    -- marked successors 935 623 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_715_completed_
      -- 
    cp_elements(936) <= cp_elements(950);
    -- CP-element group 937 transition  bypass 
    -- predecessors 945 
    -- successors 934 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_word_address_calculated
      -- 
    cp_elements(937) <= cp_elements(945);
    -- CP-element group 938 join  transition  bypass 
    -- predecessors 943 
    -- marked predecessors 935 
    -- successors 944 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_root_address_calculated
      -- 
    cpelement_group_938 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(943);
      marked_predecessors(0) <= cp_elements(935);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(938)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(938),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 939 transition  bypass 
    -- predecessors 941 
    -- successors 942 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_address_resized
      -- 
    cp_elements(939) <= cp_elements(941);
    -- CP-element group 940 transition  output  bypass 
    -- predecessors 931 
    -- successors 941 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_addr_resize/$entry
      -- 
    cp_elements(940) <= cp_elements(931);
    base_resize_req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(940), ack => ptr_deref_713_base_resize_req_0); -- 
    -- CP-element group 941 transition  input  bypass 
    -- predecessors 940 
    -- successors 939 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_addr_resize/$exit
      -- 
    base_resize_ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_base_resize_ack_0, ack => cp_elements(941)); -- 
    -- CP-element group 942 transition  output  bypass 
    -- predecessors 939 
    -- successors 943 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_plus_offset/$entry
      -- 
    cp_elements(942) <= cp_elements(939);
    sum_rename_req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(942), ack => ptr_deref_713_root_address_inst_req_0); -- 
    -- CP-element group 943 transition  input  bypass 
    -- predecessors 942 
    -- successors 938 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_base_plus_offset/$exit
      -- 
    sum_rename_ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_root_address_inst_ack_0, ack => cp_elements(943)); -- 
    -- CP-element group 944 transition  output  bypass 
    -- predecessors 938 
    -- successors 945 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_word_addrgen/root_register_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_word_addrgen/$entry
      -- 
    cp_elements(944) <= cp_elements(938);
    root_register_req_3706_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(944), ack => ptr_deref_713_addr_0_req_0); -- 
    -- CP-element group 945 transition  input  bypass 
    -- predecessors 944 
    -- successors 937 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_word_addrgen/root_register_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_word_addrgen/$exit
      -- 
    root_register_ack_3707_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_addr_0_ack_0, ack => cp_elements(945)); -- 
    -- CP-element group 946 transition  output  bypass 
    -- predecessors 934 
    -- successors 947 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/split_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/$entry
      -- 
    cp_elements(946) <= cp_elements(934);
    split_req_3711_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(946), ack => ptr_deref_713_gather_scatter_req_0); -- 
    -- CP-element group 947 transition  input  output  bypass 
    -- predecessors 946 
    -- successors 948 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/split_ack
      -- 
    split_ack_3712_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_gather_scatter_ack_0, ack => cp_elements(947)); -- 
    rr_3719_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(947), ack => ptr_deref_713_store_0_req_0); -- 
    -- CP-element group 948 transition  input  bypass 
    -- predecessors 947 
    -- successors 935 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_request/$exit
      -- 
    ra_3720_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_store_0_ack_0, ack => cp_elements(948)); -- 
    -- CP-element group 949 transition  output  bypass 
    -- predecessors 935 
    -- successors 950 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/word_access_0/cr
      -- 
    cp_elements(949) <= cp_elements(935);
    cr_3730_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(949), ack => ptr_deref_713_store_0_req_1); -- 
    -- CP-element group 950 transition  input  bypass 
    -- predecessors 949 
    -- successors 936 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_713_complete/word_access/word_access_0/ca
      -- 
    ca_3731_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_713_store_0_ack_1, ack => cp_elements(950)); -- 
    -- CP-element group 951 join  fork  transition  bypass 
    -- predecessors 953 
    -- marked predecessors 957 
    -- successors 955 
    -- marked successors 371 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_720_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_720_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_720_completed_
      -- 
    cpelement_group_951 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(953);
      marked_predecessors(0) <= cp_elements(957);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(951)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(951),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 952 transition  output  bypass 
    -- predecessors 372 
    -- successors 953 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_register/req
      -- 
    cp_elements(952) <= cp_elements(372);
    req_3741_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(952), ack => simple_obj_ref_716_inst_req_0); -- 
    -- CP-element group 953 transition  input  bypass 
    -- predecessors 952 
    -- successors 951 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_718_register/ack
      -- 
    ack_3742_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_716_inst_ack_0, ack => cp_elements(953)); -- 
    -- CP-element group 954 join  fork  transition  bypass 
    -- predecessors 956 
    -- marked predecessors 960 
    -- successors 958 
    -- marked successors 372 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_723_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_723_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_723_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_completed_
      -- 
    cpelement_group_954 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(956);
      marked_predecessors(0) <= cp_elements(960);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(954)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(954),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 955 transition  output  bypass 
    -- predecessors 951 
    -- successors 956 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_register/$entry
      -- 
    cp_elements(955) <= cp_elements(951);
    req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(955), ack => simple_obj_ref_719_inst_req_0); -- 
    -- CP-element group 956 transition  input  bypass 
    -- predecessors 955 
    -- successors 954 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_721_register/$exit
      -- 
    ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_719_inst_ack_0, ack => cp_elements(956)); -- 
    -- CP-element group 957 join  fork  transition  bypass 
    -- predecessors 959 
    -- marked predecessors 963 
    -- successors 961 
    -- marked successors 951 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_726_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_726_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_726_trigger_
      -- 
    cpelement_group_957 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(959);
      marked_predecessors(0) <= cp_elements(963);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(957)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(957),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 958 transition  output  bypass 
    -- predecessors 954 
    -- successors 959 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_register/$entry
      -- 
    cp_elements(958) <= cp_elements(954);
    req_3763_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(958), ack => simple_obj_ref_722_inst_req_0); -- 
    -- CP-element group 959 transition  input  bypass 
    -- predecessors 958 
    -- successors 957 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_724_register/$exit
      -- 
    ack_3764_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_722_inst_ack_0, ack => cp_elements(959)); -- 
    -- CP-element group 960 join  fork  transition  bypass 
    -- predecessors 962 
    -- marked predecessors 967 
    -- successors 964 
    -- marked successors 954 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_729_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_729_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_729_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_active_
      -- 
    cpelement_group_960 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(962);
      marked_predecessors(0) <= cp_elements(967);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(960)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(960),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 961 transition  output  bypass 
    -- predecessors 957 
    -- successors 962 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_register/$entry
      -- 
    cp_elements(961) <= cp_elements(957);
    req_3774_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(961), ack => simple_obj_ref_725_inst_req_0); -- 
    -- CP-element group 962 transition  input  bypass 
    -- predecessors 961 
    -- successors 960 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_727_register/$exit
      -- 
    ack_3775_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_725_inst_ack_0, ack => cp_elements(962)); -- 
    -- CP-element group 963 fork  transition  bypass 
    -- predecessors 965 
    -- successors 972 
    -- marked successors 957 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_731_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_731_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_731_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_active_
      -- 
    cp_elements(963) <= cp_elements(965);
    -- CP-element group 964 transition  output  bypass 
    -- predecessors 960 
    -- successors 965 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_register/req
      -- 
    cp_elements(964) <= cp_elements(960);
    req_3785_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(964), ack => simple_obj_ref_728_inst_req_0); -- 
    -- CP-element group 965 transition  input  bypass 
    -- predecessors 964 
    -- successors 963 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_730_register/ack
      -- 
    ack_3786_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_728_inst_ack_0, ack => cp_elements(965)); -- 
    -- CP-element group 966 join  transition  bypass 
    -- predecessors 935 969 663 
    -- marked predecessors 967 
    -- successors 978 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_trigger_
      -- 
    cpelement_group_966 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(935);
      predecessors(1) <= cp_elements(969);
      predecessors(2) <= cp_elements(663);
      marked_predecessors(0) <= cp_elements(967);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(966)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(966),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 967 join  fork  transition  bypass 
    -- predecessors 980 
    -- marked predecessors 968 
    -- successors 981 998 
    -- marked successors 960 966 970 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_active_
      -- 
    cpelement_group_967 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(980);
      marked_predecessors(0) <= cp_elements(968);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(967)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(967),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 968 fork  transition  bypass 
    -- predecessors 982 
    -- successors 1175 
    -- marked successors 967 666 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_734_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_completed_
      -- 
    cp_elements(968) <= cp_elements(982);
    -- CP-element group 969 transition  bypass 
    -- predecessors 977 
    -- successors 966 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_word_address_calculated
      -- 
    cp_elements(969) <= cp_elements(977);
    -- CP-element group 970 join  transition  bypass 
    -- predecessors 975 
    -- marked predecessors 967 
    -- successors 976 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_root_address_calculated
      -- 
    cpelement_group_970 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(975);
      marked_predecessors(0) <= cp_elements(967);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(970)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(970),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 971 transition  bypass 
    -- predecessors 973 
    -- successors 974 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_address_resized
      -- 
    cp_elements(971) <= cp_elements(973);
    -- CP-element group 972 transition  output  bypass 
    -- predecessors 963 
    -- successors 973 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_addr_resize/base_resize_req
      -- 
    cp_elements(972) <= cp_elements(963);
    base_resize_req_3806_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(972), ack => ptr_deref_732_base_resize_req_0); -- 
    -- CP-element group 973 transition  input  bypass 
    -- predecessors 972 
    -- successors 971 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_3807_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_base_resize_ack_0, ack => cp_elements(973)); -- 
    -- CP-element group 974 transition  output  bypass 
    -- predecessors 971 
    -- successors 975 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_plus_offset/$entry
      -- 
    cp_elements(974) <= cp_elements(971);
    sum_rename_req_3811_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(974), ack => ptr_deref_732_root_address_inst_req_0); -- 
    -- CP-element group 975 transition  input  bypass 
    -- predecessors 974 
    -- successors 970 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_plus_offset/sum_rename_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_base_plus_offset/$exit
      -- 
    sum_rename_ack_3812_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_root_address_inst_ack_0, ack => cp_elements(975)); -- 
    -- CP-element group 976 transition  output  bypass 
    -- predecessors 970 
    -- successors 977 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_word_addrgen/root_register_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_word_addrgen/$entry
      -- 
    cp_elements(976) <= cp_elements(970);
    root_register_req_3816_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(976), ack => ptr_deref_732_addr_0_req_0); -- 
    -- CP-element group 977 transition  input  bypass 
    -- predecessors 976 
    -- successors 969 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_word_addrgen/root_register_ack
      -- 
    root_register_ack_3817_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_addr_0_ack_0, ack => cp_elements(977)); -- 
    -- CP-element group 978 transition  output  bypass 
    -- predecessors 966 
    -- successors 979 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/split_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/$entry
      -- 
    cp_elements(978) <= cp_elements(966);
    split_req_3821_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(978), ack => ptr_deref_732_gather_scatter_req_0); -- 
    -- CP-element group 979 transition  input  output  bypass 
    -- predecessors 978 
    -- successors 980 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/$entry
      -- 
    split_ack_3822_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_gather_scatter_ack_0, ack => cp_elements(979)); -- 
    rr_3829_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(979), ack => ptr_deref_732_store_0_req_0); -- 
    -- CP-element group 980 transition  input  bypass 
    -- predecessors 979 
    -- successors 967 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_request/word_access/$exit
      -- 
    ra_3830_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_store_0_ack_0, ack => cp_elements(980)); -- 
    -- CP-element group 981 transition  output  bypass 
    -- predecessors 967 
    -- successors 982 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/word_access_0/cr
      -- 
    cp_elements(981) <= cp_elements(967);
    cr_3840_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(981), ack => ptr_deref_732_store_0_req_1); -- 
    -- CP-element group 982 transition  input  bypass 
    -- predecessors 981 
    -- successors 968 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_732_complete/word_access/word_access_0/ca
      -- 
    ca_3841_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_732_store_0_ack_1, ack => cp_elements(982)); -- 
    -- CP-element group 983 join  fork  transition  bypass 
    -- predecessors 985 
    -- marked predecessors 989 
    -- successors 987 
    -- marked successors 306 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_739_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_739_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_739_completed_
      -- 
    cpelement_group_983 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(985);
      marked_predecessors(0) <= cp_elements(989);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(983)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(983),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 984 transition  output  bypass 
    -- predecessors 307 
    -- successors 985 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_register/$entry
      -- 
    cp_elements(984) <= cp_elements(307);
    req_3851_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(984), ack => simple_obj_ref_735_inst_req_0); -- 
    -- CP-element group 985 transition  input  bypass 
    -- predecessors 984 
    -- successors 983 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_737_register/$exit
      -- 
    ack_3852_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_735_inst_ack_0, ack => cp_elements(985)); -- 
    -- CP-element group 986 join  fork  transition  bypass 
    -- predecessors 988 
    -- marked predecessors 992 
    -- successors 990 
    -- marked successors 307 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_742_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_742_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_742_completed_
      -- 
    cpelement_group_986 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(988);
      marked_predecessors(0) <= cp_elements(992);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(986)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(986),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 987 transition  output  bypass 
    -- predecessors 983 
    -- successors 988 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_register/req
      -- 
    cp_elements(987) <= cp_elements(983);
    req_3862_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(987), ack => simple_obj_ref_738_inst_req_0); -- 
    -- CP-element group 988 transition  input  bypass 
    -- predecessors 987 
    -- successors 986 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_740_register/$exit
      -- 
    ack_3863_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_738_inst_ack_0, ack => cp_elements(988)); -- 
    -- CP-element group 989 join  fork  transition  bypass 
    -- predecessors 991 
    -- marked predecessors 995 
    -- successors 993 
    -- marked successors 983 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_745_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_745_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_745_trigger_
      -- 
    cpelement_group_989 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(991);
      marked_predecessors(0) <= cp_elements(995);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(989)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(989),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 990 transition  output  bypass 
    -- predecessors 986 
    -- successors 991 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_register/req
      -- 
    cp_elements(990) <= cp_elements(986);
    req_3873_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(990), ack => simple_obj_ref_741_inst_req_0); -- 
    -- CP-element group 991 transition  input  bypass 
    -- predecessors 990 
    -- successors 989 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_743_register/ack
      -- 
    ack_3874_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_741_inst_ack_0, ack => cp_elements(991)); -- 
    -- CP-element group 992 join  fork  transition  bypass 
    -- predecessors 994 
    -- marked predecessors 999 
    -- successors 996 
    -- marked successors 986 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_748_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_748_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_748_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_completed_
      -- 
    cpelement_group_992 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(994);
      marked_predecessors(0) <= cp_elements(999);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(992)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(992),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 993 transition  output  bypass 
    -- predecessors 989 
    -- successors 994 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_register/req
      -- 
    cp_elements(993) <= cp_elements(989);
    req_3884_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(993), ack => simple_obj_ref_744_inst_req_0); -- 
    -- CP-element group 994 transition  input  bypass 
    -- predecessors 993 
    -- successors 992 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_746_register/ack
      -- 
    ack_3885_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_744_inst_ack_0, ack => cp_elements(994)); -- 
    -- CP-element group 995 fork  transition  bypass 
    -- predecessors 997 
    -- successors 1004 
    -- marked successors 989 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_750_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_750_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_750_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_active_
      -- 
    cp_elements(995) <= cp_elements(997);
    -- CP-element group 996 transition  output  bypass 
    -- predecessors 992 
    -- successors 997 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_register/req
      -- 
    cp_elements(996) <= cp_elements(992);
    req_3895_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(996), ack => simple_obj_ref_747_inst_req_0); -- 
    -- CP-element group 997 transition  input  bypass 
    -- predecessors 996 
    -- successors 995 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_749_register/ack
      -- 
    ack_3896_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_747_inst_ack_0, ack => cp_elements(997)); -- 
    -- CP-element group 998 join  transition  bypass 
    -- predecessors 967 1001 706 
    -- marked predecessors 999 
    -- successors 1010 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_trigger_
      -- 
    cpelement_group_998 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(967);
      predecessors(1) <= cp_elements(1001);
      predecessors(2) <= cp_elements(706);
      marked_predecessors(0) <= cp_elements(999);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(998)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(998),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 999 join  fork  transition  bypass 
    -- predecessors 1012 
    -- marked predecessors 1000 
    -- successors 1013 1030 
    -- marked successors 992 998 1002 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_active_
      -- 
    cpelement_group_999 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1012);
      marked_predecessors(0) <= cp_elements(1000);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(999)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(999),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1000 fork  transition  bypass 
    -- predecessors 1014 
    -- successors 1175 
    -- marked successors 999 709 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_753_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_completed_
      -- 
    cp_elements(1000) <= cp_elements(1014);
    -- CP-element group 1001 transition  bypass 
    -- predecessors 1009 
    -- successors 998 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_word_address_calculated
      -- 
    cp_elements(1001) <= cp_elements(1009);
    -- CP-element group 1002 join  transition  bypass 
    -- predecessors 1007 
    -- marked predecessors 999 
    -- successors 1008 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_root_address_calculated
      -- 
    cpelement_group_1002 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1007);
      marked_predecessors(0) <= cp_elements(999);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1002)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1002),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1003 transition  bypass 
    -- predecessors 1005 
    -- successors 1006 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_address_resized
      -- 
    cp_elements(1003) <= cp_elements(1005);
    -- CP-element group 1004 transition  output  bypass 
    -- predecessors 995 
    -- successors 1005 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_addr_resize/base_resize_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_addr_resize/$entry
      -- 
    cp_elements(1004) <= cp_elements(995);
    base_resize_req_3916_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1004), ack => ptr_deref_751_base_resize_req_0); -- 
    -- CP-element group 1005 transition  input  bypass 
    -- predecessors 1004 
    -- successors 1003 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_addr_resize/base_resize_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_addr_resize/$exit
      -- 
    base_resize_ack_3917_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_base_resize_ack_0, ack => cp_elements(1005)); -- 
    -- CP-element group 1006 transition  output  bypass 
    -- predecessors 1003 
    -- successors 1007 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_plus_offset/sum_rename_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_plus_offset/$entry
      -- 
    cp_elements(1006) <= cp_elements(1003);
    sum_rename_req_3921_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1006), ack => ptr_deref_751_root_address_inst_req_0); -- 
    -- CP-element group 1007 transition  input  bypass 
    -- predecessors 1006 
    -- successors 1002 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_3922_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_root_address_inst_ack_0, ack => cp_elements(1007)); -- 
    -- CP-element group 1008 transition  output  bypass 
    -- predecessors 1002 
    -- successors 1009 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_word_addrgen/root_register_req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_word_addrgen/$entry
      -- 
    cp_elements(1008) <= cp_elements(1002);
    root_register_req_3926_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1008), ack => ptr_deref_751_addr_0_req_0); -- 
    -- CP-element group 1009 transition  input  bypass 
    -- predecessors 1008 
    -- successors 1001 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_word_addrgen/root_register_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_word_addrgen/$exit
      -- 
    root_register_ack_3927_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_addr_0_ack_0, ack => cp_elements(1009)); -- 
    -- CP-element group 1010 transition  output  bypass 
    -- predecessors 998 
    -- successors 1011 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/split_req
      -- 
    cp_elements(1010) <= cp_elements(998);
    split_req_3931_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1010), ack => ptr_deref_751_gather_scatter_req_0); -- 
    -- CP-element group 1011 transition  input  output  bypass 
    -- predecessors 1010 
    -- successors 1012 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/word_access_0/rr
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/split_ack
      -- 
    split_ack_3932_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_gather_scatter_ack_0, ack => cp_elements(1011)); -- 
    rr_3939_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1011), ack => ptr_deref_751_store_0_req_0); -- 
    -- CP-element group 1012 transition  input  bypass 
    -- predecessors 1011 
    -- successors 999 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/word_access_0/ra
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_request/word_access/word_access_0/$exit
      -- 
    ra_3940_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_store_0_ack_0, ack => cp_elements(1012)); -- 
    -- CP-element group 1013 transition  output  bypass 
    -- predecessors 999 
    -- successors 1014 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/word_access_0/cr
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/$entry
      -- 
    cp_elements(1013) <= cp_elements(999);
    cr_3950_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1013), ack => ptr_deref_751_store_0_req_1); -- 
    -- CP-element group 1014 transition  input  bypass 
    -- predecessors 1013 
    -- successors 1000 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/word_access_0/ca
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_751_complete/word_access/word_access_0/$exit
      -- 
    ca_3951_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_751_store_0_ack_1, ack => cp_elements(1014)); -- 
    -- CP-element group 1015 join  fork  transition  bypass 
    -- predecessors 1017 
    -- marked predecessors 1021 
    -- successors 1019 
    -- marked successors 241 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_758_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_758_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_758_completed_
      -- 
    cpelement_group_1015 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1017);
      marked_predecessors(0) <= cp_elements(1021);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1015)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1015),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1016 transition  output  bypass 
    -- predecessors 242 
    -- successors 1017 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_register/$entry
      -- 
    cp_elements(1016) <= cp_elements(242);
    req_3961_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1016), ack => simple_obj_ref_754_inst_req_0); -- 
    -- CP-element group 1017 transition  input  bypass 
    -- predecessors 1016 
    -- successors 1015 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_756_register/$exit
      -- 
    ack_3962_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_754_inst_ack_0, ack => cp_elements(1017)); -- 
    -- CP-element group 1018 join  fork  transition  bypass 
    -- predecessors 1020 
    -- marked predecessors 1024 
    -- successors 1022 
    -- marked successors 242 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_761_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_761_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_761_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_trigger_
      -- 
    cpelement_group_1018 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1020);
      marked_predecessors(0) <= cp_elements(1024);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1018)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1018),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1019 transition  output  bypass 
    -- predecessors 1015 
    -- successors 1020 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_register/$entry
      -- 
    cp_elements(1019) <= cp_elements(1015);
    req_3972_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1019), ack => simple_obj_ref_757_inst_req_0); -- 
    -- CP-element group 1020 transition  input  bypass 
    -- predecessors 1019 
    -- successors 1018 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_759_register/ack
      -- 
    ack_3973_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_757_inst_ack_0, ack => cp_elements(1020)); -- 
    -- CP-element group 1021 join  fork  transition  bypass 
    -- predecessors 1023 
    -- marked predecessors 1027 
    -- successors 1025 
    -- marked successors 1015 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_764_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_764_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_764_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_active_
      -- 
    cpelement_group_1021 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1023);
      marked_predecessors(0) <= cp_elements(1027);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1021)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1021),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1022 transition  output  bypass 
    -- predecessors 1018 
    -- successors 1023 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_register/$entry
      -- 
    cp_elements(1022) <= cp_elements(1018);
    req_3983_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1022), ack => simple_obj_ref_760_inst_req_0); -- 
    -- CP-element group 1023 transition  input  bypass 
    -- predecessors 1022 
    -- successors 1021 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_register/ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_762_register/$exit
      -- 
    ack_3984_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_760_inst_ack_0, ack => cp_elements(1023)); -- 
    -- CP-element group 1024 join  fork  transition  bypass 
    -- predecessors 1026 
    -- marked predecessors 1031 
    -- successors 1028 
    -- marked successors 1018 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_767_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_767_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_767_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_active_
      -- 
    cpelement_group_1024 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1026);
      marked_predecessors(0) <= cp_elements(1031);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1024)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1024),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1025 transition  output  bypass 
    -- predecessors 1021 
    -- successors 1026 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_register/req
      -- 
    cp_elements(1025) <= cp_elements(1021);
    req_3994_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1025), ack => simple_obj_ref_763_inst_req_0); -- 
    -- CP-element group 1026 transition  input  bypass 
    -- predecessors 1025 
    -- successors 1024 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_765_register/ack
      -- 
    ack_3995_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_763_inst_ack_0, ack => cp_elements(1026)); -- 
    -- CP-element group 1027 fork  transition  bypass 
    -- predecessors 1029 
    -- successors 1036 
    -- marked successors 1021 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_769_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_769_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_769_completed_
      -- 
    cp_elements(1027) <= cp_elements(1029);
    -- CP-element group 1028 transition  output  bypass 
    -- predecessors 1024 
    -- successors 1029 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_register/req
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_register/$entry
      -- 
    cp_elements(1028) <= cp_elements(1024);
    req_4005_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1028), ack => simple_obj_ref_766_inst_req_0); -- 
    -- CP-element group 1029 transition  input  bypass 
    -- predecessors 1028 
    -- successors 1027 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_768_register/ack
      -- 
    ack_4006_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_766_inst_ack_0, ack => cp_elements(1029)); -- 
    -- CP-element group 1030 join  transition  bypass 
    -- predecessors 999 1033 749 
    -- marked predecessors 1031 
    -- successors 1042 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_trigger_
      -- 
    cpelement_group_1030 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(999);
      predecessors(1) <= cp_elements(1033);
      predecessors(2) <= cp_elements(749);
      marked_predecessors(0) <= cp_elements(1031);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1030)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1030),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1031 join  fork  transition  bypass 
    -- predecessors 1044 
    -- marked predecessors 1032 
    -- successors 1045 1062 
    -- marked successors 1024 1030 1034 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_active_
      -- 
    cpelement_group_1031 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1044);
      marked_predecessors(0) <= cp_elements(1032);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1031)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1031),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1032 fork  transition  bypass 
    -- predecessors 1046 
    -- successors 1175 
    -- marked successors 752 1031 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_772_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_completed_
      -- 
    cp_elements(1032) <= cp_elements(1046);
    -- CP-element group 1033 transition  bypass 
    -- predecessors 1041 
    -- successors 1030 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_word_address_calculated
      -- 
    cp_elements(1033) <= cp_elements(1041);
    -- CP-element group 1034 join  transition  bypass 
    -- predecessors 1039 
    -- marked predecessors 1031 
    -- successors 1040 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_root_address_calculated
      -- 
    cpelement_group_1034 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1039);
      marked_predecessors(0) <= cp_elements(1031);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1034)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1034),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1035 transition  bypass 
    -- predecessors 1037 
    -- successors 1038 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_address_resized
      -- 
    cp_elements(1035) <= cp_elements(1037);
    -- CP-element group 1036 transition  output  bypass 
    -- predecessors 1027 
    -- successors 1037 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_addr_resize/base_resize_req
      -- 
    cp_elements(1036) <= cp_elements(1027);
    base_resize_req_4026_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1036), ack => ptr_deref_770_base_resize_req_0); -- 
    -- CP-element group 1037 transition  input  bypass 
    -- predecessors 1036 
    -- successors 1035 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_4027_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_base_resize_ack_0, ack => cp_elements(1037)); -- 
    -- CP-element group 1038 transition  output  bypass 
    -- predecessors 1035 
    -- successors 1039 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_plus_offset/sum_rename_req
      -- 
    cp_elements(1038) <= cp_elements(1035);
    sum_rename_req_4031_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1038), ack => ptr_deref_770_root_address_inst_req_0); -- 
    -- CP-element group 1039 transition  input  bypass 
    -- predecessors 1038 
    -- successors 1034 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4032_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_root_address_inst_ack_0, ack => cp_elements(1039)); -- 
    -- CP-element group 1040 transition  output  bypass 
    -- predecessors 1034 
    -- successors 1041 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_word_addrgen/root_register_req
      -- 
    cp_elements(1040) <= cp_elements(1034);
    root_register_req_4036_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1040), ack => ptr_deref_770_addr_0_req_0); -- 
    -- CP-element group 1041 transition  input  bypass 
    -- predecessors 1040 
    -- successors 1033 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_word_addrgen/root_register_ack
      -- 
    root_register_ack_4037_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_addr_0_ack_0, ack => cp_elements(1041)); -- 
    -- CP-element group 1042 transition  output  bypass 
    -- predecessors 1030 
    -- successors 1043 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/split_req
      -- 
    cp_elements(1042) <= cp_elements(1030);
    split_req_4041_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1042), ack => ptr_deref_770_gather_scatter_req_0); -- 
    -- CP-element group 1043 transition  input  output  bypass 
    -- predecessors 1042 
    -- successors 1044 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/word_access_0/rr
      -- 
    split_ack_4042_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_gather_scatter_ack_0, ack => cp_elements(1043)); -- 
    rr_4049_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1043), ack => ptr_deref_770_store_0_req_0); -- 
    -- CP-element group 1044 transition  input  bypass 
    -- predecessors 1043 
    -- successors 1031 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_request/word_access/word_access_0/ra
      -- 
    ra_4050_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_store_0_ack_0, ack => cp_elements(1044)); -- 
    -- CP-element group 1045 transition  output  bypass 
    -- predecessors 1031 
    -- successors 1046 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1045) <= cp_elements(1031);
    cr_4060_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1045), ack => ptr_deref_770_store_0_req_1); -- 
    -- CP-element group 1046 transition  input  bypass 
    -- predecessors 1045 
    -- successors 1032 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_770_complete/word_access/word_access_0/ca
      -- 
    ca_4061_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_770_store_0_ack_1, ack => cp_elements(1046)); -- 
    -- CP-element group 1047 join  fork  transition  bypass 
    -- predecessors 1049 
    -- marked predecessors 1053 
    -- successors 1051 
    -- marked successors 176 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_777_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_777_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_777_completed_
      -- 
    cpelement_group_1047 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1049);
      marked_predecessors(0) <= cp_elements(1053);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1047)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1047),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1048 transition  output  bypass 
    -- predecessors 177 
    -- successors 1049 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_register/req
      -- 
    cp_elements(1048) <= cp_elements(177);
    req_4071_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1048), ack => simple_obj_ref_773_inst_req_0); -- 
    -- CP-element group 1049 transition  input  bypass 
    -- predecessors 1048 
    -- successors 1047 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_775_register/ack
      -- 
    ack_4072_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_773_inst_ack_0, ack => cp_elements(1049)); -- 
    -- CP-element group 1050 join  fork  transition  bypass 
    -- predecessors 1052 
    -- marked predecessors 1056 
    -- successors 1054 
    -- marked successors 177 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_780_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_780_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_780_completed_
      -- 
    cpelement_group_1050 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1052);
      marked_predecessors(0) <= cp_elements(1056);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1050)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1050),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1051 transition  output  bypass 
    -- predecessors 1047 
    -- successors 1052 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_register/req
      -- 
    cp_elements(1051) <= cp_elements(1047);
    req_4082_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1051), ack => simple_obj_ref_776_inst_req_0); -- 
    -- CP-element group 1052 transition  input  bypass 
    -- predecessors 1051 
    -- successors 1050 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_778_register/ack
      -- 
    ack_4083_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_776_inst_ack_0, ack => cp_elements(1052)); -- 
    -- CP-element group 1053 join  fork  transition  bypass 
    -- predecessors 1055 
    -- marked predecessors 1059 
    -- successors 1057 
    -- marked successors 1047 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_783_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_783_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_783_completed_
      -- 
    cpelement_group_1053 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1055);
      marked_predecessors(0) <= cp_elements(1059);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1053)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1053),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1054 transition  output  bypass 
    -- predecessors 1050 
    -- successors 1055 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_register/req
      -- 
    cp_elements(1054) <= cp_elements(1050);
    req_4093_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1054), ack => simple_obj_ref_779_inst_req_0); -- 
    -- CP-element group 1055 transition  input  bypass 
    -- predecessors 1054 
    -- successors 1053 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_781_register/ack
      -- 
    ack_4094_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_779_inst_ack_0, ack => cp_elements(1055)); -- 
    -- CP-element group 1056 join  fork  transition  bypass 
    -- predecessors 1058 
    -- marked predecessors 1063 
    -- successors 1060 
    -- marked successors 1050 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_786_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_786_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_786_completed_
      -- 
    cpelement_group_1056 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1058);
      marked_predecessors(0) <= cp_elements(1063);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1056)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1056),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1057 transition  output  bypass 
    -- predecessors 1053 
    -- successors 1058 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_register/req
      -- 
    cp_elements(1057) <= cp_elements(1053);
    req_4104_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1057), ack => simple_obj_ref_782_inst_req_0); -- 
    -- CP-element group 1058 transition  input  bypass 
    -- predecessors 1057 
    -- successors 1056 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_784_register/ack
      -- 
    ack_4105_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_782_inst_ack_0, ack => cp_elements(1058)); -- 
    -- CP-element group 1059 fork  transition  bypass 
    -- predecessors 1061 
    -- successors 1068 
    -- marked successors 1053 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_788_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_788_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_788_completed_
      -- 
    cp_elements(1059) <= cp_elements(1061);
    -- CP-element group 1060 transition  output  bypass 
    -- predecessors 1056 
    -- successors 1061 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_register/req
      -- 
    cp_elements(1060) <= cp_elements(1056);
    req_4115_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1060), ack => simple_obj_ref_785_inst_req_0); -- 
    -- CP-element group 1061 transition  input  bypass 
    -- predecessors 1060 
    -- successors 1059 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_787_register/ack
      -- 
    ack_4116_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_785_inst_ack_0, ack => cp_elements(1061)); -- 
    -- CP-element group 1062 join  transition  bypass 
    -- predecessors 792 1031 1065 
    -- marked predecessors 1063 
    -- successors 1074 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_trigger_
      -- 
    cpelement_group_1062 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(792);
      predecessors(1) <= cp_elements(1031);
      predecessors(2) <= cp_elements(1065);
      marked_predecessors(0) <= cp_elements(1063);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1062)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1062),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1063 join  fork  transition  bypass 
    -- predecessors 1076 
    -- marked predecessors 1064 
    -- successors 1094 1077 
    -- marked successors 1056 1062 1066 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_active_
      -- 
    cpelement_group_1063 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1076);
      marked_predecessors(0) <= cp_elements(1064);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1063)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1063),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1064 fork  transition  bypass 
    -- predecessors 1078 
    -- successors 1175 
    -- marked successors 795 1063 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_791_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_completed_
      -- 
    cp_elements(1064) <= cp_elements(1078);
    -- CP-element group 1065 transition  bypass 
    -- predecessors 1073 
    -- successors 1062 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_word_address_calculated
      -- 
    cp_elements(1065) <= cp_elements(1073);
    -- CP-element group 1066 join  transition  bypass 
    -- predecessors 1071 
    -- marked predecessors 1063 
    -- successors 1072 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_root_address_calculated
      -- 
    cpelement_group_1066 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1071);
      marked_predecessors(0) <= cp_elements(1063);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1066)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1066),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1067 transition  bypass 
    -- predecessors 1069 
    -- successors 1070 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_address_resized
      -- 
    cp_elements(1067) <= cp_elements(1069);
    -- CP-element group 1068 transition  output  bypass 
    -- predecessors 1059 
    -- successors 1069 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_addr_resize/base_resize_req
      -- 
    cp_elements(1068) <= cp_elements(1059);
    base_resize_req_4136_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1068), ack => ptr_deref_789_base_resize_req_0); -- 
    -- CP-element group 1069 transition  input  bypass 
    -- predecessors 1068 
    -- successors 1067 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_4137_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_base_resize_ack_0, ack => cp_elements(1069)); -- 
    -- CP-element group 1070 transition  output  bypass 
    -- predecessors 1067 
    -- successors 1071 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_plus_offset/sum_rename_req
      -- 
    cp_elements(1070) <= cp_elements(1067);
    sum_rename_req_4141_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1070), ack => ptr_deref_789_root_address_inst_req_0); -- 
    -- CP-element group 1071 transition  input  bypass 
    -- predecessors 1070 
    -- successors 1066 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4142_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_root_address_inst_ack_0, ack => cp_elements(1071)); -- 
    -- CP-element group 1072 transition  output  bypass 
    -- predecessors 1066 
    -- successors 1073 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_word_addrgen/root_register_req
      -- 
    cp_elements(1072) <= cp_elements(1066);
    root_register_req_4146_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1072), ack => ptr_deref_789_addr_0_req_0); -- 
    -- CP-element group 1073 transition  input  bypass 
    -- predecessors 1072 
    -- successors 1065 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_word_addrgen/root_register_ack
      -- 
    root_register_ack_4147_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_addr_0_ack_0, ack => cp_elements(1073)); -- 
    -- CP-element group 1074 transition  output  bypass 
    -- predecessors 1062 
    -- successors 1075 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/split_req
      -- 
    cp_elements(1074) <= cp_elements(1062);
    split_req_4151_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1074), ack => ptr_deref_789_gather_scatter_req_0); -- 
    -- CP-element group 1075 transition  input  output  bypass 
    -- predecessors 1074 
    -- successors 1076 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/word_access_0/rr
      -- 
    split_ack_4152_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_gather_scatter_ack_0, ack => cp_elements(1075)); -- 
    rr_4159_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1075), ack => ptr_deref_789_store_0_req_0); -- 
    -- CP-element group 1076 transition  input  bypass 
    -- predecessors 1075 
    -- successors 1063 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_request/word_access/word_access_0/ra
      -- 
    ra_4160_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_store_0_ack_0, ack => cp_elements(1076)); -- 
    -- CP-element group 1077 transition  output  bypass 
    -- predecessors 1063 
    -- successors 1078 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1077) <= cp_elements(1063);
    cr_4170_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1077), ack => ptr_deref_789_store_0_req_1); -- 
    -- CP-element group 1078 transition  input  bypass 
    -- predecessors 1077 
    -- successors 1064 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_789_complete/word_access/word_access_0/ca
      -- 
    ca_4171_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_789_store_0_ack_1, ack => cp_elements(1078)); -- 
    -- CP-element group 1079 join  fork  transition  bypass 
    -- predecessors 1081 
    -- marked predecessors 1085 
    -- successors 1083 
    -- marked successors 111 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_796_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_796_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_796_completed_
      -- 
    cpelement_group_1079 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1081);
      marked_predecessors(0) <= cp_elements(1085);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1079)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1079),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1080 transition  output  bypass 
    -- predecessors 112 
    -- successors 1081 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_register/req
      -- 
    cp_elements(1080) <= cp_elements(112);
    req_4181_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1080), ack => simple_obj_ref_792_inst_req_0); -- 
    -- CP-element group 1081 transition  input  bypass 
    -- predecessors 1080 
    -- successors 1079 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_794_register/ack
      -- 
    ack_4182_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_792_inst_ack_0, ack => cp_elements(1081)); -- 
    -- CP-element group 1082 join  fork  transition  bypass 
    -- predecessors 1084 
    -- marked predecessors 1088 
    -- successors 1086 
    -- marked successors 112 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_799_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_799_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_799_completed_
      -- 
    cpelement_group_1082 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1084);
      marked_predecessors(0) <= cp_elements(1088);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1082)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1082),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1083 transition  output  bypass 
    -- predecessors 1079 
    -- successors 1084 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_register/req
      -- 
    cp_elements(1083) <= cp_elements(1079);
    req_4192_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1083), ack => simple_obj_ref_795_inst_req_0); -- 
    -- CP-element group 1084 transition  input  bypass 
    -- predecessors 1083 
    -- successors 1082 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_797_register/ack
      -- 
    ack_4193_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_795_inst_ack_0, ack => cp_elements(1084)); -- 
    -- CP-element group 1085 join  fork  transition  bypass 
    -- predecessors 1087 
    -- marked predecessors 1091 
    -- successors 1089 
    -- marked successors 1079 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_802_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_802_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_802_completed_
      -- 
    cpelement_group_1085 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1087);
      marked_predecessors(0) <= cp_elements(1091);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1085)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1085),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1086 transition  output  bypass 
    -- predecessors 1082 
    -- successors 1087 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_register/req
      -- 
    cp_elements(1086) <= cp_elements(1082);
    req_4203_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1086), ack => simple_obj_ref_798_inst_req_0); -- 
    -- CP-element group 1087 transition  input  bypass 
    -- predecessors 1086 
    -- successors 1085 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_800_register/ack
      -- 
    ack_4204_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_798_inst_ack_0, ack => cp_elements(1087)); -- 
    -- CP-element group 1088 join  fork  transition  bypass 
    -- predecessors 1090 
    -- marked predecessors 1095 
    -- successors 1092 
    -- marked successors 1082 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_805_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_805_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_805_completed_
      -- 
    cpelement_group_1088 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1090);
      marked_predecessors(0) <= cp_elements(1095);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1088)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1088),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1089 transition  output  bypass 
    -- predecessors 1085 
    -- successors 1090 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_register/req
      -- 
    cp_elements(1089) <= cp_elements(1085);
    req_4214_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1089), ack => simple_obj_ref_801_inst_req_0); -- 
    -- CP-element group 1090 transition  input  bypass 
    -- predecessors 1089 
    -- successors 1088 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_803_register/ack
      -- 
    ack_4215_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_801_inst_ack_0, ack => cp_elements(1090)); -- 
    -- CP-element group 1091 fork  transition  bypass 
    -- predecessors 1093 
    -- successors 1100 
    -- marked successors 1085 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_807_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_807_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_807_completed_
      -- 
    cp_elements(1091) <= cp_elements(1093);
    -- CP-element group 1092 transition  output  bypass 
    -- predecessors 1088 
    -- successors 1093 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_register/req
      -- 
    cp_elements(1092) <= cp_elements(1088);
    req_4225_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1092), ack => simple_obj_ref_804_inst_req_0); -- 
    -- CP-element group 1093 transition  input  bypass 
    -- predecessors 1092 
    -- successors 1091 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_806_register/ack
      -- 
    ack_4226_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_804_inst_ack_0, ack => cp_elements(1093)); -- 
    -- CP-element group 1094 join  transition  bypass 
    -- predecessors 1097 835 1063 
    -- marked predecessors 1095 
    -- successors 1106 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_trigger_
      -- 
    cpelement_group_1094 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1097);
      predecessors(1) <= cp_elements(835);
      predecessors(2) <= cp_elements(1063);
      marked_predecessors(0) <= cp_elements(1095);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1094)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1094),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1095 join  fork  transition  bypass 
    -- predecessors 1108 
    -- marked predecessors 1096 
    -- successors 1109 1126 
    -- marked successors 1094 1098 1088 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_active_
      -- 
    cpelement_group_1095 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1108);
      marked_predecessors(0) <= cp_elements(1096);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1095)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1095),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1096 fork  transition  bypass 
    -- predecessors 1110 
    -- successors 1175 
    -- marked successors 1095 838 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_810_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_completed_
      -- 
    cp_elements(1096) <= cp_elements(1110);
    -- CP-element group 1097 transition  bypass 
    -- predecessors 1105 
    -- successors 1094 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_word_address_calculated
      -- 
    cp_elements(1097) <= cp_elements(1105);
    -- CP-element group 1098 join  transition  bypass 
    -- predecessors 1103 
    -- marked predecessors 1095 
    -- successors 1104 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_root_address_calculated
      -- 
    cpelement_group_1098 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1103);
      marked_predecessors(0) <= cp_elements(1095);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1098)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1098),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1099 transition  bypass 
    -- predecessors 1101 
    -- successors 1102 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_address_resized
      -- 
    cp_elements(1099) <= cp_elements(1101);
    -- CP-element group 1100 transition  output  bypass 
    -- predecessors 1091 
    -- successors 1101 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_addr_resize/base_resize_req
      -- 
    cp_elements(1100) <= cp_elements(1091);
    base_resize_req_4246_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1100), ack => ptr_deref_808_base_resize_req_0); -- 
    -- CP-element group 1101 transition  input  bypass 
    -- predecessors 1100 
    -- successors 1099 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_4247_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_base_resize_ack_0, ack => cp_elements(1101)); -- 
    -- CP-element group 1102 transition  output  bypass 
    -- predecessors 1099 
    -- successors 1103 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_plus_offset/sum_rename_req
      -- 
    cp_elements(1102) <= cp_elements(1099);
    sum_rename_req_4251_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1102), ack => ptr_deref_808_root_address_inst_req_0); -- 
    -- CP-element group 1103 transition  input  bypass 
    -- predecessors 1102 
    -- successors 1098 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4252_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_root_address_inst_ack_0, ack => cp_elements(1103)); -- 
    -- CP-element group 1104 transition  output  bypass 
    -- predecessors 1098 
    -- successors 1105 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_word_addrgen/root_register_req
      -- 
    cp_elements(1104) <= cp_elements(1098);
    root_register_req_4256_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1104), ack => ptr_deref_808_addr_0_req_0); -- 
    -- CP-element group 1105 transition  input  bypass 
    -- predecessors 1104 
    -- successors 1097 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_word_addrgen/root_register_ack
      -- 
    root_register_ack_4257_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_addr_0_ack_0, ack => cp_elements(1105)); -- 
    -- CP-element group 1106 transition  output  bypass 
    -- predecessors 1094 
    -- successors 1107 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/split_req
      -- 
    cp_elements(1106) <= cp_elements(1094);
    split_req_4261_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1106), ack => ptr_deref_808_gather_scatter_req_0); -- 
    -- CP-element group 1107 transition  input  output  bypass 
    -- predecessors 1106 
    -- successors 1108 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/word_access_0/rr
      -- 
    split_ack_4262_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_gather_scatter_ack_0, ack => cp_elements(1107)); -- 
    rr_4269_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1107), ack => ptr_deref_808_store_0_req_0); -- 
    -- CP-element group 1108 transition  input  bypass 
    -- predecessors 1107 
    -- successors 1095 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_request/word_access/word_access_0/ra
      -- 
    ra_4270_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_store_0_ack_0, ack => cp_elements(1108)); -- 
    -- CP-element group 1109 transition  output  bypass 
    -- predecessors 1095 
    -- successors 1110 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1109) <= cp_elements(1095);
    cr_4280_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1109), ack => ptr_deref_808_store_0_req_1); -- 
    -- CP-element group 1110 transition  input  bypass 
    -- predecessors 1109 
    -- successors 1096 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_808_complete/word_access/word_access_0/ca
      -- 
    ca_4281_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_808_store_0_ack_1, ack => cp_elements(1110)); -- 
    -- CP-element group 1111 join  fork  transition  bypass 
    -- predecessors 1113 
    -- marked predecessors 1117 
    -- successors 1115 
    -- marked successors 46 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_815_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_815_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_815_completed_
      -- 
    cpelement_group_1111 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1113);
      marked_predecessors(0) <= cp_elements(1117);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1111)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1111),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1112 transition  output  bypass 
    -- predecessors 47 
    -- successors 1113 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_register/req
      -- 
    cp_elements(1112) <= cp_elements(47);
    req_4291_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1112), ack => simple_obj_ref_811_inst_req_0); -- 
    -- CP-element group 1113 transition  input  bypass 
    -- predecessors 1112 
    -- successors 1111 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_813_register/ack
      -- 
    ack_4292_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_811_inst_ack_0, ack => cp_elements(1113)); -- 
    -- CP-element group 1114 join  fork  transition  bypass 
    -- predecessors 1116 
    -- marked predecessors 1120 
    -- successors 1118 
    -- marked successors 47 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_818_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_818_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_818_completed_
      -- 
    cpelement_group_1114 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1116);
      marked_predecessors(0) <= cp_elements(1120);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1114)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1114),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1115 transition  output  bypass 
    -- predecessors 1111 
    -- successors 1116 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_register/req
      -- 
    cp_elements(1115) <= cp_elements(1111);
    req_4302_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1115), ack => simple_obj_ref_814_inst_req_0); -- 
    -- CP-element group 1116 transition  input  bypass 
    -- predecessors 1115 
    -- successors 1114 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_816_register/ack
      -- 
    ack_4303_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_814_inst_ack_0, ack => cp_elements(1116)); -- 
    -- CP-element group 1117 join  fork  transition  bypass 
    -- predecessors 1119 
    -- marked predecessors 1123 
    -- successors 1121 
    -- marked successors 1111 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_821_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_821_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_821_completed_
      -- 
    cpelement_group_1117 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1119);
      marked_predecessors(0) <= cp_elements(1123);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1117)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1117),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1118 transition  output  bypass 
    -- predecessors 1114 
    -- successors 1119 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_register/req
      -- 
    cp_elements(1118) <= cp_elements(1114);
    req_4313_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1118), ack => simple_obj_ref_817_inst_req_0); -- 
    -- CP-element group 1119 transition  input  bypass 
    -- predecessors 1118 
    -- successors 1117 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_819_register/ack
      -- 
    ack_4314_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_817_inst_ack_0, ack => cp_elements(1119)); -- 
    -- CP-element group 1120 join  fork  transition  bypass 
    -- predecessors 1122 
    -- marked predecessors 1127 
    -- successors 1124 
    -- marked successors 1114 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_824_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_824_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_824_completed_
      -- 
    cpelement_group_1120 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1122);
      marked_predecessors(0) <= cp_elements(1127);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1120)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1120),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1121 transition  output  bypass 
    -- predecessors 1117 
    -- successors 1122 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_register/req
      -- 
    cp_elements(1121) <= cp_elements(1117);
    req_4324_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1121), ack => simple_obj_ref_820_inst_req_0); -- 
    -- CP-element group 1122 transition  input  bypass 
    -- predecessors 1121 
    -- successors 1120 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_822_register/ack
      -- 
    ack_4325_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_820_inst_ack_0, ack => cp_elements(1122)); -- 
    -- CP-element group 1123 fork  transition  bypass 
    -- predecessors 1125 
    -- successors 1132 
    -- marked successors 1117 
    -- members (6) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_address_calculated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_826_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_826_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_826_completed_
      -- 
    cp_elements(1123) <= cp_elements(1125);
    -- CP-element group 1124 transition  output  bypass 
    -- predecessors 1120 
    -- successors 1125 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_register/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_register/req
      -- 
    cp_elements(1124) <= cp_elements(1120);
    req_4335_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1124), ack => simple_obj_ref_823_inst_req_0); -- 
    -- CP-element group 1125 transition  input  bypass 
    -- predecessors 1124 
    -- successors 1123 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_register/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_825_register/ack
      -- 
    ack_4336_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => simple_obj_ref_823_inst_ack_0, ack => cp_elements(1125)); -- 
    -- CP-element group 1126 join  transition  bypass 
    -- predecessors 878 1095 1129 
    -- marked predecessors 1127 
    -- successors 1138 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_trigger_
      -- 
    cpelement_group_1126 : Block -- 
      signal predecessors: BooleanArray(2 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(878);
      predecessors(1) <= cp_elements(1095);
      predecessors(2) <= cp_elements(1129);
      marked_predecessors(0) <= cp_elements(1127);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1126)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1126),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1127 join  fork  transition  bypass 
    -- predecessors 1140 
    -- marked predecessors 1128 
    -- successors 1141 1174 
    -- marked successors 1120 1126 1130 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_active_
      -- 
    cpelement_group_1127 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1140);
      marked_predecessors(0) <= cp_elements(1128);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1127)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1127),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1128 fork  transition  bypass 
    -- predecessors 1142 
    -- successors 1175 
    -- marked successors 881 1127 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_829_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_completed_
      -- 
    cp_elements(1128) <= cp_elements(1142);
    -- CP-element group 1129 transition  bypass 
    -- predecessors 1137 
    -- successors 1126 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_word_address_calculated
      -- 
    cp_elements(1129) <= cp_elements(1137);
    -- CP-element group 1130 join  transition  bypass 
    -- predecessors 1135 
    -- marked predecessors 1127 
    -- successors 1136 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_root_address_calculated
      -- 
    cpelement_group_1130 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1135);
      marked_predecessors(0) <= cp_elements(1127);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1130)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1130),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1131 transition  bypass 
    -- predecessors 1133 
    -- successors 1134 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_address_resized
      -- 
    cp_elements(1131) <= cp_elements(1133);
    -- CP-element group 1132 transition  output  bypass 
    -- predecessors 1123 
    -- successors 1133 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_addr_resize/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_addr_resize/base_resize_req
      -- 
    cp_elements(1132) <= cp_elements(1123);
    base_resize_req_4356_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1132), ack => ptr_deref_827_base_resize_req_0); -- 
    -- CP-element group 1133 transition  input  bypass 
    -- predecessors 1132 
    -- successors 1131 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_addr_resize/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_addr_resize/base_resize_ack
      -- 
    base_resize_ack_4357_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_base_resize_ack_0, ack => cp_elements(1133)); -- 
    -- CP-element group 1134 transition  output  bypass 
    -- predecessors 1131 
    -- successors 1135 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_plus_offset/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_plus_offset/sum_rename_req
      -- 
    cp_elements(1134) <= cp_elements(1131);
    sum_rename_req_4361_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1134), ack => ptr_deref_827_root_address_inst_req_0); -- 
    -- CP-element group 1135 transition  input  bypass 
    -- predecessors 1134 
    -- successors 1130 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_plus_offset/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_base_plus_offset/sum_rename_ack
      -- 
    sum_rename_ack_4362_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_root_address_inst_ack_0, ack => cp_elements(1135)); -- 
    -- CP-element group 1136 transition  output  bypass 
    -- predecessors 1130 
    -- successors 1137 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_word_addrgen/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_word_addrgen/root_register_req
      -- 
    cp_elements(1136) <= cp_elements(1130);
    root_register_req_4366_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1136), ack => ptr_deref_827_addr_0_req_0); -- 
    -- CP-element group 1137 transition  input  bypass 
    -- predecessors 1136 
    -- successors 1129 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_word_addrgen/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_word_addrgen/root_register_ack
      -- 
    root_register_ack_4367_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_addr_0_ack_0, ack => cp_elements(1137)); -- 
    -- CP-element group 1138 transition  output  bypass 
    -- predecessors 1126 
    -- successors 1139 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/split_req
      -- 
    cp_elements(1138) <= cp_elements(1126);
    split_req_4371_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1138), ack => ptr_deref_827_gather_scatter_req_0); -- 
    -- CP-element group 1139 transition  input  output  bypass 
    -- predecessors 1138 
    -- successors 1140 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/split_ack
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/word_access_0/rr
      -- 
    split_ack_4372_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_gather_scatter_ack_0, ack => cp_elements(1139)); -- 
    rr_4379_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1139), ack => ptr_deref_827_store_0_req_0); -- 
    -- CP-element group 1140 transition  input  bypass 
    -- predecessors 1139 
    -- successors 1127 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_request/word_access/word_access_0/ra
      -- 
    ra_4380_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_store_0_ack_0, ack => cp_elements(1140)); -- 
    -- CP-element group 1141 transition  output  bypass 
    -- predecessors 1127 
    -- successors 1142 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/word_access_0/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/word_access_0/cr
      -- 
    cp_elements(1141) <= cp_elements(1127);
    cr_4390_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1141), ack => ptr_deref_827_store_0_req_1); -- 
    -- CP-element group 1142 transition  input  bypass 
    -- predecessors 1141 
    -- successors 1128 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/word_access_0/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ptr_deref_827_complete/word_access/word_access_0/ca
      -- 
    ca_4391_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => ptr_deref_827_store_0_ack_1, ack => cp_elements(1142)); -- 
    -- CP-element group 1143 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_active_
      -- 
    cp_elements(1143) <= cp_elements(7);
    -- CP-element group 1144 join  fork  transition  bypass 
    -- predecessors 1146 1148 
    -- successors 1156 1158 
    -- marked successors 19 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_835_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_835_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_835_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_837_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_837_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_837_completed_
      -- 
    cpelement_group_1144 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1146);
      predecessors(1) <= cp_elements(1148);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1144)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1144),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1145 join  transition  bypass 
    -- predecessors 1149 
    -- marked predecessors 1146 
    -- successors 1150 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_sample_start_
      -- 
    cpelement_group_1145 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1149);
      marked_predecessors(0) <= cp_elements(1146);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1145)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1145),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1146 fork  transition  bypass 
    -- predecessors 1151 
    -- successors 1144 
    -- marked successors 17 1145 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_sample_completed_
      -- 
    cp_elements(1146) <= cp_elements(1151);
    -- CP-element group 1147 join  transition  bypass 
    -- predecessors 1149 
    -- marked predecessors 1157 
    -- successors 1152 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_update_start_
      -- 
    cpelement_group_1147 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1149);
      marked_predecessors(0) <= cp_elements(1157);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1147)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1147),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1148 transition  bypass 
    -- predecessors 1153 
    -- successors 1144 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_update_completed_
      -- 
    cp_elements(1148) <= cp_elements(1153);
    -- CP-element group 1149 fork  transition  bypass 
    -- predecessors 15 
    -- successors 1145 1147 
    -- members (4) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_831_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_831_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_831_completed_
      -- 
    cp_elements(1149) <= cp_elements(15);
    -- CP-element group 1150 transition  output  bypass 
    -- predecessors 1145 
    -- successors 1151 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Sample/rr
      -- 
    cp_elements(1150) <= cp_elements(1145);
    rr_4408_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1150), ack => binary_834_inst_req_0); -- 
    -- CP-element group 1151 transition  input  bypass 
    -- predecessors 1150 
    -- successors 1146 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Sample/ra
      -- 
    ra_4409_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_834_inst_ack_0, ack => cp_elements(1151)); -- 
    -- CP-element group 1152 transition  output  bypass 
    -- predecessors 1147 
    -- successors 1153 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Update/cr
      -- 
    cp_elements(1152) <= cp_elements(1147);
    cr_4413_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1152), ack => binary_834_inst_req_1); -- 
    -- CP-element group 1153 transition  input  bypass 
    -- predecessors 1152 
    -- successors 1148 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_834_Update/ca
      -- 
    ca_4414_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_834_inst_ack_1, ack => cp_elements(1153)); -- 
    -- CP-element group 1154 transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_active_
      -- 
    cp_elements(1154) <= cp_elements(7);
    -- CP-element group 1155 join  fork  transition  bypass 
    -- predecessors 1157 1159 
    -- successors 1166 1168 
    -- marked successors 1158 
    -- members (8) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_841_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_841_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/assign_stmt_841_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_completed_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_843_trigger_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_843_active_
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/simple_obj_ref_843_completed_
      -- 
    cpelement_group_1155 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1157);
      predecessors(1) <= cp_elements(1159);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1155)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1155),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1156 join  transition  bypass 
    -- predecessors 1144 
    -- marked predecessors 1157 
    -- successors 1160 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_sample_start_
      -- 
    cpelement_group_1156 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1144);
      marked_predecessors(0) <= cp_elements(1157);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1156)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1156),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1157 fork  transition  bypass 
    -- predecessors 1161 
    -- successors 1155 
    -- marked successors 1147 1156 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_sample_completed_
      -- 
    cp_elements(1157) <= cp_elements(1161);
    -- CP-element group 1158 join  transition  bypass 
    -- predecessors 1144 
    -- marked predecessors 1155 1164 
    -- successors 1162 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_update_start_
      -- 
    cpelement_group_1158 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1144);
      marked_predecessors(0) <= cp_elements(1155);
      marked_predecessors(1) <= cp_elements(1164);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1158)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1158),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1159 transition  bypass 
    -- predecessors 1163 
    -- successors 1155 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_update_completed_
      -- 
    cp_elements(1159) <= cp_elements(1163);
    -- CP-element group 1160 transition  output  bypass 
    -- predecessors 1156 
    -- successors 1161 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Sample/rr
      -- 
    cp_elements(1160) <= cp_elements(1156);
    rr_4431_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1160), ack => binary_840_inst_req_0); -- 
    -- CP-element group 1161 transition  input  bypass 
    -- predecessors 1160 
    -- successors 1157 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Sample/ra
      -- 
    ra_4432_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_840_inst_ack_0, ack => cp_elements(1161)); -- 
    -- CP-element group 1162 transition  output  bypass 
    -- predecessors 1158 
    -- successors 1163 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Update/cr
      -- 
    cp_elements(1162) <= cp_elements(1158);
    cr_4436_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1162), ack => binary_840_inst_req_1); -- 
    -- CP-element group 1163 transition  input  bypass 
    -- predecessors 1162 
    -- successors 1159 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/binary_840_Update/ca
      -- 
    ca_4437_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => binary_840_inst_ack_1, ack => cp_elements(1163)); -- 
    -- CP-element group 1164 fork  transition  bypass 
    -- predecessors 7 
    -- successors 1175 
    -- marked successors 1158 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_active_
      -- 
    cp_elements(1164) <= cp_elements(7);
    -- CP-element group 1165 join  transition  output  bypass 
    -- predecessors 1167 1169 
    -- successors 3 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/condition_evaluated
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_completed_
      -- 
    cpelement_group_1165 : Block -- 
      signal predecessors: BooleanArray(1 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1167);
      predecessors(1) <= cp_elements(1169);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1165)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1165),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    condition_evaluated_4438_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1165), ack => do_while_stmt_398_branch_req_0); -- 
    -- CP-element group 1166 join  transition  bypass 
    -- predecessors 1155 
    -- marked predecessors 1167 
    -- successors 1170 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_sample_start_
      -- 
    cpelement_group_1166 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1155);
      marked_predecessors(0) <= cp_elements(1167);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1166)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1166),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1167 fork  transition  bypass 
    -- predecessors 1171 
    -- successors 1165 
    -- marked successors 1166 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_sample_completed_
      -- 
    cp_elements(1167) <= cp_elements(1171);
    -- CP-element group 1168 join  transition  bypass 
    -- predecessors 1155 
    -- marked predecessors 1169 
    -- successors 1172 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_update_start_
      -- 
    cpelement_group_1168 : Block -- 
      signal predecessors: BooleanArray(0 downto 0);
      signal marked_predecessors: BooleanArray(0 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(1155);
      marked_predecessors(0) <= cp_elements(1169);
      jNoI: marked_join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1168)_join")
        port map( -- 
          preds => predecessors,
          marked_preds => marked_predecessors,
          symbol_out => cp_elements(1168),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1169 fork  transition  bypass 
    -- predecessors 1173 
    -- successors 1165 
    -- marked successors 1168 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_update_completed_
      -- 
    cp_elements(1169) <= cp_elements(1173);
    -- CP-element group 1170 transition  output  bypass 
    -- predecessors 1166 
    -- successors 1171 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Sample/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Sample/rr
      -- 
    cp_elements(1170) <= cp_elements(1166);
    rr_4452_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1170), ack => unary_844_inst_req_0); -- 
    -- CP-element group 1171 transition  input  bypass 
    -- predecessors 1170 
    -- successors 1167 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Sample/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Sample/ra
      -- 
    ra_4453_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => unary_844_inst_ack_0, ack => cp_elements(1171)); -- 
    -- CP-element group 1172 transition  output  bypass 
    -- predecessors 1168 
    -- successors 1173 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Update/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Update/cr
      -- 
    cp_elements(1172) <= cp_elements(1168);
    cr_4457_symbol_link_to_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => cp_elements(1172), ack => unary_844_inst_req_1); -- 
    -- CP-element group 1173 transition  input  bypass 
    -- predecessors 1172 
    -- successors 1169 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Update/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/unary_844_Update/ca
      -- 
    ca_4458_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => unary_844_inst_ack_1, ack => cp_elements(1173)); -- 
    -- CP-element group 1174 fork  transition  bypass 
    -- predecessors 1127 
    -- successors 1175 
    -- marked successors 902 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/ring_reenable_memory_space_2
      -- 
    cp_elements(1174) <= cp_elements(1127);
    -- CP-element group 1175 join  transition  bypass 
    -- predecessors 99 164 877 904 936 968 1096 1128 1143 791 1000 1032 834 705 748 1064 1154 1164 1174 359 23 34 576 619 662 424 229 294 
    -- successors 4 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398_loop_body/$exit
      -- 
    cpelement_group_1175 : Block -- 
      signal predecessors: BooleanArray(27 downto 0);
      -- 
    begin -- 
      predecessors(0) <= cp_elements(99);
      predecessors(1) <= cp_elements(164);
      predecessors(2) <= cp_elements(877);
      predecessors(3) <= cp_elements(904);
      predecessors(4) <= cp_elements(936);
      predecessors(5) <= cp_elements(968);
      predecessors(6) <= cp_elements(1096);
      predecessors(7) <= cp_elements(1128);
      predecessors(8) <= cp_elements(1143);
      predecessors(9) <= cp_elements(791);
      predecessors(10) <= cp_elements(1000);
      predecessors(11) <= cp_elements(1032);
      predecessors(12) <= cp_elements(834);
      predecessors(13) <= cp_elements(705);
      predecessors(14) <= cp_elements(748);
      predecessors(15) <= cp_elements(1064);
      predecessors(16) <= cp_elements(1154);
      predecessors(17) <= cp_elements(1164);
      predecessors(18) <= cp_elements(1174);
      predecessors(19) <= cp_elements(359);
      predecessors(20) <= cp_elements(23);
      predecessors(21) <= cp_elements(34);
      predecessors(22) <= cp_elements(576);
      predecessors(23) <= cp_elements(619);
      predecessors(24) <= cp_elements(662);
      predecessors(25) <= cp_elements(424);
      predecessors(26) <= cp_elements(229);
      predecessors(27) <= cp_elements(294);
      jNoI: join -- 
        generic map(place_capacity => 16,
        bypass => true,
        name => " cp_elements(1175)_join")
        port map( -- 
          preds => predecessors,
          symbol_out => cp_elements(1175),
          clk => clk,
          reset => reset); -- 
      -- 
    end Block;
    -- CP-element group 1176 transition  bypass 
    -- predecessors 3 
    -- successors 1177 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_exit/$entry
      -- 
    cp_elements(1176) <= cp_elements(3);
    -- CP-element group 1177 transition  input  bypass 
    -- predecessors 1176 
    -- successors 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_exit/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_exit/ack
      -- 
    ack_4463_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_398_branch_ack_0, ack => cp_elements(1177)); -- 
    -- CP-element group 1178 transition  bypass 
    -- predecessors 3 
    -- successors 1179 
    -- members (1) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_taken/$entry
      -- 
    cp_elements(1178) <= cp_elements(3);
    -- CP-element group 1179 transition  input  bypass 
    -- predecessors 1178 
    -- successors 
    -- members (2) 
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_taken/$exit
      -- 	branch_block_stmt_389/do_while_stmt_398/loop_taken/ack
      -- 
    ack_4467_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_398_branch_ack_1, ack => cp_elements(1179)); -- 
    -- CP-element group 1180 transition  place  bypass 
    -- predecessors 1 
    -- successors 
    -- members (21) 
      -- 	$exit
      -- 	branch_block_stmt_389/$exit
      -- 	branch_block_stmt_389/branch_block_stmt_389__exit__
      -- 	branch_block_stmt_389/do_while_stmt_398__exit__
      -- 	branch_block_stmt_389/bb_1_xx_x_crit_edge
      -- 	branch_block_stmt_389/merge_stmt_846__exit__
      -- 	branch_block_stmt_389/return__
      -- 	branch_block_stmt_389/merge_stmt_848__exit__
      -- 	branch_block_stmt_389/do_while_stmt_398/$exit
      -- 	branch_block_stmt_389/bb_1_xx_x_crit_edge_PhiReq/$entry
      -- 	branch_block_stmt_389/bb_1_xx_x_crit_edge_PhiReq/$exit
      -- 	branch_block_stmt_389/merge_stmt_846_PhiReqMerge
      -- 	branch_block_stmt_389/merge_stmt_846_PhiAck/$entry
      -- 	branch_block_stmt_389/merge_stmt_846_PhiAck/$exit
      -- 	branch_block_stmt_389/merge_stmt_846_PhiAck/dummy
      -- 	branch_block_stmt_389/return___PhiReq/$entry
      -- 	branch_block_stmt_389/return___PhiReq/$exit
      -- 	branch_block_stmt_389/merge_stmt_848_PhiReqMerge
      -- 	branch_block_stmt_389/merge_stmt_848_PhiAck/$entry
      -- 	branch_block_stmt_389/merge_stmt_848_PhiAck/$exit
      -- 	branch_block_stmt_389/merge_stmt_848_PhiAck/dummy
      -- 
    cp_elements(1180) <= cp_elements(1);
    -- CP-element group 1181 transition  place  input  bypass 
    -- predecessors 0 
    -- successors 6 
    -- members (6) 
      -- 	branch_block_stmt_389/merge_stmt_391__exit__
      -- 	branch_block_stmt_389/do_while_stmt_398__entry__
      -- 	branch_block_stmt_389/do_while_stmt_398/$entry
      -- 	branch_block_stmt_389/do_while_stmt_398/do_while_stmt_398__entry__
      -- 	branch_block_stmt_389/merge_stmt_391_PhiAck/$exit
      -- 	branch_block_stmt_389/merge_stmt_391_PhiAck/phi_stmt_392_ack
      -- 
    phi_stmt_392_ack_4483_symbol_link_from_dp: control_delay_element -- 
      generic map (delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_392_ack_0, ack => cp_elements(1181)); -- 
    do_while_stmt_398_terminator_4468: loop_terminator -- 
      generic map (max_iterations_in_flight =>16) 
      port map(loop_body_exit => cp_elements(4),loop_continue => cp_elements(1179),loop_terminate => cp_elements(1177),loop_back => cp_elements(2),loop_exit => cp_elements(1),clk => clk, reset => reset); -- 
    phi_stmt_400_phi_seq_1336_block : block -- 
      signal reqs, selects : BooleanArray(0 to 1);
      signal enables : BooleanArray(0 to 0); -- 
    begin -- 
      selects(0)  <= cp_elements(10);
      cp_elements(8) <= reqs(0);
      selects(1)  <= cp_elements(13);
      cp_elements(11) <= reqs(1);
      enables(0)  <= cp_elements(17);
      phi_stmt_400_phi_seq_1336 : phi_sequencer -- 
        generic map (place_capacity => 16, nreqs => 2, nenables => 1, name => "phi_stmt_400_phi_seq_1336") 
        port map (selects => selects, reqs => reqs, enables => enables, ack => cp_elements(16), done => cp_elements(15), clk => clk, reset => reset);
        -- 
    end block;
    entry_tmerge_1322_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= cp_elements(5);
        preds(1)  <= cp_elements(6);
        entry_tmerge_1322 : transition_merge -- 
          port map (preds => preds, symbol_out => cp_elements(7));
          -- 
    end block;
    phi_stmt_400_req_merger_1337_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= cp_elements(9);
        preds(1)  <= cp_elements(12);
        phi_stmt_400_req_merger_1337 : transition_merge -- 
          port map (preds => preds, symbol_out => cp_elements(14));
          -- 
    end block;
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal array_obj_ref_420_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_420_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_420_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_420_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_425_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_425_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_425_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_425_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_430_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_430_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_430_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_430_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_441_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_441_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_441_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_441_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_446_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_446_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_446_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_446_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_451_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_451_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_451_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_451_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_462_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_462_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_462_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_462_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_467_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_467_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_467_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_467_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_472_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_472_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_472_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_472_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_483_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_483_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_483_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_483_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_488_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_488_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_488_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_488_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_493_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_493_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_493_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_493_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_504_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_504_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_504_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_504_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_509_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_509_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_509_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_509_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_514_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_514_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_514_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_514_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_525_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_525_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_525_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_525_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_530_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_530_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_530_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_530_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_535_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_535_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_535_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_535_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_546_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_546_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_546_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_546_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_551_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_551_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_551_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_551_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_556_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_556_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_556_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_556_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_561_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_561_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_561_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_561_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_566_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_566_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_566_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_566_root_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_571_final_offset : std_logic_vector(6 downto 0);
    signal array_obj_ref_571_offset_scale_factor_0 : std_logic_vector(6 downto 0);
    signal array_obj_ref_571_resized_base_address : std_logic_vector(6 downto 0);
    signal array_obj_ref_571_root_address : std_logic_vector(6 downto 0);
    signal exitcond1_841 : std_logic_vector(0 downto 0);
    signal iNsTr_10_612 : std_logic_vector(31 downto 0);
    signal iNsTr_11_616 : std_logic_vector(31 downto 0);
    signal iNsTr_12_620 : std_logic_vector(31 downto 0);
    signal iNsTr_13_625 : std_logic_vector(31 downto 0);
    signal iNsTr_14_629 : std_logic_vector(31 downto 0);
    signal iNsTr_15_633 : std_logic_vector(31 downto 0);
    signal iNsTr_16_638 : std_logic_vector(31 downto 0);
    signal iNsTr_17_642 : std_logic_vector(31 downto 0);
    signal iNsTr_18_646 : std_logic_vector(31 downto 0);
    signal iNsTr_19_651 : std_logic_vector(31 downto 0);
    signal iNsTr_20_655 : std_logic_vector(31 downto 0);
    signal iNsTr_21_659 : std_logic_vector(31 downto 0);
    signal iNsTr_22_664 : std_logic_vector(31 downto 0);
    signal iNsTr_23_668 : std_logic_vector(31 downto 0);
    signal iNsTr_24_672 : std_logic_vector(31 downto 0);
    signal iNsTr_25_677 : std_logic_vector(31 downto 0);
    signal iNsTr_2_577 : std_logic_vector(31 downto 0);
    signal iNsTr_3_581 : std_logic_vector(31 downto 0);
    signal iNsTr_4_586 : std_logic_vector(31 downto 0);
    signal iNsTr_5_590 : std_logic_vector(31 downto 0);
    signal iNsTr_6_594 : std_logic_vector(31 downto 0);
    signal iNsTr_7_599 : std_logic_vector(31 downto 0);
    signal iNsTr_8_603 : std_logic_vector(31 downto 0);
    signal iNsTr_9_607 : std_logic_vector(31 downto 0);
    signal indvar_400 : std_logic_vector(31 downto 0);
    signal indvar_at_entry_392 : std_logic_vector(31 downto 0);
    signal indvarx_xnext_835 : std_logic_vector(31 downto 0);
    signal ptr_deref_576_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_576_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_576_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_576_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_576_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_580_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_580_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_580_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_580_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_580_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_589_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_589_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_589_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_589_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_589_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_593_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_593_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_593_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_593_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_593_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_602_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_602_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_602_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_602_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_602_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_606_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_606_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_606_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_606_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_606_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_615_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_615_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_615_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_615_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_615_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_619_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_619_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_619_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_619_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_619_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_628_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_628_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_628_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_628_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_628_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_632_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_632_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_632_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_632_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_632_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_641_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_641_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_641_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_641_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_641_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_645_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_645_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_645_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_645_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_645_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_654_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_654_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_654_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_654_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_654_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_658_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_658_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_658_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_658_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_658_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_667_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_667_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_667_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_667_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_667_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_671_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_671_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_671_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_671_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_671_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_694_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_694_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_694_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_694_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_694_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_694_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_713_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_713_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_713_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_713_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_713_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_713_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_732_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_732_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_732_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_732_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_732_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_732_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_751_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_751_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_751_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_751_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_751_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_751_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_770_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_770_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_770_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_770_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_770_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_770_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_789_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_789_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_789_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_789_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_789_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_789_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_808_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_808_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_808_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_808_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_808_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_808_word_offset_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_827_data_0 : std_logic_vector(31 downto 0);
    signal ptr_deref_827_resized_base_address : std_logic_vector(6 downto 0);
    signal ptr_deref_827_root_address : std_logic_vector(6 downto 0);
    signal ptr_deref_827_wire : std_logic_vector(31 downto 0);
    signal ptr_deref_827_word_address_0 : std_logic_vector(6 downto 0);
    signal ptr_deref_827_word_offset_0 : std_logic_vector(6 downto 0);
    signal scevgep10_532 : std_logic_vector(31 downto 0);
    signal scevgep11_527 : std_logic_vector(31 downto 0);
    signal scevgep11_686_718 : std_logic_vector(31 downto 0);
    signal scevgep11_686_delayed_1_721 : std_logic_vector(31 downto 0);
    signal scevgep11_686_delayed_2_724 : std_logic_vector(31 downto 0);
    signal scevgep11_686_delayed_3_727 : std_logic_vector(31 downto 0);
    signal scevgep11_686_delayed_4_730 : std_logic_vector(31 downto 0);
    signal scevgep13_516 : std_logic_vector(31 downto 0);
    signal scevgep14_511 : std_logic_vector(31 downto 0);
    signal scevgep15_506 : std_logic_vector(31 downto 0);
    signal scevgep15_690_737 : std_logic_vector(31 downto 0);
    signal scevgep15_690_delayed_1_740 : std_logic_vector(31 downto 0);
    signal scevgep15_690_delayed_2_743 : std_logic_vector(31 downto 0);
    signal scevgep15_690_delayed_3_746 : std_logic_vector(31 downto 0);
    signal scevgep15_690_delayed_4_749 : std_logic_vector(31 downto 0);
    signal scevgep17_495 : std_logic_vector(31 downto 0);
    signal scevgep18_490 : std_logic_vector(31 downto 0);
    signal scevgep19_485 : std_logic_vector(31 downto 0);
    signal scevgep19_694_756 : std_logic_vector(31 downto 0);
    signal scevgep19_694_delayed_1_759 : std_logic_vector(31 downto 0);
    signal scevgep19_694_delayed_2_762 : std_logic_vector(31 downto 0);
    signal scevgep19_694_delayed_3_765 : std_logic_vector(31 downto 0);
    signal scevgep19_694_delayed_4_768 : std_logic_vector(31 downto 0);
    signal scevgep21_474 : std_logic_vector(31 downto 0);
    signal scevgep22_469 : std_logic_vector(31 downto 0);
    signal scevgep23_464 : std_logic_vector(31 downto 0);
    signal scevgep23_698_775 : std_logic_vector(31 downto 0);
    signal scevgep23_698_delayed_1_778 : std_logic_vector(31 downto 0);
    signal scevgep23_698_delayed_2_781 : std_logic_vector(31 downto 0);
    signal scevgep23_698_delayed_3_784 : std_logic_vector(31 downto 0);
    signal scevgep23_698_delayed_4_787 : std_logic_vector(31 downto 0);
    signal scevgep25_453 : std_logic_vector(31 downto 0);
    signal scevgep26_448 : std_logic_vector(31 downto 0);
    signal scevgep27_443 : std_logic_vector(31 downto 0);
    signal scevgep27_702_794 : std_logic_vector(31 downto 0);
    signal scevgep27_702_delayed_1_797 : std_logic_vector(31 downto 0);
    signal scevgep27_702_delayed_2_800 : std_logic_vector(31 downto 0);
    signal scevgep27_702_delayed_3_803 : std_logic_vector(31 downto 0);
    signal scevgep27_702_delayed_4_806 : std_logic_vector(31 downto 0);
    signal scevgep29_432 : std_logic_vector(31 downto 0);
    signal scevgep2_568 : std_logic_vector(31 downto 0);
    signal scevgep30_427 : std_logic_vector(31 downto 0);
    signal scevgep31_422 : std_logic_vector(31 downto 0);
    signal scevgep31_706_813 : std_logic_vector(31 downto 0);
    signal scevgep31_706_delayed_1_816 : std_logic_vector(31 downto 0);
    signal scevgep31_706_delayed_2_819 : std_logic_vector(31 downto 0);
    signal scevgep31_706_delayed_3_822 : std_logic_vector(31 downto 0);
    signal scevgep31_706_delayed_4_825 : std_logic_vector(31 downto 0);
    signal scevgep3_563 : std_logic_vector(31 downto 0);
    signal scevgep3_678_680 : std_logic_vector(31 downto 0);
    signal scevgep3_678_delayed_1_683 : std_logic_vector(31 downto 0);
    signal scevgep3_678_delayed_2_686 : std_logic_vector(31 downto 0);
    signal scevgep3_678_delayed_3_689 : std_logic_vector(31 downto 0);
    signal scevgep3_678_delayed_4_692 : std_logic_vector(31 downto 0);
    signal scevgep5_558 : std_logic_vector(31 downto 0);
    signal scevgep6_553 : std_logic_vector(31 downto 0);
    signal scevgep7_548 : std_logic_vector(31 downto 0);
    signal scevgep7_682_699 : std_logic_vector(31 downto 0);
    signal scevgep7_682_delayed_1_702 : std_logic_vector(31 downto 0);
    signal scevgep7_682_delayed_2_705 : std_logic_vector(31 downto 0);
    signal scevgep7_682_delayed_3_708 : std_logic_vector(31 downto 0);
    signal scevgep7_682_delayed_4_711 : std_logic_vector(31 downto 0);
    signal scevgep9_537 : std_logic_vector(31 downto 0);
    signal scevgep_573 : std_logic_vector(31 downto 0);
    signal simple_obj_ref_419_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_419_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_424_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_424_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_429_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_429_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_440_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_440_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_445_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_445_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_450_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_450_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_461_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_461_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_466_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_466_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_471_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_471_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_482_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_482_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_487_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_487_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_492_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_492_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_503_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_503_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_508_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_508_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_513_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_513_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_524_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_524_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_529_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_529_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_534_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_534_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_545_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_545_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_550_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_550_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_555_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_555_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_560_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_560_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_565_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_565_scaled : std_logic_vector(6 downto 0);
    signal simple_obj_ref_570_resized : std_logic_vector(6 downto 0);
    signal simple_obj_ref_570_scaled : std_logic_vector(6 downto 0);
    signal tmp13_438 : std_logic_vector(31 downto 0);
    signal tmp25_459 : std_logic_vector(31 downto 0);
    signal tmp2_411 : std_logic_vector(31 downto 0);
    signal tmp34_480 : std_logic_vector(31 downto 0);
    signal tmp38_501 : std_logic_vector(31 downto 0);
    signal tmp3_417 : std_logic_vector(31 downto 0);
    signal tmp42_522 : std_logic_vector(31 downto 0);
    signal tmp46_543 : std_logic_vector(31 downto 0);
    signal type_cast_396_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_403_wire : std_logic_vector(31 downto 0);
    signal type_cast_409_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_415_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_436_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_457_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_478_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_520_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_541_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_833_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_839_wire_constant : std_logic_vector(31 downto 0);
    signal unary_844_wire : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    array_obj_ref_420_offset_scale_factor_0 <= "0000001";
    array_obj_ref_420_resized_base_address <= "0000000";
    array_obj_ref_425_offset_scale_factor_0 <= "0000001";
    array_obj_ref_425_resized_base_address <= "0000000";
    array_obj_ref_430_offset_scale_factor_0 <= "0000001";
    array_obj_ref_430_resized_base_address <= "0000000";
    array_obj_ref_441_offset_scale_factor_0 <= "0000001";
    array_obj_ref_441_resized_base_address <= "0000000";
    array_obj_ref_446_offset_scale_factor_0 <= "0000001";
    array_obj_ref_446_resized_base_address <= "0000000";
    array_obj_ref_451_offset_scale_factor_0 <= "0000001";
    array_obj_ref_451_resized_base_address <= "0000000";
    array_obj_ref_462_offset_scale_factor_0 <= "0000001";
    array_obj_ref_462_resized_base_address <= "0000000";
    array_obj_ref_467_offset_scale_factor_0 <= "0000001";
    array_obj_ref_467_resized_base_address <= "0000000";
    array_obj_ref_472_offset_scale_factor_0 <= "0000001";
    array_obj_ref_472_resized_base_address <= "0000000";
    array_obj_ref_483_offset_scale_factor_0 <= "0000001";
    array_obj_ref_483_resized_base_address <= "0000000";
    array_obj_ref_488_offset_scale_factor_0 <= "0000001";
    array_obj_ref_488_resized_base_address <= "0000000";
    array_obj_ref_493_offset_scale_factor_0 <= "0000001";
    array_obj_ref_493_resized_base_address <= "0000000";
    array_obj_ref_504_offset_scale_factor_0 <= "0000001";
    array_obj_ref_504_resized_base_address <= "0000000";
    array_obj_ref_509_offset_scale_factor_0 <= "0000001";
    array_obj_ref_509_resized_base_address <= "0000000";
    array_obj_ref_514_offset_scale_factor_0 <= "0000001";
    array_obj_ref_514_resized_base_address <= "0000000";
    array_obj_ref_525_offset_scale_factor_0 <= "0000001";
    array_obj_ref_525_resized_base_address <= "0000000";
    array_obj_ref_530_offset_scale_factor_0 <= "0000001";
    array_obj_ref_530_resized_base_address <= "0000000";
    array_obj_ref_535_offset_scale_factor_0 <= "0000001";
    array_obj_ref_535_resized_base_address <= "0000000";
    array_obj_ref_546_offset_scale_factor_0 <= "0000001";
    array_obj_ref_546_resized_base_address <= "0000000";
    array_obj_ref_551_offset_scale_factor_0 <= "0000001";
    array_obj_ref_551_resized_base_address <= "0000000";
    array_obj_ref_556_offset_scale_factor_0 <= "0000001";
    array_obj_ref_556_resized_base_address <= "0000000";
    array_obj_ref_561_offset_scale_factor_0 <= "0000001";
    array_obj_ref_561_resized_base_address <= "0000000";
    array_obj_ref_566_offset_scale_factor_0 <= "0000001";
    array_obj_ref_566_resized_base_address <= "0000000";
    array_obj_ref_571_offset_scale_factor_0 <= "0000001";
    array_obj_ref_571_resized_base_address <= "0000000";
    ptr_deref_576_word_offset_0 <= "0000000";
    ptr_deref_580_word_offset_0 <= "0000000";
    ptr_deref_589_word_offset_0 <= "0000000";
    ptr_deref_593_word_offset_0 <= "0000000";
    ptr_deref_602_word_offset_0 <= "0000000";
    ptr_deref_606_word_offset_0 <= "0000000";
    ptr_deref_615_word_offset_0 <= "0000000";
    ptr_deref_619_word_offset_0 <= "0000000";
    ptr_deref_628_word_offset_0 <= "0000000";
    ptr_deref_632_word_offset_0 <= "0000000";
    ptr_deref_641_word_offset_0 <= "0000000";
    ptr_deref_645_word_offset_0 <= "0000000";
    ptr_deref_654_word_offset_0 <= "0000000";
    ptr_deref_658_word_offset_0 <= "0000000";
    ptr_deref_667_word_offset_0 <= "0000000";
    ptr_deref_671_word_offset_0 <= "0000000";
    ptr_deref_694_word_offset_0 <= "0000000";
    ptr_deref_713_word_offset_0 <= "0000000";
    ptr_deref_732_word_offset_0 <= "0000000";
    ptr_deref_751_word_offset_0 <= "0000000";
    ptr_deref_770_word_offset_0 <= "0000000";
    ptr_deref_789_word_offset_0 <= "0000000";
    ptr_deref_808_word_offset_0 <= "0000000";
    ptr_deref_827_word_offset_0 <= "0000000";
    type_cast_396_wire_constant <= "00000000000000000000000000000000";
    type_cast_409_wire_constant <= "00000000000000000000000000001000";
    type_cast_415_wire_constant <= "00000000000000000000000000000111";
    type_cast_436_wire_constant <= "00000000000000000000000000000110";
    type_cast_457_wire_constant <= "00000000000000000000000000000101";
    type_cast_478_wire_constant <= "00000000000000000000000000000100";
    type_cast_499_wire_constant <= "00000000000000000000000000000011";
    type_cast_520_wire_constant <= "00000000000000000000000000000010";
    type_cast_541_wire_constant <= "00000000000000000000000000000001";
    type_cast_833_wire_constant <= "00000000000000000000000000000001";
    type_cast_839_wire_constant <= "00000000000000000000000000001000";
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_392_req_0," req0 phi_stmt_392");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_392_ack_0," ack0 phi_stmt_392");
    phi_stmt_392: Block -- phi operator 
      signal idata: std_logic_vector(31 downto 0);
      signal req: BooleanArray(0 downto 0);
      --
    begin -- 
      idata <= type_cast_396_wire_constant;
      req(0) <= phi_stmt_392_req_0;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 1,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_392_ack_0,
          idata => idata,
          odata => indvar_at_entry_392,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_392
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_400_req_0," req0 phi_stmt_400");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_400_req_1," req1 phi_stmt_400");
    LogCPEvent(clk, reset, global_clock_cycle_count,phi_stmt_400_ack_0," ack0 phi_stmt_400");
    phi_stmt_400: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_403_wire & indvar_at_entry_392;
      req <= phi_stmt_400_req_0 & phi_stmt_400_req_1;
      phi: PhiBase -- 
        generic map( -- 
          num_reqs => 2,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_400_ack_0,
          idata => idata,
          odata => indvar_400,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_400
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_421_final_reg_req_0,addr_of_421_final_reg_ack_0,sl_one,"addr_of_421_final_reg ",false,array_obj_ref_420_root_address,
    false,scevgep31_422);
    register_block_0 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_421_final_reg_req_0;
      addr_of_421_final_reg_ack_0 <= ack; 
      addr_of_421_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_420_root_address, dout => scevgep31_422, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_426_final_reg_req_0,addr_of_426_final_reg_ack_0,sl_one,"addr_of_426_final_reg ",false,array_obj_ref_425_root_address,
    false,scevgep30_427);
    register_block_1 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_426_final_reg_req_0;
      addr_of_426_final_reg_ack_0 <= ack; 
      addr_of_426_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_425_root_address, dout => scevgep30_427, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_431_final_reg_req_0,addr_of_431_final_reg_ack_0,sl_one,"addr_of_431_final_reg ",false,array_obj_ref_430_root_address,
    false,scevgep29_432);
    register_block_2 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_431_final_reg_req_0;
      addr_of_431_final_reg_ack_0 <= ack; 
      addr_of_431_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_430_root_address, dout => scevgep29_432, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_442_final_reg_req_0,addr_of_442_final_reg_ack_0,sl_one,"addr_of_442_final_reg ",false,array_obj_ref_441_root_address,
    false,scevgep27_443);
    register_block_3 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_442_final_reg_req_0;
      addr_of_442_final_reg_ack_0 <= ack; 
      addr_of_442_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_441_root_address, dout => scevgep27_443, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_447_final_reg_req_0,addr_of_447_final_reg_ack_0,sl_one,"addr_of_447_final_reg ",false,array_obj_ref_446_root_address,
    false,scevgep26_448);
    register_block_4 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_447_final_reg_req_0;
      addr_of_447_final_reg_ack_0 <= ack; 
      addr_of_447_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_446_root_address, dout => scevgep26_448, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_452_final_reg_req_0,addr_of_452_final_reg_ack_0,sl_one,"addr_of_452_final_reg ",false,array_obj_ref_451_root_address,
    false,scevgep25_453);
    register_block_5 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_452_final_reg_req_0;
      addr_of_452_final_reg_ack_0 <= ack; 
      addr_of_452_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_451_root_address, dout => scevgep25_453, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_463_final_reg_req_0,addr_of_463_final_reg_ack_0,sl_one,"addr_of_463_final_reg ",false,array_obj_ref_462_root_address,
    false,scevgep23_464);
    register_block_6 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_463_final_reg_req_0;
      addr_of_463_final_reg_ack_0 <= ack; 
      addr_of_463_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_462_root_address, dout => scevgep23_464, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_468_final_reg_req_0,addr_of_468_final_reg_ack_0,sl_one,"addr_of_468_final_reg ",false,array_obj_ref_467_root_address,
    false,scevgep22_469);
    register_block_7 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_468_final_reg_req_0;
      addr_of_468_final_reg_ack_0 <= ack; 
      addr_of_468_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_467_root_address, dout => scevgep22_469, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_473_final_reg_req_0,addr_of_473_final_reg_ack_0,sl_one,"addr_of_473_final_reg ",false,array_obj_ref_472_root_address,
    false,scevgep21_474);
    register_block_8 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_473_final_reg_req_0;
      addr_of_473_final_reg_ack_0 <= ack; 
      addr_of_473_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_472_root_address, dout => scevgep21_474, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_484_final_reg_req_0,addr_of_484_final_reg_ack_0,sl_one,"addr_of_484_final_reg ",false,array_obj_ref_483_root_address,
    false,scevgep19_485);
    register_block_9 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_484_final_reg_req_0;
      addr_of_484_final_reg_ack_0 <= ack; 
      addr_of_484_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_483_root_address, dout => scevgep19_485, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_489_final_reg_req_0,addr_of_489_final_reg_ack_0,sl_one,"addr_of_489_final_reg ",false,array_obj_ref_488_root_address,
    false,scevgep18_490);
    register_block_10 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_489_final_reg_req_0;
      addr_of_489_final_reg_ack_0 <= ack; 
      addr_of_489_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_488_root_address, dout => scevgep18_490, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_494_final_reg_req_0,addr_of_494_final_reg_ack_0,sl_one,"addr_of_494_final_reg ",false,array_obj_ref_493_root_address,
    false,scevgep17_495);
    register_block_11 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_494_final_reg_req_0;
      addr_of_494_final_reg_ack_0 <= ack; 
      addr_of_494_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_493_root_address, dout => scevgep17_495, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_505_final_reg_req_0,addr_of_505_final_reg_ack_0,sl_one,"addr_of_505_final_reg ",false,array_obj_ref_504_root_address,
    false,scevgep15_506);
    register_block_12 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_505_final_reg_req_0;
      addr_of_505_final_reg_ack_0 <= ack; 
      addr_of_505_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_504_root_address, dout => scevgep15_506, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_510_final_reg_req_0,addr_of_510_final_reg_ack_0,sl_one,"addr_of_510_final_reg ",false,array_obj_ref_509_root_address,
    false,scevgep14_511);
    register_block_13 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_510_final_reg_req_0;
      addr_of_510_final_reg_ack_0 <= ack; 
      addr_of_510_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_509_root_address, dout => scevgep14_511, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_515_final_reg_req_0,addr_of_515_final_reg_ack_0,sl_one,"addr_of_515_final_reg ",false,array_obj_ref_514_root_address,
    false,scevgep13_516);
    register_block_14 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_515_final_reg_req_0;
      addr_of_515_final_reg_ack_0 <= ack; 
      addr_of_515_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_514_root_address, dout => scevgep13_516, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_526_final_reg_req_0,addr_of_526_final_reg_ack_0,sl_one,"addr_of_526_final_reg ",false,array_obj_ref_525_root_address,
    false,scevgep11_527);
    register_block_15 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_526_final_reg_req_0;
      addr_of_526_final_reg_ack_0 <= ack; 
      addr_of_526_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_525_root_address, dout => scevgep11_527, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_531_final_reg_req_0,addr_of_531_final_reg_ack_0,sl_one,"addr_of_531_final_reg ",false,array_obj_ref_530_root_address,
    false,scevgep10_532);
    register_block_16 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_531_final_reg_req_0;
      addr_of_531_final_reg_ack_0 <= ack; 
      addr_of_531_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_530_root_address, dout => scevgep10_532, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_536_final_reg_req_0,addr_of_536_final_reg_ack_0,sl_one,"addr_of_536_final_reg ",false,array_obj_ref_535_root_address,
    false,scevgep9_537);
    register_block_17 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_536_final_reg_req_0;
      addr_of_536_final_reg_ack_0 <= ack; 
      addr_of_536_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_535_root_address, dout => scevgep9_537, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_547_final_reg_req_0,addr_of_547_final_reg_ack_0,sl_one,"addr_of_547_final_reg ",false,array_obj_ref_546_root_address,
    false,scevgep7_548);
    register_block_18 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_547_final_reg_req_0;
      addr_of_547_final_reg_ack_0 <= ack; 
      addr_of_547_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_546_root_address, dout => scevgep7_548, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_552_final_reg_req_0,addr_of_552_final_reg_ack_0,sl_one,"addr_of_552_final_reg ",false,array_obj_ref_551_root_address,
    false,scevgep6_553);
    register_block_19 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_552_final_reg_req_0;
      addr_of_552_final_reg_ack_0 <= ack; 
      addr_of_552_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_551_root_address, dout => scevgep6_553, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_557_final_reg_req_0,addr_of_557_final_reg_ack_0,sl_one,"addr_of_557_final_reg ",false,array_obj_ref_556_root_address,
    false,scevgep5_558);
    register_block_20 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_557_final_reg_req_0;
      addr_of_557_final_reg_ack_0 <= ack; 
      addr_of_557_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_556_root_address, dout => scevgep5_558, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_562_final_reg_req_0,addr_of_562_final_reg_ack_0,sl_one,"addr_of_562_final_reg ",false,array_obj_ref_561_root_address,
    false,scevgep3_563);
    register_block_21 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_562_final_reg_req_0;
      addr_of_562_final_reg_ack_0 <= ack; 
      addr_of_562_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_561_root_address, dout => scevgep3_563, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_567_final_reg_req_0,addr_of_567_final_reg_ack_0,sl_one,"addr_of_567_final_reg ",false,array_obj_ref_566_root_address,
    false,scevgep2_568);
    register_block_22 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_567_final_reg_req_0;
      addr_of_567_final_reg_ack_0 <= ack; 
      addr_of_567_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_566_root_address, dout => scevgep2_568, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,addr_of_572_final_reg_req_0,addr_of_572_final_reg_ack_0,sl_one,"addr_of_572_final_reg ",false,array_obj_ref_571_root_address,
    false,scevgep_573);
    register_block_23 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= addr_of_572_final_reg_req_0;
      addr_of_572_final_reg_ack_0 <= ack; 
      addr_of_572_final_reg: RegisterBase --
        generic map(in_data_width => 7,out_data_width => 32) 
        port map( din => array_obj_ref_571_root_address, dout => scevgep_573, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_678_inst_req_0,simple_obj_ref_678_inst_ack_0,sl_one,"simple_obj_ref_678_inst ",false,scevgep3_563,
    false,scevgep3_678_680);
    register_block_24 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_678_inst_req_0;
      simple_obj_ref_678_inst_ack_0 <= ack; 
      simple_obj_ref_678_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep3_563, dout => scevgep3_678_680, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_681_inst_req_0,simple_obj_ref_681_inst_ack_0,sl_one,"simple_obj_ref_681_inst ",false,scevgep3_678_680,
    false,scevgep3_678_delayed_1_683);
    register_block_25 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_681_inst_req_0;
      simple_obj_ref_681_inst_ack_0 <= ack; 
      simple_obj_ref_681_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep3_678_680, dout => scevgep3_678_delayed_1_683, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_684_inst_req_0,simple_obj_ref_684_inst_ack_0,sl_one,"simple_obj_ref_684_inst ",false,scevgep3_678_delayed_1_683,
    false,scevgep3_678_delayed_2_686);
    register_block_26 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_684_inst_req_0;
      simple_obj_ref_684_inst_ack_0 <= ack; 
      simple_obj_ref_684_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep3_678_delayed_1_683, dout => scevgep3_678_delayed_2_686, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_687_inst_req_0,simple_obj_ref_687_inst_ack_0,sl_one,"simple_obj_ref_687_inst ",false,scevgep3_678_delayed_2_686,
    false,scevgep3_678_delayed_3_689);
    register_block_27 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_687_inst_req_0;
      simple_obj_ref_687_inst_ack_0 <= ack; 
      simple_obj_ref_687_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep3_678_delayed_2_686, dout => scevgep3_678_delayed_3_689, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_690_inst_req_0,simple_obj_ref_690_inst_ack_0,sl_one,"simple_obj_ref_690_inst ",false,scevgep3_678_delayed_3_689,
    false,scevgep3_678_delayed_4_692);
    register_block_28 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_690_inst_req_0;
      simple_obj_ref_690_inst_ack_0 <= ack; 
      simple_obj_ref_690_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep3_678_delayed_3_689, dout => scevgep3_678_delayed_4_692, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_697_inst_req_0,simple_obj_ref_697_inst_ack_0,sl_one,"simple_obj_ref_697_inst ",false,scevgep7_548,
    false,scevgep7_682_699);
    register_block_29 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_697_inst_req_0;
      simple_obj_ref_697_inst_ack_0 <= ack; 
      simple_obj_ref_697_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep7_548, dout => scevgep7_682_699, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_700_inst_req_0,simple_obj_ref_700_inst_ack_0,sl_one,"simple_obj_ref_700_inst ",false,scevgep7_682_699,
    false,scevgep7_682_delayed_1_702);
    register_block_30 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_700_inst_req_0;
      simple_obj_ref_700_inst_ack_0 <= ack; 
      simple_obj_ref_700_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep7_682_699, dout => scevgep7_682_delayed_1_702, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_703_inst_req_0,simple_obj_ref_703_inst_ack_0,sl_one,"simple_obj_ref_703_inst ",false,scevgep7_682_delayed_1_702,
    false,scevgep7_682_delayed_2_705);
    register_block_31 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_703_inst_req_0;
      simple_obj_ref_703_inst_ack_0 <= ack; 
      simple_obj_ref_703_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep7_682_delayed_1_702, dout => scevgep7_682_delayed_2_705, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_706_inst_req_0,simple_obj_ref_706_inst_ack_0,sl_one,"simple_obj_ref_706_inst ",false,scevgep7_682_delayed_2_705,
    false,scevgep7_682_delayed_3_708);
    register_block_32 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_706_inst_req_0;
      simple_obj_ref_706_inst_ack_0 <= ack; 
      simple_obj_ref_706_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep7_682_delayed_2_705, dout => scevgep7_682_delayed_3_708, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_709_inst_req_0,simple_obj_ref_709_inst_ack_0,sl_one,"simple_obj_ref_709_inst ",false,scevgep7_682_delayed_3_708,
    false,scevgep7_682_delayed_4_711);
    register_block_33 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_709_inst_req_0;
      simple_obj_ref_709_inst_ack_0 <= ack; 
      simple_obj_ref_709_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep7_682_delayed_3_708, dout => scevgep7_682_delayed_4_711, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_716_inst_req_0,simple_obj_ref_716_inst_ack_0,sl_one,"simple_obj_ref_716_inst ",false,scevgep11_527,
    false,scevgep11_686_718);
    register_block_34 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_716_inst_req_0;
      simple_obj_ref_716_inst_ack_0 <= ack; 
      simple_obj_ref_716_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep11_527, dout => scevgep11_686_718, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_719_inst_req_0,simple_obj_ref_719_inst_ack_0,sl_one,"simple_obj_ref_719_inst ",false,scevgep11_686_718,
    false,scevgep11_686_delayed_1_721);
    register_block_35 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_719_inst_req_0;
      simple_obj_ref_719_inst_ack_0 <= ack; 
      simple_obj_ref_719_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep11_686_718, dout => scevgep11_686_delayed_1_721, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_722_inst_req_0,simple_obj_ref_722_inst_ack_0,sl_one,"simple_obj_ref_722_inst ",false,scevgep11_686_delayed_1_721,
    false,scevgep11_686_delayed_2_724);
    register_block_36 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_722_inst_req_0;
      simple_obj_ref_722_inst_ack_0 <= ack; 
      simple_obj_ref_722_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep11_686_delayed_1_721, dout => scevgep11_686_delayed_2_724, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_725_inst_req_0,simple_obj_ref_725_inst_ack_0,sl_one,"simple_obj_ref_725_inst ",false,scevgep11_686_delayed_2_724,
    false,scevgep11_686_delayed_3_727);
    register_block_37 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_725_inst_req_0;
      simple_obj_ref_725_inst_ack_0 <= ack; 
      simple_obj_ref_725_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep11_686_delayed_2_724, dout => scevgep11_686_delayed_3_727, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_728_inst_req_0,simple_obj_ref_728_inst_ack_0,sl_one,"simple_obj_ref_728_inst ",false,scevgep11_686_delayed_3_727,
    false,scevgep11_686_delayed_4_730);
    register_block_38 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_728_inst_req_0;
      simple_obj_ref_728_inst_ack_0 <= ack; 
      simple_obj_ref_728_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep11_686_delayed_3_727, dout => scevgep11_686_delayed_4_730, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_735_inst_req_0,simple_obj_ref_735_inst_ack_0,sl_one,"simple_obj_ref_735_inst ",false,scevgep15_506,
    false,scevgep15_690_737);
    register_block_39 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_735_inst_req_0;
      simple_obj_ref_735_inst_ack_0 <= ack; 
      simple_obj_ref_735_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep15_506, dout => scevgep15_690_737, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_738_inst_req_0,simple_obj_ref_738_inst_ack_0,sl_one,"simple_obj_ref_738_inst ",false,scevgep15_690_737,
    false,scevgep15_690_delayed_1_740);
    register_block_40 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_738_inst_req_0;
      simple_obj_ref_738_inst_ack_0 <= ack; 
      simple_obj_ref_738_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep15_690_737, dout => scevgep15_690_delayed_1_740, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_741_inst_req_0,simple_obj_ref_741_inst_ack_0,sl_one,"simple_obj_ref_741_inst ",false,scevgep15_690_delayed_1_740,
    false,scevgep15_690_delayed_2_743);
    register_block_41 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_741_inst_req_0;
      simple_obj_ref_741_inst_ack_0 <= ack; 
      simple_obj_ref_741_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep15_690_delayed_1_740, dout => scevgep15_690_delayed_2_743, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_744_inst_req_0,simple_obj_ref_744_inst_ack_0,sl_one,"simple_obj_ref_744_inst ",false,scevgep15_690_delayed_2_743,
    false,scevgep15_690_delayed_3_746);
    register_block_42 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_744_inst_req_0;
      simple_obj_ref_744_inst_ack_0 <= ack; 
      simple_obj_ref_744_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep15_690_delayed_2_743, dout => scevgep15_690_delayed_3_746, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_747_inst_req_0,simple_obj_ref_747_inst_ack_0,sl_one,"simple_obj_ref_747_inst ",false,scevgep15_690_delayed_3_746,
    false,scevgep15_690_delayed_4_749);
    register_block_43 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_747_inst_req_0;
      simple_obj_ref_747_inst_ack_0 <= ack; 
      simple_obj_ref_747_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep15_690_delayed_3_746, dout => scevgep15_690_delayed_4_749, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_754_inst_req_0,simple_obj_ref_754_inst_ack_0,sl_one,"simple_obj_ref_754_inst ",false,scevgep19_485,
    false,scevgep19_694_756);
    register_block_44 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_754_inst_req_0;
      simple_obj_ref_754_inst_ack_0 <= ack; 
      simple_obj_ref_754_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep19_485, dout => scevgep19_694_756, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_757_inst_req_0,simple_obj_ref_757_inst_ack_0,sl_one,"simple_obj_ref_757_inst ",false,scevgep19_694_756,
    false,scevgep19_694_delayed_1_759);
    register_block_45 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_757_inst_req_0;
      simple_obj_ref_757_inst_ack_0 <= ack; 
      simple_obj_ref_757_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep19_694_756, dout => scevgep19_694_delayed_1_759, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_760_inst_req_0,simple_obj_ref_760_inst_ack_0,sl_one,"simple_obj_ref_760_inst ",false,scevgep19_694_delayed_1_759,
    false,scevgep19_694_delayed_2_762);
    register_block_46 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_760_inst_req_0;
      simple_obj_ref_760_inst_ack_0 <= ack; 
      simple_obj_ref_760_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep19_694_delayed_1_759, dout => scevgep19_694_delayed_2_762, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_763_inst_req_0,simple_obj_ref_763_inst_ack_0,sl_one,"simple_obj_ref_763_inst ",false,scevgep19_694_delayed_2_762,
    false,scevgep19_694_delayed_3_765);
    register_block_47 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_763_inst_req_0;
      simple_obj_ref_763_inst_ack_0 <= ack; 
      simple_obj_ref_763_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep19_694_delayed_2_762, dout => scevgep19_694_delayed_3_765, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_766_inst_req_0,simple_obj_ref_766_inst_ack_0,sl_one,"simple_obj_ref_766_inst ",false,scevgep19_694_delayed_3_765,
    false,scevgep19_694_delayed_4_768);
    register_block_48 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_766_inst_req_0;
      simple_obj_ref_766_inst_ack_0 <= ack; 
      simple_obj_ref_766_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep19_694_delayed_3_765, dout => scevgep19_694_delayed_4_768, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_773_inst_req_0,simple_obj_ref_773_inst_ack_0,sl_one,"simple_obj_ref_773_inst ",false,scevgep23_464,
    false,scevgep23_698_775);
    register_block_49 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_773_inst_req_0;
      simple_obj_ref_773_inst_ack_0 <= ack; 
      simple_obj_ref_773_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep23_464, dout => scevgep23_698_775, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_776_inst_req_0,simple_obj_ref_776_inst_ack_0,sl_one,"simple_obj_ref_776_inst ",false,scevgep23_698_775,
    false,scevgep23_698_delayed_1_778);
    register_block_50 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_776_inst_req_0;
      simple_obj_ref_776_inst_ack_0 <= ack; 
      simple_obj_ref_776_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep23_698_775, dout => scevgep23_698_delayed_1_778, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_779_inst_req_0,simple_obj_ref_779_inst_ack_0,sl_one,"simple_obj_ref_779_inst ",false,scevgep23_698_delayed_1_778,
    false,scevgep23_698_delayed_2_781);
    register_block_51 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_779_inst_req_0;
      simple_obj_ref_779_inst_ack_0 <= ack; 
      simple_obj_ref_779_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep23_698_delayed_1_778, dout => scevgep23_698_delayed_2_781, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_782_inst_req_0,simple_obj_ref_782_inst_ack_0,sl_one,"simple_obj_ref_782_inst ",false,scevgep23_698_delayed_2_781,
    false,scevgep23_698_delayed_3_784);
    register_block_52 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_782_inst_req_0;
      simple_obj_ref_782_inst_ack_0 <= ack; 
      simple_obj_ref_782_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep23_698_delayed_2_781, dout => scevgep23_698_delayed_3_784, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_785_inst_req_0,simple_obj_ref_785_inst_ack_0,sl_one,"simple_obj_ref_785_inst ",false,scevgep23_698_delayed_3_784,
    false,scevgep23_698_delayed_4_787);
    register_block_53 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_785_inst_req_0;
      simple_obj_ref_785_inst_ack_0 <= ack; 
      simple_obj_ref_785_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep23_698_delayed_3_784, dout => scevgep23_698_delayed_4_787, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_792_inst_req_0,simple_obj_ref_792_inst_ack_0,sl_one,"simple_obj_ref_792_inst ",false,scevgep27_443,
    false,scevgep27_702_794);
    register_block_54 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_792_inst_req_0;
      simple_obj_ref_792_inst_ack_0 <= ack; 
      simple_obj_ref_792_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep27_443, dout => scevgep27_702_794, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_795_inst_req_0,simple_obj_ref_795_inst_ack_0,sl_one,"simple_obj_ref_795_inst ",false,scevgep27_702_794,
    false,scevgep27_702_delayed_1_797);
    register_block_55 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_795_inst_req_0;
      simple_obj_ref_795_inst_ack_0 <= ack; 
      simple_obj_ref_795_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep27_702_794, dout => scevgep27_702_delayed_1_797, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_798_inst_req_0,simple_obj_ref_798_inst_ack_0,sl_one,"simple_obj_ref_798_inst ",false,scevgep27_702_delayed_1_797,
    false,scevgep27_702_delayed_2_800);
    register_block_56 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_798_inst_req_0;
      simple_obj_ref_798_inst_ack_0 <= ack; 
      simple_obj_ref_798_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep27_702_delayed_1_797, dout => scevgep27_702_delayed_2_800, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_801_inst_req_0,simple_obj_ref_801_inst_ack_0,sl_one,"simple_obj_ref_801_inst ",false,scevgep27_702_delayed_2_800,
    false,scevgep27_702_delayed_3_803);
    register_block_57 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_801_inst_req_0;
      simple_obj_ref_801_inst_ack_0 <= ack; 
      simple_obj_ref_801_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep27_702_delayed_2_800, dout => scevgep27_702_delayed_3_803, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_804_inst_req_0,simple_obj_ref_804_inst_ack_0,sl_one,"simple_obj_ref_804_inst ",false,scevgep27_702_delayed_3_803,
    false,scevgep27_702_delayed_4_806);
    register_block_58 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_804_inst_req_0;
      simple_obj_ref_804_inst_ack_0 <= ack; 
      simple_obj_ref_804_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep27_702_delayed_3_803, dout => scevgep27_702_delayed_4_806, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_811_inst_req_0,simple_obj_ref_811_inst_ack_0,sl_one,"simple_obj_ref_811_inst ",false,scevgep31_422,
    false,scevgep31_706_813);
    register_block_59 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_811_inst_req_0;
      simple_obj_ref_811_inst_ack_0 <= ack; 
      simple_obj_ref_811_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep31_422, dout => scevgep31_706_813, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_814_inst_req_0,simple_obj_ref_814_inst_ack_0,sl_one,"simple_obj_ref_814_inst ",false,scevgep31_706_813,
    false,scevgep31_706_delayed_1_816);
    register_block_60 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_814_inst_req_0;
      simple_obj_ref_814_inst_ack_0 <= ack; 
      simple_obj_ref_814_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep31_706_813, dout => scevgep31_706_delayed_1_816, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_817_inst_req_0,simple_obj_ref_817_inst_ack_0,sl_one,"simple_obj_ref_817_inst ",false,scevgep31_706_delayed_1_816,
    false,scevgep31_706_delayed_2_819);
    register_block_61 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_817_inst_req_0;
      simple_obj_ref_817_inst_ack_0 <= ack; 
      simple_obj_ref_817_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep31_706_delayed_1_816, dout => scevgep31_706_delayed_2_819, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_820_inst_req_0,simple_obj_ref_820_inst_ack_0,sl_one,"simple_obj_ref_820_inst ",false,scevgep31_706_delayed_2_819,
    false,scevgep31_706_delayed_3_822);
    register_block_62 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_820_inst_req_0;
      simple_obj_ref_820_inst_ack_0 <= ack; 
      simple_obj_ref_820_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep31_706_delayed_2_819, dout => scevgep31_706_delayed_3_822, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,simple_obj_ref_823_inst_req_0,simple_obj_ref_823_inst_ack_0,sl_one,"simple_obj_ref_823_inst ",false,scevgep31_706_delayed_3_822,
    false,scevgep31_706_delayed_4_825);
    register_block_63 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= simple_obj_ref_823_inst_req_0;
      simple_obj_ref_823_inst_ack_0 <= ack; 
      simple_obj_ref_823_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => scevgep31_706_delayed_3_822, dout => scevgep31_706_delayed_4_825, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,type_cast_403_inst_req_0,type_cast_403_inst_ack_0,sl_one,"type_cast_403_inst ",false,indvarx_xnext_835,
    false,type_cast_403_wire);
    register_block_64 : block -- 
      signal req, ack: boolean; --
    begin -- 
      req <= type_cast_403_inst_req_0;
      type_cast_403_inst_ack_0 <= ack; 
      type_cast_403_inst: RegisterBase --
        generic map(in_data_width => 32,out_data_width => 32) 
        port map( din => indvarx_xnext_835, dout => type_cast_403_wire, req => req,  ack => ack,  clk => clk, reset => reset); -- 
      -- 
    end block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_420_index_0_rename_req_0,array_obj_ref_420_index_0_rename_ack_0,sl_one,"array_obj_ref_420_index_0_rename ",false,simple_obj_ref_419_resized,
    false,simple_obj_ref_419_scaled);
    array_obj_ref_420_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_420_index_0_rename_ack_0 <= array_obj_ref_420_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_419_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_419_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_420_index_0_resize_req_0,array_obj_ref_420_index_0_resize_ack_0,sl_one,"array_obj_ref_420_index_0_resize ",false,tmp3_417,
    false,simple_obj_ref_419_resized);
    array_obj_ref_420_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_420_index_0_resize_ack_0 <= array_obj_ref_420_index_0_resize_req_0;
      in_aggregated_sig <= tmp3_417;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_419_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_420_offset_inst_req_0,array_obj_ref_420_offset_inst_ack_0,sl_one,"array_obj_ref_420_offset_inst ",false,simple_obj_ref_419_scaled,
    false,array_obj_ref_420_final_offset);
    array_obj_ref_420_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_420_offset_inst_ack_0 <= array_obj_ref_420_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_419_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_420_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_420_root_address_inst_req_0,array_obj_ref_420_root_address_inst_ack_0,sl_one,"array_obj_ref_420_root_address_inst ",false,array_obj_ref_420_final_offset,
    false,array_obj_ref_420_root_address);
    array_obj_ref_420_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_420_root_address_inst_ack_0 <= array_obj_ref_420_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_420_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_420_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_425_index_0_rename_req_0,array_obj_ref_425_index_0_rename_ack_0,sl_one,"array_obj_ref_425_index_0_rename ",false,simple_obj_ref_424_resized,
    false,simple_obj_ref_424_scaled);
    array_obj_ref_425_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_425_index_0_rename_ack_0 <= array_obj_ref_425_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_424_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_424_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_425_index_0_resize_req_0,array_obj_ref_425_index_0_resize_ack_0,sl_one,"array_obj_ref_425_index_0_resize ",false,tmp3_417,
    false,simple_obj_ref_424_resized);
    array_obj_ref_425_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_425_index_0_resize_ack_0 <= array_obj_ref_425_index_0_resize_req_0;
      in_aggregated_sig <= tmp3_417;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_424_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_425_offset_inst_req_0,array_obj_ref_425_offset_inst_ack_0,sl_one,"array_obj_ref_425_offset_inst ",false,simple_obj_ref_424_scaled,
    false,array_obj_ref_425_final_offset);
    array_obj_ref_425_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_425_offset_inst_ack_0 <= array_obj_ref_425_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_424_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_425_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_425_root_address_inst_req_0,array_obj_ref_425_root_address_inst_ack_0,sl_one,"array_obj_ref_425_root_address_inst ",false,array_obj_ref_425_final_offset,
    false,array_obj_ref_425_root_address);
    array_obj_ref_425_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_425_root_address_inst_ack_0 <= array_obj_ref_425_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_425_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_425_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_430_index_0_rename_req_0,array_obj_ref_430_index_0_rename_ack_0,sl_one,"array_obj_ref_430_index_0_rename ",false,simple_obj_ref_429_resized,
    false,simple_obj_ref_429_scaled);
    array_obj_ref_430_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_430_index_0_rename_ack_0 <= array_obj_ref_430_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_429_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_429_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_430_index_0_resize_req_0,array_obj_ref_430_index_0_resize_ack_0,sl_one,"array_obj_ref_430_index_0_resize ",false,tmp3_417,
    false,simple_obj_ref_429_resized);
    array_obj_ref_430_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_430_index_0_resize_ack_0 <= array_obj_ref_430_index_0_resize_req_0;
      in_aggregated_sig <= tmp3_417;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_429_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_430_offset_inst_req_0,array_obj_ref_430_offset_inst_ack_0,sl_one,"array_obj_ref_430_offset_inst ",false,simple_obj_ref_429_scaled,
    false,array_obj_ref_430_final_offset);
    array_obj_ref_430_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_430_offset_inst_ack_0 <= array_obj_ref_430_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_429_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_430_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_430_root_address_inst_req_0,array_obj_ref_430_root_address_inst_ack_0,sl_one,"array_obj_ref_430_root_address_inst ",false,array_obj_ref_430_final_offset,
    false,array_obj_ref_430_root_address);
    array_obj_ref_430_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_430_root_address_inst_ack_0 <= array_obj_ref_430_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_430_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_430_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_441_index_0_rename_req_0,array_obj_ref_441_index_0_rename_ack_0,sl_one,"array_obj_ref_441_index_0_rename ",false,simple_obj_ref_440_resized,
    false,simple_obj_ref_440_scaled);
    array_obj_ref_441_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_441_index_0_rename_ack_0 <= array_obj_ref_441_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_440_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_440_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_441_index_0_resize_req_0,array_obj_ref_441_index_0_resize_ack_0,sl_one,"array_obj_ref_441_index_0_resize ",false,tmp13_438,
    false,simple_obj_ref_440_resized);
    array_obj_ref_441_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_441_index_0_resize_ack_0 <= array_obj_ref_441_index_0_resize_req_0;
      in_aggregated_sig <= tmp13_438;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_440_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_441_offset_inst_req_0,array_obj_ref_441_offset_inst_ack_0,sl_one,"array_obj_ref_441_offset_inst ",false,simple_obj_ref_440_scaled,
    false,array_obj_ref_441_final_offset);
    array_obj_ref_441_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_441_offset_inst_ack_0 <= array_obj_ref_441_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_440_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_441_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_441_root_address_inst_req_0,array_obj_ref_441_root_address_inst_ack_0,sl_one,"array_obj_ref_441_root_address_inst ",false,array_obj_ref_441_final_offset,
    false,array_obj_ref_441_root_address);
    array_obj_ref_441_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_441_root_address_inst_ack_0 <= array_obj_ref_441_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_441_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_441_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_446_index_0_rename_req_0,array_obj_ref_446_index_0_rename_ack_0,sl_one,"array_obj_ref_446_index_0_rename ",false,simple_obj_ref_445_resized,
    false,simple_obj_ref_445_scaled);
    array_obj_ref_446_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_446_index_0_rename_ack_0 <= array_obj_ref_446_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_445_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_445_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_446_index_0_resize_req_0,array_obj_ref_446_index_0_resize_ack_0,sl_one,"array_obj_ref_446_index_0_resize ",false,tmp13_438,
    false,simple_obj_ref_445_resized);
    array_obj_ref_446_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_446_index_0_resize_ack_0 <= array_obj_ref_446_index_0_resize_req_0;
      in_aggregated_sig <= tmp13_438;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_445_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_446_offset_inst_req_0,array_obj_ref_446_offset_inst_ack_0,sl_one,"array_obj_ref_446_offset_inst ",false,simple_obj_ref_445_scaled,
    false,array_obj_ref_446_final_offset);
    array_obj_ref_446_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_446_offset_inst_ack_0 <= array_obj_ref_446_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_445_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_446_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_446_root_address_inst_req_0,array_obj_ref_446_root_address_inst_ack_0,sl_one,"array_obj_ref_446_root_address_inst ",false,array_obj_ref_446_final_offset,
    false,array_obj_ref_446_root_address);
    array_obj_ref_446_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_446_root_address_inst_ack_0 <= array_obj_ref_446_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_446_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_446_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_451_index_0_rename_req_0,array_obj_ref_451_index_0_rename_ack_0,sl_one,"array_obj_ref_451_index_0_rename ",false,simple_obj_ref_450_resized,
    false,simple_obj_ref_450_scaled);
    array_obj_ref_451_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_451_index_0_rename_ack_0 <= array_obj_ref_451_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_450_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_450_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_451_index_0_resize_req_0,array_obj_ref_451_index_0_resize_ack_0,sl_one,"array_obj_ref_451_index_0_resize ",false,tmp13_438,
    false,simple_obj_ref_450_resized);
    array_obj_ref_451_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_451_index_0_resize_ack_0 <= array_obj_ref_451_index_0_resize_req_0;
      in_aggregated_sig <= tmp13_438;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_450_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_451_offset_inst_req_0,array_obj_ref_451_offset_inst_ack_0,sl_one,"array_obj_ref_451_offset_inst ",false,simple_obj_ref_450_scaled,
    false,array_obj_ref_451_final_offset);
    array_obj_ref_451_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_451_offset_inst_ack_0 <= array_obj_ref_451_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_450_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_451_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_451_root_address_inst_req_0,array_obj_ref_451_root_address_inst_ack_0,sl_one,"array_obj_ref_451_root_address_inst ",false,array_obj_ref_451_final_offset,
    false,array_obj_ref_451_root_address);
    array_obj_ref_451_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_451_root_address_inst_ack_0 <= array_obj_ref_451_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_451_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_451_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_462_index_0_rename_req_0,array_obj_ref_462_index_0_rename_ack_0,sl_one,"array_obj_ref_462_index_0_rename ",false,simple_obj_ref_461_resized,
    false,simple_obj_ref_461_scaled);
    array_obj_ref_462_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_462_index_0_rename_ack_0 <= array_obj_ref_462_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_461_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_461_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_462_index_0_resize_req_0,array_obj_ref_462_index_0_resize_ack_0,sl_one,"array_obj_ref_462_index_0_resize ",false,tmp25_459,
    false,simple_obj_ref_461_resized);
    array_obj_ref_462_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_462_index_0_resize_ack_0 <= array_obj_ref_462_index_0_resize_req_0;
      in_aggregated_sig <= tmp25_459;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_461_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_462_offset_inst_req_0,array_obj_ref_462_offset_inst_ack_0,sl_one,"array_obj_ref_462_offset_inst ",false,simple_obj_ref_461_scaled,
    false,array_obj_ref_462_final_offset);
    array_obj_ref_462_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_462_offset_inst_ack_0 <= array_obj_ref_462_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_461_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_462_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_462_root_address_inst_req_0,array_obj_ref_462_root_address_inst_ack_0,sl_one,"array_obj_ref_462_root_address_inst ",false,array_obj_ref_462_final_offset,
    false,array_obj_ref_462_root_address);
    array_obj_ref_462_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_462_root_address_inst_ack_0 <= array_obj_ref_462_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_462_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_462_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_467_index_0_rename_req_0,array_obj_ref_467_index_0_rename_ack_0,sl_one,"array_obj_ref_467_index_0_rename ",false,simple_obj_ref_466_resized,
    false,simple_obj_ref_466_scaled);
    array_obj_ref_467_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_467_index_0_rename_ack_0 <= array_obj_ref_467_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_466_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_466_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_467_index_0_resize_req_0,array_obj_ref_467_index_0_resize_ack_0,sl_one,"array_obj_ref_467_index_0_resize ",false,tmp25_459,
    false,simple_obj_ref_466_resized);
    array_obj_ref_467_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_467_index_0_resize_ack_0 <= array_obj_ref_467_index_0_resize_req_0;
      in_aggregated_sig <= tmp25_459;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_466_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_467_offset_inst_req_0,array_obj_ref_467_offset_inst_ack_0,sl_one,"array_obj_ref_467_offset_inst ",false,simple_obj_ref_466_scaled,
    false,array_obj_ref_467_final_offset);
    array_obj_ref_467_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_467_offset_inst_ack_0 <= array_obj_ref_467_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_466_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_467_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_467_root_address_inst_req_0,array_obj_ref_467_root_address_inst_ack_0,sl_one,"array_obj_ref_467_root_address_inst ",false,array_obj_ref_467_final_offset,
    false,array_obj_ref_467_root_address);
    array_obj_ref_467_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_467_root_address_inst_ack_0 <= array_obj_ref_467_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_467_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_467_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_472_index_0_rename_req_0,array_obj_ref_472_index_0_rename_ack_0,sl_one,"array_obj_ref_472_index_0_rename ",false,simple_obj_ref_471_resized,
    false,simple_obj_ref_471_scaled);
    array_obj_ref_472_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_472_index_0_rename_ack_0 <= array_obj_ref_472_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_471_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_471_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_472_index_0_resize_req_0,array_obj_ref_472_index_0_resize_ack_0,sl_one,"array_obj_ref_472_index_0_resize ",false,tmp25_459,
    false,simple_obj_ref_471_resized);
    array_obj_ref_472_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_472_index_0_resize_ack_0 <= array_obj_ref_472_index_0_resize_req_0;
      in_aggregated_sig <= tmp25_459;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_471_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_472_offset_inst_req_0,array_obj_ref_472_offset_inst_ack_0,sl_one,"array_obj_ref_472_offset_inst ",false,simple_obj_ref_471_scaled,
    false,array_obj_ref_472_final_offset);
    array_obj_ref_472_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_472_offset_inst_ack_0 <= array_obj_ref_472_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_471_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_472_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_472_root_address_inst_req_0,array_obj_ref_472_root_address_inst_ack_0,sl_one,"array_obj_ref_472_root_address_inst ",false,array_obj_ref_472_final_offset,
    false,array_obj_ref_472_root_address);
    array_obj_ref_472_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_472_root_address_inst_ack_0 <= array_obj_ref_472_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_472_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_472_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_483_index_0_rename_req_0,array_obj_ref_483_index_0_rename_ack_0,sl_one,"array_obj_ref_483_index_0_rename ",false,simple_obj_ref_482_resized,
    false,simple_obj_ref_482_scaled);
    array_obj_ref_483_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_483_index_0_rename_ack_0 <= array_obj_ref_483_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_482_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_482_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_483_index_0_resize_req_0,array_obj_ref_483_index_0_resize_ack_0,sl_one,"array_obj_ref_483_index_0_resize ",false,tmp34_480,
    false,simple_obj_ref_482_resized);
    array_obj_ref_483_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_483_index_0_resize_ack_0 <= array_obj_ref_483_index_0_resize_req_0;
      in_aggregated_sig <= tmp34_480;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_482_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_483_offset_inst_req_0,array_obj_ref_483_offset_inst_ack_0,sl_one,"array_obj_ref_483_offset_inst ",false,simple_obj_ref_482_scaled,
    false,array_obj_ref_483_final_offset);
    array_obj_ref_483_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_483_offset_inst_ack_0 <= array_obj_ref_483_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_482_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_483_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_483_root_address_inst_req_0,array_obj_ref_483_root_address_inst_ack_0,sl_one,"array_obj_ref_483_root_address_inst ",false,array_obj_ref_483_final_offset,
    false,array_obj_ref_483_root_address);
    array_obj_ref_483_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_483_root_address_inst_ack_0 <= array_obj_ref_483_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_483_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_483_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_488_index_0_rename_req_0,array_obj_ref_488_index_0_rename_ack_0,sl_one,"array_obj_ref_488_index_0_rename ",false,simple_obj_ref_487_resized,
    false,simple_obj_ref_487_scaled);
    array_obj_ref_488_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_488_index_0_rename_ack_0 <= array_obj_ref_488_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_487_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_487_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_488_index_0_resize_req_0,array_obj_ref_488_index_0_resize_ack_0,sl_one,"array_obj_ref_488_index_0_resize ",false,tmp34_480,
    false,simple_obj_ref_487_resized);
    array_obj_ref_488_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_488_index_0_resize_ack_0 <= array_obj_ref_488_index_0_resize_req_0;
      in_aggregated_sig <= tmp34_480;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_487_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_488_offset_inst_req_0,array_obj_ref_488_offset_inst_ack_0,sl_one,"array_obj_ref_488_offset_inst ",false,simple_obj_ref_487_scaled,
    false,array_obj_ref_488_final_offset);
    array_obj_ref_488_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_488_offset_inst_ack_0 <= array_obj_ref_488_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_487_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_488_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_488_root_address_inst_req_0,array_obj_ref_488_root_address_inst_ack_0,sl_one,"array_obj_ref_488_root_address_inst ",false,array_obj_ref_488_final_offset,
    false,array_obj_ref_488_root_address);
    array_obj_ref_488_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_488_root_address_inst_ack_0 <= array_obj_ref_488_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_488_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_488_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_493_index_0_rename_req_0,array_obj_ref_493_index_0_rename_ack_0,sl_one,"array_obj_ref_493_index_0_rename ",false,simple_obj_ref_492_resized,
    false,simple_obj_ref_492_scaled);
    array_obj_ref_493_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_493_index_0_rename_ack_0 <= array_obj_ref_493_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_492_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_492_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_493_index_0_resize_req_0,array_obj_ref_493_index_0_resize_ack_0,sl_one,"array_obj_ref_493_index_0_resize ",false,tmp34_480,
    false,simple_obj_ref_492_resized);
    array_obj_ref_493_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_493_index_0_resize_ack_0 <= array_obj_ref_493_index_0_resize_req_0;
      in_aggregated_sig <= tmp34_480;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_492_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_493_offset_inst_req_0,array_obj_ref_493_offset_inst_ack_0,sl_one,"array_obj_ref_493_offset_inst ",false,simple_obj_ref_492_scaled,
    false,array_obj_ref_493_final_offset);
    array_obj_ref_493_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_493_offset_inst_ack_0 <= array_obj_ref_493_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_492_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_493_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_493_root_address_inst_req_0,array_obj_ref_493_root_address_inst_ack_0,sl_one,"array_obj_ref_493_root_address_inst ",false,array_obj_ref_493_final_offset,
    false,array_obj_ref_493_root_address);
    array_obj_ref_493_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_493_root_address_inst_ack_0 <= array_obj_ref_493_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_493_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_493_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_504_index_0_rename_req_0,array_obj_ref_504_index_0_rename_ack_0,sl_one,"array_obj_ref_504_index_0_rename ",false,simple_obj_ref_503_resized,
    false,simple_obj_ref_503_scaled);
    array_obj_ref_504_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_504_index_0_rename_ack_0 <= array_obj_ref_504_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_503_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_503_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_504_index_0_resize_req_0,array_obj_ref_504_index_0_resize_ack_0,sl_one,"array_obj_ref_504_index_0_resize ",false,tmp38_501,
    false,simple_obj_ref_503_resized);
    array_obj_ref_504_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_504_index_0_resize_ack_0 <= array_obj_ref_504_index_0_resize_req_0;
      in_aggregated_sig <= tmp38_501;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_503_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_504_offset_inst_req_0,array_obj_ref_504_offset_inst_ack_0,sl_one,"array_obj_ref_504_offset_inst ",false,simple_obj_ref_503_scaled,
    false,array_obj_ref_504_final_offset);
    array_obj_ref_504_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_504_offset_inst_ack_0 <= array_obj_ref_504_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_503_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_504_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_504_root_address_inst_req_0,array_obj_ref_504_root_address_inst_ack_0,sl_one,"array_obj_ref_504_root_address_inst ",false,array_obj_ref_504_final_offset,
    false,array_obj_ref_504_root_address);
    array_obj_ref_504_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_504_root_address_inst_ack_0 <= array_obj_ref_504_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_504_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_504_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_509_index_0_rename_req_0,array_obj_ref_509_index_0_rename_ack_0,sl_one,"array_obj_ref_509_index_0_rename ",false,simple_obj_ref_508_resized,
    false,simple_obj_ref_508_scaled);
    array_obj_ref_509_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_509_index_0_rename_ack_0 <= array_obj_ref_509_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_508_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_508_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_509_index_0_resize_req_0,array_obj_ref_509_index_0_resize_ack_0,sl_one,"array_obj_ref_509_index_0_resize ",false,tmp38_501,
    false,simple_obj_ref_508_resized);
    array_obj_ref_509_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_509_index_0_resize_ack_0 <= array_obj_ref_509_index_0_resize_req_0;
      in_aggregated_sig <= tmp38_501;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_508_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_509_offset_inst_req_0,array_obj_ref_509_offset_inst_ack_0,sl_one,"array_obj_ref_509_offset_inst ",false,simple_obj_ref_508_scaled,
    false,array_obj_ref_509_final_offset);
    array_obj_ref_509_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_509_offset_inst_ack_0 <= array_obj_ref_509_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_508_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_509_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_509_root_address_inst_req_0,array_obj_ref_509_root_address_inst_ack_0,sl_one,"array_obj_ref_509_root_address_inst ",false,array_obj_ref_509_final_offset,
    false,array_obj_ref_509_root_address);
    array_obj_ref_509_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_509_root_address_inst_ack_0 <= array_obj_ref_509_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_509_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_509_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_514_index_0_rename_req_0,array_obj_ref_514_index_0_rename_ack_0,sl_one,"array_obj_ref_514_index_0_rename ",false,simple_obj_ref_513_resized,
    false,simple_obj_ref_513_scaled);
    array_obj_ref_514_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_514_index_0_rename_ack_0 <= array_obj_ref_514_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_513_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_513_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_514_index_0_resize_req_0,array_obj_ref_514_index_0_resize_ack_0,sl_one,"array_obj_ref_514_index_0_resize ",false,tmp38_501,
    false,simple_obj_ref_513_resized);
    array_obj_ref_514_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_514_index_0_resize_ack_0 <= array_obj_ref_514_index_0_resize_req_0;
      in_aggregated_sig <= tmp38_501;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_513_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_514_offset_inst_req_0,array_obj_ref_514_offset_inst_ack_0,sl_one,"array_obj_ref_514_offset_inst ",false,simple_obj_ref_513_scaled,
    false,array_obj_ref_514_final_offset);
    array_obj_ref_514_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_514_offset_inst_ack_0 <= array_obj_ref_514_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_513_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_514_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_514_root_address_inst_req_0,array_obj_ref_514_root_address_inst_ack_0,sl_one,"array_obj_ref_514_root_address_inst ",false,array_obj_ref_514_final_offset,
    false,array_obj_ref_514_root_address);
    array_obj_ref_514_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_514_root_address_inst_ack_0 <= array_obj_ref_514_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_514_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_514_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_525_index_0_rename_req_0,array_obj_ref_525_index_0_rename_ack_0,sl_one,"array_obj_ref_525_index_0_rename ",false,simple_obj_ref_524_resized,
    false,simple_obj_ref_524_scaled);
    array_obj_ref_525_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_525_index_0_rename_ack_0 <= array_obj_ref_525_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_524_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_524_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_525_index_0_resize_req_0,array_obj_ref_525_index_0_resize_ack_0,sl_one,"array_obj_ref_525_index_0_resize ",false,tmp42_522,
    false,simple_obj_ref_524_resized);
    array_obj_ref_525_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_525_index_0_resize_ack_0 <= array_obj_ref_525_index_0_resize_req_0;
      in_aggregated_sig <= tmp42_522;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_524_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_525_offset_inst_req_0,array_obj_ref_525_offset_inst_ack_0,sl_one,"array_obj_ref_525_offset_inst ",false,simple_obj_ref_524_scaled,
    false,array_obj_ref_525_final_offset);
    array_obj_ref_525_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_525_offset_inst_ack_0 <= array_obj_ref_525_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_524_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_525_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_525_root_address_inst_req_0,array_obj_ref_525_root_address_inst_ack_0,sl_one,"array_obj_ref_525_root_address_inst ",false,array_obj_ref_525_final_offset,
    false,array_obj_ref_525_root_address);
    array_obj_ref_525_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_525_root_address_inst_ack_0 <= array_obj_ref_525_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_525_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_525_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_530_index_0_rename_req_0,array_obj_ref_530_index_0_rename_ack_0,sl_one,"array_obj_ref_530_index_0_rename ",false,simple_obj_ref_529_resized,
    false,simple_obj_ref_529_scaled);
    array_obj_ref_530_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_530_index_0_rename_ack_0 <= array_obj_ref_530_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_529_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_529_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_530_index_0_resize_req_0,array_obj_ref_530_index_0_resize_ack_0,sl_one,"array_obj_ref_530_index_0_resize ",false,tmp42_522,
    false,simple_obj_ref_529_resized);
    array_obj_ref_530_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_530_index_0_resize_ack_0 <= array_obj_ref_530_index_0_resize_req_0;
      in_aggregated_sig <= tmp42_522;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_529_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_530_offset_inst_req_0,array_obj_ref_530_offset_inst_ack_0,sl_one,"array_obj_ref_530_offset_inst ",false,simple_obj_ref_529_scaled,
    false,array_obj_ref_530_final_offset);
    array_obj_ref_530_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_530_offset_inst_ack_0 <= array_obj_ref_530_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_529_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_530_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_530_root_address_inst_req_0,array_obj_ref_530_root_address_inst_ack_0,sl_one,"array_obj_ref_530_root_address_inst ",false,array_obj_ref_530_final_offset,
    false,array_obj_ref_530_root_address);
    array_obj_ref_530_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_530_root_address_inst_ack_0 <= array_obj_ref_530_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_530_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_530_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_535_index_0_rename_req_0,array_obj_ref_535_index_0_rename_ack_0,sl_one,"array_obj_ref_535_index_0_rename ",false,simple_obj_ref_534_resized,
    false,simple_obj_ref_534_scaled);
    array_obj_ref_535_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_535_index_0_rename_ack_0 <= array_obj_ref_535_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_534_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_534_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_535_index_0_resize_req_0,array_obj_ref_535_index_0_resize_ack_0,sl_one,"array_obj_ref_535_index_0_resize ",false,tmp42_522,
    false,simple_obj_ref_534_resized);
    array_obj_ref_535_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_535_index_0_resize_ack_0 <= array_obj_ref_535_index_0_resize_req_0;
      in_aggregated_sig <= tmp42_522;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_534_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_535_offset_inst_req_0,array_obj_ref_535_offset_inst_ack_0,sl_one,"array_obj_ref_535_offset_inst ",false,simple_obj_ref_534_scaled,
    false,array_obj_ref_535_final_offset);
    array_obj_ref_535_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_535_offset_inst_ack_0 <= array_obj_ref_535_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_534_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_535_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_535_root_address_inst_req_0,array_obj_ref_535_root_address_inst_ack_0,sl_one,"array_obj_ref_535_root_address_inst ",false,array_obj_ref_535_final_offset,
    false,array_obj_ref_535_root_address);
    array_obj_ref_535_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_535_root_address_inst_ack_0 <= array_obj_ref_535_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_535_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_535_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_546_index_0_rename_req_0,array_obj_ref_546_index_0_rename_ack_0,sl_one,"array_obj_ref_546_index_0_rename ",false,simple_obj_ref_545_resized,
    false,simple_obj_ref_545_scaled);
    array_obj_ref_546_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_546_index_0_rename_ack_0 <= array_obj_ref_546_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_545_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_545_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_546_index_0_resize_req_0,array_obj_ref_546_index_0_resize_ack_0,sl_one,"array_obj_ref_546_index_0_resize ",false,tmp46_543,
    false,simple_obj_ref_545_resized);
    array_obj_ref_546_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_546_index_0_resize_ack_0 <= array_obj_ref_546_index_0_resize_req_0;
      in_aggregated_sig <= tmp46_543;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_545_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_546_offset_inst_req_0,array_obj_ref_546_offset_inst_ack_0,sl_one,"array_obj_ref_546_offset_inst ",false,simple_obj_ref_545_scaled,
    false,array_obj_ref_546_final_offset);
    array_obj_ref_546_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_546_offset_inst_ack_0 <= array_obj_ref_546_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_545_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_546_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_546_root_address_inst_req_0,array_obj_ref_546_root_address_inst_ack_0,sl_one,"array_obj_ref_546_root_address_inst ",false,array_obj_ref_546_final_offset,
    false,array_obj_ref_546_root_address);
    array_obj_ref_546_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_546_root_address_inst_ack_0 <= array_obj_ref_546_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_546_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_546_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_551_index_0_rename_req_0,array_obj_ref_551_index_0_rename_ack_0,sl_one,"array_obj_ref_551_index_0_rename ",false,simple_obj_ref_550_resized,
    false,simple_obj_ref_550_scaled);
    array_obj_ref_551_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_551_index_0_rename_ack_0 <= array_obj_ref_551_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_550_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_550_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_551_index_0_resize_req_0,array_obj_ref_551_index_0_resize_ack_0,sl_one,"array_obj_ref_551_index_0_resize ",false,tmp46_543,
    false,simple_obj_ref_550_resized);
    array_obj_ref_551_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_551_index_0_resize_ack_0 <= array_obj_ref_551_index_0_resize_req_0;
      in_aggregated_sig <= tmp46_543;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_550_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_551_offset_inst_req_0,array_obj_ref_551_offset_inst_ack_0,sl_one,"array_obj_ref_551_offset_inst ",false,simple_obj_ref_550_scaled,
    false,array_obj_ref_551_final_offset);
    array_obj_ref_551_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_551_offset_inst_ack_0 <= array_obj_ref_551_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_550_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_551_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_551_root_address_inst_req_0,array_obj_ref_551_root_address_inst_ack_0,sl_one,"array_obj_ref_551_root_address_inst ",false,array_obj_ref_551_final_offset,
    false,array_obj_ref_551_root_address);
    array_obj_ref_551_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_551_root_address_inst_ack_0 <= array_obj_ref_551_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_551_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_551_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_556_index_0_rename_req_0,array_obj_ref_556_index_0_rename_ack_0,sl_one,"array_obj_ref_556_index_0_rename ",false,simple_obj_ref_555_resized,
    false,simple_obj_ref_555_scaled);
    array_obj_ref_556_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_556_index_0_rename_ack_0 <= array_obj_ref_556_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_555_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_555_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_556_index_0_resize_req_0,array_obj_ref_556_index_0_resize_ack_0,sl_one,"array_obj_ref_556_index_0_resize ",false,tmp46_543,
    false,simple_obj_ref_555_resized);
    array_obj_ref_556_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_556_index_0_resize_ack_0 <= array_obj_ref_556_index_0_resize_req_0;
      in_aggregated_sig <= tmp46_543;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_555_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_556_offset_inst_req_0,array_obj_ref_556_offset_inst_ack_0,sl_one,"array_obj_ref_556_offset_inst ",false,simple_obj_ref_555_scaled,
    false,array_obj_ref_556_final_offset);
    array_obj_ref_556_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_556_offset_inst_ack_0 <= array_obj_ref_556_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_555_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_556_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_556_root_address_inst_req_0,array_obj_ref_556_root_address_inst_ack_0,sl_one,"array_obj_ref_556_root_address_inst ",false,array_obj_ref_556_final_offset,
    false,array_obj_ref_556_root_address);
    array_obj_ref_556_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_556_root_address_inst_ack_0 <= array_obj_ref_556_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_556_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_556_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_561_index_0_rename_req_0,array_obj_ref_561_index_0_rename_ack_0,sl_one,"array_obj_ref_561_index_0_rename ",false,simple_obj_ref_560_resized,
    false,simple_obj_ref_560_scaled);
    array_obj_ref_561_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_561_index_0_rename_ack_0 <= array_obj_ref_561_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_560_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_560_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_561_index_0_resize_req_0,array_obj_ref_561_index_0_resize_ack_0,sl_one,"array_obj_ref_561_index_0_resize ",false,tmp2_411,
    false,simple_obj_ref_560_resized);
    array_obj_ref_561_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_561_index_0_resize_ack_0 <= array_obj_ref_561_index_0_resize_req_0;
      in_aggregated_sig <= tmp2_411;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_560_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_561_offset_inst_req_0,array_obj_ref_561_offset_inst_ack_0,sl_one,"array_obj_ref_561_offset_inst ",false,simple_obj_ref_560_scaled,
    false,array_obj_ref_561_final_offset);
    array_obj_ref_561_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_561_offset_inst_ack_0 <= array_obj_ref_561_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_560_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_561_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_561_root_address_inst_req_0,array_obj_ref_561_root_address_inst_ack_0,sl_one,"array_obj_ref_561_root_address_inst ",false,array_obj_ref_561_final_offset,
    false,array_obj_ref_561_root_address);
    array_obj_ref_561_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_561_root_address_inst_ack_0 <= array_obj_ref_561_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_561_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_561_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_566_index_0_rename_req_0,array_obj_ref_566_index_0_rename_ack_0,sl_one,"array_obj_ref_566_index_0_rename ",false,simple_obj_ref_565_resized,
    false,simple_obj_ref_565_scaled);
    array_obj_ref_566_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_566_index_0_rename_ack_0 <= array_obj_ref_566_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_565_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_565_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_566_index_0_resize_req_0,array_obj_ref_566_index_0_resize_ack_0,sl_one,"array_obj_ref_566_index_0_resize ",false,tmp2_411,
    false,simple_obj_ref_565_resized);
    array_obj_ref_566_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_566_index_0_resize_ack_0 <= array_obj_ref_566_index_0_resize_req_0;
      in_aggregated_sig <= tmp2_411;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_565_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_566_offset_inst_req_0,array_obj_ref_566_offset_inst_ack_0,sl_one,"array_obj_ref_566_offset_inst ",false,simple_obj_ref_565_scaled,
    false,array_obj_ref_566_final_offset);
    array_obj_ref_566_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_566_offset_inst_ack_0 <= array_obj_ref_566_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_565_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_566_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_566_root_address_inst_req_0,array_obj_ref_566_root_address_inst_ack_0,sl_one,"array_obj_ref_566_root_address_inst ",false,array_obj_ref_566_final_offset,
    false,array_obj_ref_566_root_address);
    array_obj_ref_566_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_566_root_address_inst_ack_0 <= array_obj_ref_566_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_566_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_566_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_571_index_0_rename_req_0,array_obj_ref_571_index_0_rename_ack_0,sl_one,"array_obj_ref_571_index_0_rename ",false,simple_obj_ref_570_resized,
    false,simple_obj_ref_570_scaled);
    array_obj_ref_571_index_0_rename: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_571_index_0_rename_ack_0 <= array_obj_ref_571_index_0_rename_req_0;
      in_aggregated_sig <= simple_obj_ref_570_resized;
      out_aggregated_sig <= in_aggregated_sig;
      simple_obj_ref_570_scaled <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_571_index_0_resize_req_0,array_obj_ref_571_index_0_resize_ack_0,sl_one,"array_obj_ref_571_index_0_resize ",false,tmp2_411,
    false,simple_obj_ref_570_resized);
    array_obj_ref_571_index_0_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_571_index_0_resize_ack_0 <= array_obj_ref_571_index_0_resize_req_0;
      in_aggregated_sig <= tmp2_411;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      simple_obj_ref_570_resized <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_571_offset_inst_req_0,array_obj_ref_571_offset_inst_ack_0,sl_one,"array_obj_ref_571_offset_inst ",false,simple_obj_ref_570_scaled,
    false,array_obj_ref_571_final_offset);
    array_obj_ref_571_offset_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_571_offset_inst_ack_0 <= array_obj_ref_571_offset_inst_req_0;
      in_aggregated_sig <= simple_obj_ref_570_scaled;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_571_final_offset <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,array_obj_ref_571_root_address_inst_req_0,array_obj_ref_571_root_address_inst_ack_0,sl_one,"array_obj_ref_571_root_address_inst ",false,array_obj_ref_571_final_offset,
    false,array_obj_ref_571_root_address);
    array_obj_ref_571_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      array_obj_ref_571_root_address_inst_ack_0 <= array_obj_ref_571_root_address_inst_req_0;
      in_aggregated_sig <= array_obj_ref_571_final_offset;
      out_aggregated_sig <= in_aggregated_sig;
      array_obj_ref_571_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_576_addr_0_req_0,ptr_deref_576_addr_0_ack_0,sl_one,"ptr_deref_576_addr_0 ",false,ptr_deref_576_root_address,
    false,ptr_deref_576_word_address_0);
    ptr_deref_576_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_576_addr_0_ack_0 <= ptr_deref_576_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_576_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_576_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_576_base_resize_req_0,ptr_deref_576_base_resize_ack_0,sl_one,"ptr_deref_576_base_resize ",false,scevgep_573,
    false,ptr_deref_576_resized_base_address);
    ptr_deref_576_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_576_base_resize_ack_0 <= ptr_deref_576_base_resize_req_0;
      in_aggregated_sig <= scevgep_573;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_576_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_576_gather_scatter_req_0,ptr_deref_576_gather_scatter_ack_0,sl_one,"ptr_deref_576_gather_scatter ",false,ptr_deref_576_data_0,
    false,iNsTr_2_577);
    ptr_deref_576_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_576_gather_scatter_ack_0 <= ptr_deref_576_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_576_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_2_577 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_576_root_address_inst_req_0,ptr_deref_576_root_address_inst_ack_0,sl_one,"ptr_deref_576_root_address_inst ",false,ptr_deref_576_resized_base_address,
    false,ptr_deref_576_root_address);
    ptr_deref_576_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_576_root_address_inst_ack_0 <= ptr_deref_576_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_576_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_576_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_580_addr_0_req_0,ptr_deref_580_addr_0_ack_0,sl_one,"ptr_deref_580_addr_0 ",false,ptr_deref_580_root_address,
    false,ptr_deref_580_word_address_0);
    ptr_deref_580_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_580_addr_0_ack_0 <= ptr_deref_580_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_580_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_580_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_580_base_resize_req_0,ptr_deref_580_base_resize_ack_0,sl_one,"ptr_deref_580_base_resize ",false,scevgep2_568,
    false,ptr_deref_580_resized_base_address);
    ptr_deref_580_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_580_base_resize_ack_0 <= ptr_deref_580_base_resize_req_0;
      in_aggregated_sig <= scevgep2_568;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_580_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_580_gather_scatter_req_0,ptr_deref_580_gather_scatter_ack_0,sl_one,"ptr_deref_580_gather_scatter ",false,ptr_deref_580_data_0,
    false,iNsTr_3_581);
    ptr_deref_580_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_580_gather_scatter_ack_0 <= ptr_deref_580_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_580_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_3_581 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_580_root_address_inst_req_0,ptr_deref_580_root_address_inst_ack_0,sl_one,"ptr_deref_580_root_address_inst ",false,ptr_deref_580_resized_base_address,
    false,ptr_deref_580_root_address);
    ptr_deref_580_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_580_root_address_inst_ack_0 <= ptr_deref_580_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_580_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_580_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_589_addr_0_req_0,ptr_deref_589_addr_0_ack_0,sl_one,"ptr_deref_589_addr_0 ",false,ptr_deref_589_root_address,
    false,ptr_deref_589_word_address_0);
    ptr_deref_589_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_589_addr_0_ack_0 <= ptr_deref_589_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_589_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_589_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_589_base_resize_req_0,ptr_deref_589_base_resize_ack_0,sl_one,"ptr_deref_589_base_resize ",false,scevgep5_558,
    false,ptr_deref_589_resized_base_address);
    ptr_deref_589_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_589_base_resize_ack_0 <= ptr_deref_589_base_resize_req_0;
      in_aggregated_sig <= scevgep5_558;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_589_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_589_gather_scatter_req_0,ptr_deref_589_gather_scatter_ack_0,sl_one,"ptr_deref_589_gather_scatter ",false,ptr_deref_589_data_0,
    false,iNsTr_5_590);
    ptr_deref_589_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_589_gather_scatter_ack_0 <= ptr_deref_589_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_589_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_5_590 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_589_root_address_inst_req_0,ptr_deref_589_root_address_inst_ack_0,sl_one,"ptr_deref_589_root_address_inst ",false,ptr_deref_589_resized_base_address,
    false,ptr_deref_589_root_address);
    ptr_deref_589_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_589_root_address_inst_ack_0 <= ptr_deref_589_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_589_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_589_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_593_addr_0_req_0,ptr_deref_593_addr_0_ack_0,sl_one,"ptr_deref_593_addr_0 ",false,ptr_deref_593_root_address,
    false,ptr_deref_593_word_address_0);
    ptr_deref_593_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_593_addr_0_ack_0 <= ptr_deref_593_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_593_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_593_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_593_base_resize_req_0,ptr_deref_593_base_resize_ack_0,sl_one,"ptr_deref_593_base_resize ",false,scevgep6_553,
    false,ptr_deref_593_resized_base_address);
    ptr_deref_593_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_593_base_resize_ack_0 <= ptr_deref_593_base_resize_req_0;
      in_aggregated_sig <= scevgep6_553;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_593_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_593_gather_scatter_req_0,ptr_deref_593_gather_scatter_ack_0,sl_one,"ptr_deref_593_gather_scatter ",false,ptr_deref_593_data_0,
    false,iNsTr_6_594);
    ptr_deref_593_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_593_gather_scatter_ack_0 <= ptr_deref_593_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_593_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_6_594 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_593_root_address_inst_req_0,ptr_deref_593_root_address_inst_ack_0,sl_one,"ptr_deref_593_root_address_inst ",false,ptr_deref_593_resized_base_address,
    false,ptr_deref_593_root_address);
    ptr_deref_593_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_593_root_address_inst_ack_0 <= ptr_deref_593_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_593_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_593_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_602_addr_0_req_0,ptr_deref_602_addr_0_ack_0,sl_one,"ptr_deref_602_addr_0 ",false,ptr_deref_602_root_address,
    false,ptr_deref_602_word_address_0);
    ptr_deref_602_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_602_addr_0_ack_0 <= ptr_deref_602_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_602_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_602_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_602_base_resize_req_0,ptr_deref_602_base_resize_ack_0,sl_one,"ptr_deref_602_base_resize ",false,scevgep9_537,
    false,ptr_deref_602_resized_base_address);
    ptr_deref_602_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_602_base_resize_ack_0 <= ptr_deref_602_base_resize_req_0;
      in_aggregated_sig <= scevgep9_537;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_602_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_602_gather_scatter_req_0,ptr_deref_602_gather_scatter_ack_0,sl_one,"ptr_deref_602_gather_scatter ",false,ptr_deref_602_data_0,
    false,iNsTr_8_603);
    ptr_deref_602_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_602_gather_scatter_ack_0 <= ptr_deref_602_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_602_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_8_603 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_602_root_address_inst_req_0,ptr_deref_602_root_address_inst_ack_0,sl_one,"ptr_deref_602_root_address_inst ",false,ptr_deref_602_resized_base_address,
    false,ptr_deref_602_root_address);
    ptr_deref_602_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_602_root_address_inst_ack_0 <= ptr_deref_602_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_602_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_602_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_606_addr_0_req_0,ptr_deref_606_addr_0_ack_0,sl_one,"ptr_deref_606_addr_0 ",false,ptr_deref_606_root_address,
    false,ptr_deref_606_word_address_0);
    ptr_deref_606_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_606_addr_0_ack_0 <= ptr_deref_606_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_606_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_606_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_606_base_resize_req_0,ptr_deref_606_base_resize_ack_0,sl_one,"ptr_deref_606_base_resize ",false,scevgep10_532,
    false,ptr_deref_606_resized_base_address);
    ptr_deref_606_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_606_base_resize_ack_0 <= ptr_deref_606_base_resize_req_0;
      in_aggregated_sig <= scevgep10_532;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_606_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_606_gather_scatter_req_0,ptr_deref_606_gather_scatter_ack_0,sl_one,"ptr_deref_606_gather_scatter ",false,ptr_deref_606_data_0,
    false,iNsTr_9_607);
    ptr_deref_606_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_606_gather_scatter_ack_0 <= ptr_deref_606_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_606_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_9_607 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_606_root_address_inst_req_0,ptr_deref_606_root_address_inst_ack_0,sl_one,"ptr_deref_606_root_address_inst ",false,ptr_deref_606_resized_base_address,
    false,ptr_deref_606_root_address);
    ptr_deref_606_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_606_root_address_inst_ack_0 <= ptr_deref_606_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_606_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_606_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_615_addr_0_req_0,ptr_deref_615_addr_0_ack_0,sl_one,"ptr_deref_615_addr_0 ",false,ptr_deref_615_root_address,
    false,ptr_deref_615_word_address_0);
    ptr_deref_615_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_615_addr_0_ack_0 <= ptr_deref_615_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_615_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_615_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_615_base_resize_req_0,ptr_deref_615_base_resize_ack_0,sl_one,"ptr_deref_615_base_resize ",false,scevgep13_516,
    false,ptr_deref_615_resized_base_address);
    ptr_deref_615_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_615_base_resize_ack_0 <= ptr_deref_615_base_resize_req_0;
      in_aggregated_sig <= scevgep13_516;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_615_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_615_gather_scatter_req_0,ptr_deref_615_gather_scatter_ack_0,sl_one,"ptr_deref_615_gather_scatter ",false,ptr_deref_615_data_0,
    false,iNsTr_11_616);
    ptr_deref_615_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_615_gather_scatter_ack_0 <= ptr_deref_615_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_615_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_11_616 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_615_root_address_inst_req_0,ptr_deref_615_root_address_inst_ack_0,sl_one,"ptr_deref_615_root_address_inst ",false,ptr_deref_615_resized_base_address,
    false,ptr_deref_615_root_address);
    ptr_deref_615_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_615_root_address_inst_ack_0 <= ptr_deref_615_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_615_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_615_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_619_addr_0_req_0,ptr_deref_619_addr_0_ack_0,sl_one,"ptr_deref_619_addr_0 ",false,ptr_deref_619_root_address,
    false,ptr_deref_619_word_address_0);
    ptr_deref_619_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_619_addr_0_ack_0 <= ptr_deref_619_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_619_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_619_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_619_base_resize_req_0,ptr_deref_619_base_resize_ack_0,sl_one,"ptr_deref_619_base_resize ",false,scevgep14_511,
    false,ptr_deref_619_resized_base_address);
    ptr_deref_619_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_619_base_resize_ack_0 <= ptr_deref_619_base_resize_req_0;
      in_aggregated_sig <= scevgep14_511;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_619_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_619_gather_scatter_req_0,ptr_deref_619_gather_scatter_ack_0,sl_one,"ptr_deref_619_gather_scatter ",false,ptr_deref_619_data_0,
    false,iNsTr_12_620);
    ptr_deref_619_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_619_gather_scatter_ack_0 <= ptr_deref_619_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_619_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_12_620 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_619_root_address_inst_req_0,ptr_deref_619_root_address_inst_ack_0,sl_one,"ptr_deref_619_root_address_inst ",false,ptr_deref_619_resized_base_address,
    false,ptr_deref_619_root_address);
    ptr_deref_619_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_619_root_address_inst_ack_0 <= ptr_deref_619_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_619_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_619_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_628_addr_0_req_0,ptr_deref_628_addr_0_ack_0,sl_one,"ptr_deref_628_addr_0 ",false,ptr_deref_628_root_address,
    false,ptr_deref_628_word_address_0);
    ptr_deref_628_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_628_addr_0_ack_0 <= ptr_deref_628_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_628_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_628_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_628_base_resize_req_0,ptr_deref_628_base_resize_ack_0,sl_one,"ptr_deref_628_base_resize ",false,scevgep17_495,
    false,ptr_deref_628_resized_base_address);
    ptr_deref_628_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_628_base_resize_ack_0 <= ptr_deref_628_base_resize_req_0;
      in_aggregated_sig <= scevgep17_495;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_628_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_628_gather_scatter_req_0,ptr_deref_628_gather_scatter_ack_0,sl_one,"ptr_deref_628_gather_scatter ",false,ptr_deref_628_data_0,
    false,iNsTr_14_629);
    ptr_deref_628_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_628_gather_scatter_ack_0 <= ptr_deref_628_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_628_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_14_629 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_628_root_address_inst_req_0,ptr_deref_628_root_address_inst_ack_0,sl_one,"ptr_deref_628_root_address_inst ",false,ptr_deref_628_resized_base_address,
    false,ptr_deref_628_root_address);
    ptr_deref_628_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_628_root_address_inst_ack_0 <= ptr_deref_628_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_628_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_628_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_632_addr_0_req_0,ptr_deref_632_addr_0_ack_0,sl_one,"ptr_deref_632_addr_0 ",false,ptr_deref_632_root_address,
    false,ptr_deref_632_word_address_0);
    ptr_deref_632_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_632_addr_0_ack_0 <= ptr_deref_632_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_632_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_632_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_632_base_resize_req_0,ptr_deref_632_base_resize_ack_0,sl_one,"ptr_deref_632_base_resize ",false,scevgep18_490,
    false,ptr_deref_632_resized_base_address);
    ptr_deref_632_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_632_base_resize_ack_0 <= ptr_deref_632_base_resize_req_0;
      in_aggregated_sig <= scevgep18_490;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_632_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_632_gather_scatter_req_0,ptr_deref_632_gather_scatter_ack_0,sl_one,"ptr_deref_632_gather_scatter ",false,ptr_deref_632_data_0,
    false,iNsTr_15_633);
    ptr_deref_632_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_632_gather_scatter_ack_0 <= ptr_deref_632_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_632_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_15_633 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_632_root_address_inst_req_0,ptr_deref_632_root_address_inst_ack_0,sl_one,"ptr_deref_632_root_address_inst ",false,ptr_deref_632_resized_base_address,
    false,ptr_deref_632_root_address);
    ptr_deref_632_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_632_root_address_inst_ack_0 <= ptr_deref_632_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_632_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_632_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_641_addr_0_req_0,ptr_deref_641_addr_0_ack_0,sl_one,"ptr_deref_641_addr_0 ",false,ptr_deref_641_root_address,
    false,ptr_deref_641_word_address_0);
    ptr_deref_641_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_641_addr_0_ack_0 <= ptr_deref_641_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_641_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_641_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_641_base_resize_req_0,ptr_deref_641_base_resize_ack_0,sl_one,"ptr_deref_641_base_resize ",false,scevgep21_474,
    false,ptr_deref_641_resized_base_address);
    ptr_deref_641_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_641_base_resize_ack_0 <= ptr_deref_641_base_resize_req_0;
      in_aggregated_sig <= scevgep21_474;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_641_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_641_gather_scatter_req_0,ptr_deref_641_gather_scatter_ack_0,sl_one,"ptr_deref_641_gather_scatter ",false,ptr_deref_641_data_0,
    false,iNsTr_17_642);
    ptr_deref_641_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_641_gather_scatter_ack_0 <= ptr_deref_641_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_641_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_17_642 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_641_root_address_inst_req_0,ptr_deref_641_root_address_inst_ack_0,sl_one,"ptr_deref_641_root_address_inst ",false,ptr_deref_641_resized_base_address,
    false,ptr_deref_641_root_address);
    ptr_deref_641_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_641_root_address_inst_ack_0 <= ptr_deref_641_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_641_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_641_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_645_addr_0_req_0,ptr_deref_645_addr_0_ack_0,sl_one,"ptr_deref_645_addr_0 ",false,ptr_deref_645_root_address,
    false,ptr_deref_645_word_address_0);
    ptr_deref_645_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_645_addr_0_ack_0 <= ptr_deref_645_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_645_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_645_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_645_base_resize_req_0,ptr_deref_645_base_resize_ack_0,sl_one,"ptr_deref_645_base_resize ",false,scevgep22_469,
    false,ptr_deref_645_resized_base_address);
    ptr_deref_645_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_645_base_resize_ack_0 <= ptr_deref_645_base_resize_req_0;
      in_aggregated_sig <= scevgep22_469;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_645_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_645_gather_scatter_req_0,ptr_deref_645_gather_scatter_ack_0,sl_one,"ptr_deref_645_gather_scatter ",false,ptr_deref_645_data_0,
    false,iNsTr_18_646);
    ptr_deref_645_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_645_gather_scatter_ack_0 <= ptr_deref_645_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_645_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_18_646 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_645_root_address_inst_req_0,ptr_deref_645_root_address_inst_ack_0,sl_one,"ptr_deref_645_root_address_inst ",false,ptr_deref_645_resized_base_address,
    false,ptr_deref_645_root_address);
    ptr_deref_645_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_645_root_address_inst_ack_0 <= ptr_deref_645_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_645_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_645_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_654_addr_0_req_0,ptr_deref_654_addr_0_ack_0,sl_one,"ptr_deref_654_addr_0 ",false,ptr_deref_654_root_address,
    false,ptr_deref_654_word_address_0);
    ptr_deref_654_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_654_addr_0_ack_0 <= ptr_deref_654_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_654_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_654_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_654_base_resize_req_0,ptr_deref_654_base_resize_ack_0,sl_one,"ptr_deref_654_base_resize ",false,scevgep25_453,
    false,ptr_deref_654_resized_base_address);
    ptr_deref_654_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_654_base_resize_ack_0 <= ptr_deref_654_base_resize_req_0;
      in_aggregated_sig <= scevgep25_453;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_654_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_654_gather_scatter_req_0,ptr_deref_654_gather_scatter_ack_0,sl_one,"ptr_deref_654_gather_scatter ",false,ptr_deref_654_data_0,
    false,iNsTr_20_655);
    ptr_deref_654_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_654_gather_scatter_ack_0 <= ptr_deref_654_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_654_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_20_655 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_654_root_address_inst_req_0,ptr_deref_654_root_address_inst_ack_0,sl_one,"ptr_deref_654_root_address_inst ",false,ptr_deref_654_resized_base_address,
    false,ptr_deref_654_root_address);
    ptr_deref_654_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_654_root_address_inst_ack_0 <= ptr_deref_654_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_654_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_654_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_658_addr_0_req_0,ptr_deref_658_addr_0_ack_0,sl_one,"ptr_deref_658_addr_0 ",false,ptr_deref_658_root_address,
    false,ptr_deref_658_word_address_0);
    ptr_deref_658_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_658_addr_0_ack_0 <= ptr_deref_658_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_658_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_658_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_658_base_resize_req_0,ptr_deref_658_base_resize_ack_0,sl_one,"ptr_deref_658_base_resize ",false,scevgep26_448,
    false,ptr_deref_658_resized_base_address);
    ptr_deref_658_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_658_base_resize_ack_0 <= ptr_deref_658_base_resize_req_0;
      in_aggregated_sig <= scevgep26_448;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_658_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_658_gather_scatter_req_0,ptr_deref_658_gather_scatter_ack_0,sl_one,"ptr_deref_658_gather_scatter ",false,ptr_deref_658_data_0,
    false,iNsTr_21_659);
    ptr_deref_658_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_658_gather_scatter_ack_0 <= ptr_deref_658_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_658_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_21_659 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_658_root_address_inst_req_0,ptr_deref_658_root_address_inst_ack_0,sl_one,"ptr_deref_658_root_address_inst ",false,ptr_deref_658_resized_base_address,
    false,ptr_deref_658_root_address);
    ptr_deref_658_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_658_root_address_inst_ack_0 <= ptr_deref_658_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_658_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_658_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_667_addr_0_req_0,ptr_deref_667_addr_0_ack_0,sl_one,"ptr_deref_667_addr_0 ",false,ptr_deref_667_root_address,
    false,ptr_deref_667_word_address_0);
    ptr_deref_667_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_667_addr_0_ack_0 <= ptr_deref_667_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_667_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_667_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_667_base_resize_req_0,ptr_deref_667_base_resize_ack_0,sl_one,"ptr_deref_667_base_resize ",false,scevgep29_432,
    false,ptr_deref_667_resized_base_address);
    ptr_deref_667_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_667_base_resize_ack_0 <= ptr_deref_667_base_resize_req_0;
      in_aggregated_sig <= scevgep29_432;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_667_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_667_gather_scatter_req_0,ptr_deref_667_gather_scatter_ack_0,sl_one,"ptr_deref_667_gather_scatter ",false,ptr_deref_667_data_0,
    false,iNsTr_23_668);
    ptr_deref_667_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_667_gather_scatter_ack_0 <= ptr_deref_667_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_667_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_23_668 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_667_root_address_inst_req_0,ptr_deref_667_root_address_inst_ack_0,sl_one,"ptr_deref_667_root_address_inst ",false,ptr_deref_667_resized_base_address,
    false,ptr_deref_667_root_address);
    ptr_deref_667_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_667_root_address_inst_ack_0 <= ptr_deref_667_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_667_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_667_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_671_addr_0_req_0,ptr_deref_671_addr_0_ack_0,sl_one,"ptr_deref_671_addr_0 ",false,ptr_deref_671_root_address,
    false,ptr_deref_671_word_address_0);
    ptr_deref_671_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_671_addr_0_ack_0 <= ptr_deref_671_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_671_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_671_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_671_base_resize_req_0,ptr_deref_671_base_resize_ack_0,sl_one,"ptr_deref_671_base_resize ",false,scevgep30_427,
    false,ptr_deref_671_resized_base_address);
    ptr_deref_671_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_671_base_resize_ack_0 <= ptr_deref_671_base_resize_req_0;
      in_aggregated_sig <= scevgep30_427;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_671_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_671_gather_scatter_req_0,ptr_deref_671_gather_scatter_ack_0,sl_one,"ptr_deref_671_gather_scatter ",false,ptr_deref_671_data_0,
    false,iNsTr_24_672);
    ptr_deref_671_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_671_gather_scatter_ack_0 <= ptr_deref_671_gather_scatter_req_0;
      in_aggregated_sig <= ptr_deref_671_data_0;
      out_aggregated_sig <= in_aggregated_sig;
      iNsTr_24_672 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_671_root_address_inst_req_0,ptr_deref_671_root_address_inst_ack_0,sl_one,"ptr_deref_671_root_address_inst ",false,ptr_deref_671_resized_base_address,
    false,ptr_deref_671_root_address);
    ptr_deref_671_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_671_root_address_inst_ack_0 <= ptr_deref_671_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_671_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_671_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_694_addr_0_req_0,ptr_deref_694_addr_0_ack_0,sl_one,"ptr_deref_694_addr_0 ",false,ptr_deref_694_root_address,
    false,ptr_deref_694_word_address_0);
    ptr_deref_694_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_694_addr_0_ack_0 <= ptr_deref_694_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_694_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_694_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_694_base_resize_req_0,ptr_deref_694_base_resize_ack_0,sl_one,"ptr_deref_694_base_resize ",false,scevgep3_678_delayed_4_692,
    false,ptr_deref_694_resized_base_address);
    ptr_deref_694_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_694_base_resize_ack_0 <= ptr_deref_694_base_resize_req_0;
      in_aggregated_sig <= scevgep3_678_delayed_4_692;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_694_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_694_gather_scatter_req_0,ptr_deref_694_gather_scatter_ack_0,sl_one,"ptr_deref_694_gather_scatter ",false,iNsTr_4_586,
    false,ptr_deref_694_data_0);
    ptr_deref_694_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_694_gather_scatter_ack_0 <= ptr_deref_694_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_4_586;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_694_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_694_root_address_inst_req_0,ptr_deref_694_root_address_inst_ack_0,sl_one,"ptr_deref_694_root_address_inst ",false,ptr_deref_694_resized_base_address,
    false,ptr_deref_694_root_address);
    ptr_deref_694_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_694_root_address_inst_ack_0 <= ptr_deref_694_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_694_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_694_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_713_addr_0_req_0,ptr_deref_713_addr_0_ack_0,sl_one,"ptr_deref_713_addr_0 ",false,ptr_deref_713_root_address,
    false,ptr_deref_713_word_address_0);
    ptr_deref_713_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_713_addr_0_ack_0 <= ptr_deref_713_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_713_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_713_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_713_base_resize_req_0,ptr_deref_713_base_resize_ack_0,sl_one,"ptr_deref_713_base_resize ",false,scevgep7_682_delayed_4_711,
    false,ptr_deref_713_resized_base_address);
    ptr_deref_713_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_713_base_resize_ack_0 <= ptr_deref_713_base_resize_req_0;
      in_aggregated_sig <= scevgep7_682_delayed_4_711;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_713_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_713_gather_scatter_req_0,ptr_deref_713_gather_scatter_ack_0,sl_one,"ptr_deref_713_gather_scatter ",false,iNsTr_7_599,
    false,ptr_deref_713_data_0);
    ptr_deref_713_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_713_gather_scatter_ack_0 <= ptr_deref_713_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_7_599;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_713_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_713_root_address_inst_req_0,ptr_deref_713_root_address_inst_ack_0,sl_one,"ptr_deref_713_root_address_inst ",false,ptr_deref_713_resized_base_address,
    false,ptr_deref_713_root_address);
    ptr_deref_713_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_713_root_address_inst_ack_0 <= ptr_deref_713_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_713_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_713_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_732_addr_0_req_0,ptr_deref_732_addr_0_ack_0,sl_one,"ptr_deref_732_addr_0 ",false,ptr_deref_732_root_address,
    false,ptr_deref_732_word_address_0);
    ptr_deref_732_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_732_addr_0_ack_0 <= ptr_deref_732_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_732_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_732_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_732_base_resize_req_0,ptr_deref_732_base_resize_ack_0,sl_one,"ptr_deref_732_base_resize ",false,scevgep11_686_delayed_4_730,
    false,ptr_deref_732_resized_base_address);
    ptr_deref_732_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_732_base_resize_ack_0 <= ptr_deref_732_base_resize_req_0;
      in_aggregated_sig <= scevgep11_686_delayed_4_730;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_732_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_732_gather_scatter_req_0,ptr_deref_732_gather_scatter_ack_0,sl_one,"ptr_deref_732_gather_scatter ",false,iNsTr_10_612,
    false,ptr_deref_732_data_0);
    ptr_deref_732_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_732_gather_scatter_ack_0 <= ptr_deref_732_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_10_612;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_732_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_732_root_address_inst_req_0,ptr_deref_732_root_address_inst_ack_0,sl_one,"ptr_deref_732_root_address_inst ",false,ptr_deref_732_resized_base_address,
    false,ptr_deref_732_root_address);
    ptr_deref_732_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_732_root_address_inst_ack_0 <= ptr_deref_732_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_732_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_732_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_751_addr_0_req_0,ptr_deref_751_addr_0_ack_0,sl_one,"ptr_deref_751_addr_0 ",false,ptr_deref_751_root_address,
    false,ptr_deref_751_word_address_0);
    ptr_deref_751_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_751_addr_0_ack_0 <= ptr_deref_751_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_751_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_751_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_751_base_resize_req_0,ptr_deref_751_base_resize_ack_0,sl_one,"ptr_deref_751_base_resize ",false,scevgep15_690_delayed_4_749,
    false,ptr_deref_751_resized_base_address);
    ptr_deref_751_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_751_base_resize_ack_0 <= ptr_deref_751_base_resize_req_0;
      in_aggregated_sig <= scevgep15_690_delayed_4_749;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_751_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_751_gather_scatter_req_0,ptr_deref_751_gather_scatter_ack_0,sl_one,"ptr_deref_751_gather_scatter ",false,iNsTr_13_625,
    false,ptr_deref_751_data_0);
    ptr_deref_751_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_751_gather_scatter_ack_0 <= ptr_deref_751_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_13_625;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_751_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_751_root_address_inst_req_0,ptr_deref_751_root_address_inst_ack_0,sl_one,"ptr_deref_751_root_address_inst ",false,ptr_deref_751_resized_base_address,
    false,ptr_deref_751_root_address);
    ptr_deref_751_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_751_root_address_inst_ack_0 <= ptr_deref_751_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_751_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_751_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_770_addr_0_req_0,ptr_deref_770_addr_0_ack_0,sl_one,"ptr_deref_770_addr_0 ",false,ptr_deref_770_root_address,
    false,ptr_deref_770_word_address_0);
    ptr_deref_770_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_770_addr_0_ack_0 <= ptr_deref_770_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_770_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_770_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_770_base_resize_req_0,ptr_deref_770_base_resize_ack_0,sl_one,"ptr_deref_770_base_resize ",false,scevgep19_694_delayed_4_768,
    false,ptr_deref_770_resized_base_address);
    ptr_deref_770_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_770_base_resize_ack_0 <= ptr_deref_770_base_resize_req_0;
      in_aggregated_sig <= scevgep19_694_delayed_4_768;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_770_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_770_gather_scatter_req_0,ptr_deref_770_gather_scatter_ack_0,sl_one,"ptr_deref_770_gather_scatter ",false,iNsTr_16_638,
    false,ptr_deref_770_data_0);
    ptr_deref_770_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_770_gather_scatter_ack_0 <= ptr_deref_770_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_16_638;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_770_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_770_root_address_inst_req_0,ptr_deref_770_root_address_inst_ack_0,sl_one,"ptr_deref_770_root_address_inst ",false,ptr_deref_770_resized_base_address,
    false,ptr_deref_770_root_address);
    ptr_deref_770_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_770_root_address_inst_ack_0 <= ptr_deref_770_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_770_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_770_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_789_addr_0_req_0,ptr_deref_789_addr_0_ack_0,sl_one,"ptr_deref_789_addr_0 ",false,ptr_deref_789_root_address,
    false,ptr_deref_789_word_address_0);
    ptr_deref_789_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_789_addr_0_ack_0 <= ptr_deref_789_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_789_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_789_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_789_base_resize_req_0,ptr_deref_789_base_resize_ack_0,sl_one,"ptr_deref_789_base_resize ",false,scevgep23_698_delayed_4_787,
    false,ptr_deref_789_resized_base_address);
    ptr_deref_789_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_789_base_resize_ack_0 <= ptr_deref_789_base_resize_req_0;
      in_aggregated_sig <= scevgep23_698_delayed_4_787;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_789_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_789_gather_scatter_req_0,ptr_deref_789_gather_scatter_ack_0,sl_one,"ptr_deref_789_gather_scatter ",false,iNsTr_19_651,
    false,ptr_deref_789_data_0);
    ptr_deref_789_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_789_gather_scatter_ack_0 <= ptr_deref_789_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_19_651;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_789_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_789_root_address_inst_req_0,ptr_deref_789_root_address_inst_ack_0,sl_one,"ptr_deref_789_root_address_inst ",false,ptr_deref_789_resized_base_address,
    false,ptr_deref_789_root_address);
    ptr_deref_789_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_789_root_address_inst_ack_0 <= ptr_deref_789_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_789_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_789_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_808_addr_0_req_0,ptr_deref_808_addr_0_ack_0,sl_one,"ptr_deref_808_addr_0 ",false,ptr_deref_808_root_address,
    false,ptr_deref_808_word_address_0);
    ptr_deref_808_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_808_addr_0_ack_0 <= ptr_deref_808_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_808_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_808_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_808_base_resize_req_0,ptr_deref_808_base_resize_ack_0,sl_one,"ptr_deref_808_base_resize ",false,scevgep27_702_delayed_4_806,
    false,ptr_deref_808_resized_base_address);
    ptr_deref_808_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_808_base_resize_ack_0 <= ptr_deref_808_base_resize_req_0;
      in_aggregated_sig <= scevgep27_702_delayed_4_806;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_808_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_808_gather_scatter_req_0,ptr_deref_808_gather_scatter_ack_0,sl_one,"ptr_deref_808_gather_scatter ",false,iNsTr_22_664,
    false,ptr_deref_808_data_0);
    ptr_deref_808_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_808_gather_scatter_ack_0 <= ptr_deref_808_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_22_664;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_808_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_808_root_address_inst_req_0,ptr_deref_808_root_address_inst_ack_0,sl_one,"ptr_deref_808_root_address_inst ",false,ptr_deref_808_resized_base_address,
    false,ptr_deref_808_root_address);
    ptr_deref_808_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_808_root_address_inst_ack_0 <= ptr_deref_808_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_808_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_808_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_827_addr_0_req_0,ptr_deref_827_addr_0_ack_0,sl_one,"ptr_deref_827_addr_0 ",false,ptr_deref_827_root_address,
    false,ptr_deref_827_word_address_0);
    ptr_deref_827_addr_0: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_827_addr_0_ack_0 <= ptr_deref_827_addr_0_req_0;
      in_aggregated_sig <= ptr_deref_827_root_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_827_word_address_0 <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_827_base_resize_req_0,ptr_deref_827_base_resize_ack_0,sl_one,"ptr_deref_827_base_resize ",false,scevgep31_706_delayed_4_825,
    false,ptr_deref_827_resized_base_address);
    ptr_deref_827_base_resize: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_827_base_resize_ack_0 <= ptr_deref_827_base_resize_req_0;
      in_aggregated_sig <= scevgep31_706_delayed_4_825;
      out_aggregated_sig <= in_aggregated_sig(6 downto 0);
      ptr_deref_827_resized_base_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_827_gather_scatter_req_0,ptr_deref_827_gather_scatter_ack_0,sl_one,"ptr_deref_827_gather_scatter ",false,iNsTr_25_677,
    false,ptr_deref_827_data_0);
    ptr_deref_827_gather_scatter: Block -- 
      signal in_aggregated_sig: std_logic_vector(31 downto 0);
      signal out_aggregated_sig: std_logic_vector(31 downto 0);
      --
    begin -- 
      ptr_deref_827_gather_scatter_ack_0 <= ptr_deref_827_gather_scatter_req_0;
      in_aggregated_sig <= iNsTr_25_677;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_827_data_0 <= out_aggregated_sig(31 downto 0);
      --
    end Block;
    LogOperator(clk,reset,global_clock_cycle_count,ptr_deref_827_root_address_inst_req_0,ptr_deref_827_root_address_inst_ack_0,sl_one,"ptr_deref_827_root_address_inst ",false,ptr_deref_827_resized_base_address,
    false,ptr_deref_827_root_address);
    ptr_deref_827_root_address_inst: Block -- 
      signal in_aggregated_sig: std_logic_vector(6 downto 0);
      signal out_aggregated_sig: std_logic_vector(6 downto 0);
      --
    begin -- 
      ptr_deref_827_root_address_inst_ack_0 <= ptr_deref_827_root_address_inst_req_0;
      in_aggregated_sig <= ptr_deref_827_resized_base_address;
      out_aggregated_sig <= in_aggregated_sig;
      ptr_deref_827_root_address <= out_aggregated_sig(6 downto 0);
      --
    end Block;
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_398_branch_req_0," req0 do_while_stmt_398_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_398_branch_ack_0," ack0 do_while_stmt_398_branch");
    LogCPEvent(clk, reset, global_clock_cycle_count,do_while_stmt_398_branch_ack_1," ack1 do_while_stmt_398_branch");
    do_while_stmt_398_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= unary_844_wire;
      branch_instance: BranchBase -- 
        generic map( condition_width => 1)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_398_branch_req_0,
          ack0 => do_while_stmt_398_branch_ack_0,
          ack1 => do_while_stmt_398_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_410_inst_req_0,binary_410_inst_ack_0,binary_410_inst_req_1,binary_410_inst_ack_1,sl_one,"binary_410_inst",false,indvar_400 & type_cast_409_wire_constant,
    false,tmp2_411);
    -- shared split operator group (0) : binary_410_inst 
    ApIntMul_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_400;
      tmp2_411 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_410_inst_req_0;
      reqR(0) <= binary_410_inst_req_1;
      binary_410_inst_ack_0 <= ackL(0); 
      binary_410_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntMul",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_416_inst_req_0,binary_416_inst_ack_0,binary_416_inst_req_1,binary_416_inst_ack_1,sl_one,"binary_416_inst",false,tmp2_411 & type_cast_415_wire_constant,
    false,tmp3_417);
    -- shared split operator group (1) : binary_416_inst 
    ApIntAdd_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp3_417 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_416_inst_req_0;
      reqR(0) <= binary_416_inst_req_1;
      binary_416_inst_ack_0 <= ackL(0); 
      binary_416_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000111",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_437_inst_req_0,binary_437_inst_ack_0,binary_437_inst_req_1,binary_437_inst_ack_1,sl_one,"binary_437_inst",false,tmp2_411 & type_cast_436_wire_constant,
    false,tmp13_438);
    -- shared split operator group (2) : binary_437_inst 
    ApIntAdd_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp13_438 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_437_inst_req_0;
      reqR(0) <= binary_437_inst_req_1;
      binary_437_inst_ack_0 <= ackL(0); 
      binary_437_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000110",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_458_inst_req_0,binary_458_inst_ack_0,binary_458_inst_req_1,binary_458_inst_ack_1,sl_one,"binary_458_inst",false,tmp2_411 & type_cast_457_wire_constant,
    false,tmp25_459);
    -- shared split operator group (3) : binary_458_inst 
    ApIntAdd_group_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp25_459 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_458_inst_req_0;
      reqR(0) <= binary_458_inst_req_1;
      binary_458_inst_ack_0 <= ackL(0); 
      binary_458_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000101",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_479_inst_req_0,binary_479_inst_ack_0,binary_479_inst_req_1,binary_479_inst_ack_1,sl_one,"binary_479_inst",false,tmp2_411 & type_cast_478_wire_constant,
    false,tmp34_480);
    -- shared split operator group (4) : binary_479_inst 
    ApIntAdd_group_4: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp34_480 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_479_inst_req_0;
      reqR(0) <= binary_479_inst_req_1;
      binary_479_inst_ack_0 <= ackL(0); 
      binary_479_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000100",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_500_inst_req_0,binary_500_inst_ack_0,binary_500_inst_req_1,binary_500_inst_ack_1,sl_one,"binary_500_inst",false,tmp2_411 & type_cast_499_wire_constant,
    false,tmp38_501);
    -- shared split operator group (5) : binary_500_inst 
    ApIntAdd_group_5: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp38_501 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_500_inst_req_0;
      reqR(0) <= binary_500_inst_req_1;
      binary_500_inst_ack_0 <= ackL(0); 
      binary_500_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000011",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_521_inst_req_0,binary_521_inst_ack_0,binary_521_inst_req_1,binary_521_inst_ack_1,sl_one,"binary_521_inst",false,tmp2_411 & type_cast_520_wire_constant,
    false,tmp42_522);
    -- shared split operator group (6) : binary_521_inst 
    ApIntAdd_group_6: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp42_522 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_521_inst_req_0;
      reqR(0) <= binary_521_inst_req_1;
      binary_521_inst_ack_0 <= ackL(0); 
      binary_521_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000010",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_542_inst_req_0,binary_542_inst_ack_0,binary_542_inst_req_1,binary_542_inst_ack_1,sl_one,"binary_542_inst",false,tmp2_411 & type_cast_541_wire_constant,
    false,tmp46_543);
    -- shared split operator group (7) : binary_542_inst 
    ApIntAdd_group_7: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= tmp2_411;
      tmp46_543 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_542_inst_req_0;
      reqR(0) <= binary_542_inst_req_1;
      binary_542_inst_ack_0 <= ackL(0); 
      binary_542_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_663_inst_req_0,binary_663_inst_ack_0,binary_663_inst_req_1,binary_663_inst_ack_1,sl_one,"binary_663_inst",false,iNsTr_20_655 & iNsTr_21_659,
    false,iNsTr_22_664);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_676_inst_req_0,binary_676_inst_ack_0,binary_676_inst_req_1,binary_676_inst_ack_1,sl_one,"binary_676_inst",false,iNsTr_23_668 & iNsTr_24_672,
    false,iNsTr_25_677);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_650_inst_req_0,binary_650_inst_ack_0,binary_650_inst_req_1,binary_650_inst_ack_1,sl_one,"binary_650_inst",false,iNsTr_17_642 & iNsTr_18_646,
    false,iNsTr_19_651);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_637_inst_req_0,binary_637_inst_ack_0,binary_637_inst_req_1,binary_637_inst_ack_1,sl_one,"binary_637_inst",false,iNsTr_14_629 & iNsTr_15_633,
    false,iNsTr_16_638);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_624_inst_req_0,binary_624_inst_ack_0,binary_624_inst_req_1,binary_624_inst_ack_1,sl_one,"binary_624_inst",false,iNsTr_11_616 & iNsTr_12_620,
    false,iNsTr_13_625);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_611_inst_req_0,binary_611_inst_ack_0,binary_611_inst_req_1,binary_611_inst_ack_1,sl_one,"binary_611_inst",false,iNsTr_8_603 & iNsTr_9_607,
    false,iNsTr_10_612);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_598_inst_req_0,binary_598_inst_ack_0,binary_598_inst_req_1,binary_598_inst_ack_1,sl_one,"binary_598_inst",false,iNsTr_5_590 & iNsTr_6_594,
    false,iNsTr_7_599);
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_585_inst_req_0,binary_585_inst_ack_0,binary_585_inst_req_1,binary_585_inst_ack_1,sl_one,"binary_585_inst",false,iNsTr_2_577 & iNsTr_3_581,
    false,iNsTr_4_586);
    -- shared split operator group (8) : binary_663_inst binary_676_inst binary_650_inst binary_637_inst binary_624_inst binary_611_inst binary_598_inst binary_585_inst 
    ApFloatAdd_group_8: Block -- 
      signal data_in: std_logic_vector(511 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      data_in <= iNsTr_20_655 & iNsTr_21_659 & iNsTr_23_668 & iNsTr_24_672 & iNsTr_17_642 & iNsTr_18_646 & iNsTr_14_629 & iNsTr_15_633 & iNsTr_11_616 & iNsTr_12_620 & iNsTr_8_603 & iNsTr_9_607 & iNsTr_5_590 & iNsTr_6_594 & iNsTr_2_577 & iNsTr_3_581;
      iNsTr_22_664 <= data_out(255 downto 224);
      iNsTr_25_677 <= data_out(223 downto 192);
      iNsTr_19_651 <= data_out(191 downto 160);
      iNsTr_16_638 <= data_out(159 downto 128);
      iNsTr_13_625 <= data_out(127 downto 96);
      iNsTr_10_612 <= data_out(95 downto 64);
      iNsTr_7_599 <= data_out(63 downto 32);
      iNsTr_4_586 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      reqL_unguarded(7) <= binary_663_inst_req_0;
      reqL_unguarded(6) <= binary_676_inst_req_0;
      reqL_unguarded(5) <= binary_650_inst_req_0;
      reqL_unguarded(4) <= binary_637_inst_req_0;
      reqL_unguarded(3) <= binary_624_inst_req_0;
      reqL_unguarded(2) <= binary_611_inst_req_0;
      reqL_unguarded(1) <= binary_598_inst_req_0;
      reqL_unguarded(0) <= binary_585_inst_req_0;
      binary_663_inst_ack_0 <= ackL_unguarded(7);
      binary_676_inst_ack_0 <= ackL_unguarded(6);
      binary_650_inst_ack_0 <= ackL_unguarded(5);
      binary_637_inst_ack_0 <= ackL_unguarded(4);
      binary_624_inst_ack_0 <= ackL_unguarded(3);
      binary_611_inst_ack_0 <= ackL_unguarded(2);
      binary_598_inst_ack_0 <= ackL_unguarded(1);
      binary_585_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= binary_663_inst_req_1;
      reqR_unguarded(6) <= binary_676_inst_req_1;
      reqR_unguarded(5) <= binary_650_inst_req_1;
      reqR_unguarded(4) <= binary_637_inst_req_1;
      reqR_unguarded(3) <= binary_624_inst_req_1;
      reqR_unguarded(2) <= binary_611_inst_req_1;
      reqR_unguarded(1) <= binary_598_inst_req_1;
      reqR_unguarded(0) <= binary_585_inst_req_1;
      binary_663_inst_ack_1 <= ackR_unguarded(7);
      binary_676_inst_ack_1 <= ackR_unguarded(6);
      binary_650_inst_ack_1 <= ackR_unguarded(5);
      binary_637_inst_ack_1 <= ackR_unguarded(4);
      binary_624_inst_ack_1 <= ackR_unguarded(3);
      binary_611_inst_ack_1 <= ackR_unguarded(2);
      binary_598_inst_ack_1 <= ackR_unguarded(1);
      binary_585_inst_ack_1 <= ackR_unguarded(0);
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      PipedFpOp: PipelinedFPOperator -- 
        generic map( -- 
          operator_id => "ApFloatAdd",
          exponent_width => 8,
          fraction_width => 23, 
          no_arbitration => false,
          num_reqs => 8 -- 
        )
        port map ( reqL => reqL , ackL => ackL, reqR => reqR, ackR => ackR, dataL => data_in, dataR => data_out, clk => clk, reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_834_inst_req_0,binary_834_inst_ack_0,binary_834_inst_req_1,binary_834_inst_ack_1,sl_one,"binary_834_inst",false,indvar_400 & type_cast_833_wire_constant,
    false,indvarx_xnext_835);
    -- shared split operator group (9) : binary_834_inst 
    ApIntAdd_group_9: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvar_400;
      indvarx_xnext_835 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_834_inst_req_0;
      reqR(0) <= binary_834_inst_req_1;
      binary_834_inst_ack_0 <= ackL(0); 
      binary_834_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 9
    LogSplitOperator(clk,reset,global_clock_cycle_count,binary_840_inst_req_0,binary_840_inst_ack_0,binary_840_inst_req_1,binary_840_inst_ack_1,sl_one,"binary_840_inst",false,indvarx_xnext_835 & type_cast_839_wire_constant,
    false,exitcond1_841);
    -- shared split operator group (10) : binary_840_inst 
    ApIntEq_group_10: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= indvarx_xnext_835;
      exitcond1_841 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= binary_840_inst_req_0;
      reqR(0) <= binary_840_inst_req_1;
      binary_840_inst_ack_0 <= ackL(0); 
      binary_840_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000001000",
          constant_width => 32,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    LogSplitOperator(clk,reset,global_clock_cycle_count,unary_844_inst_req_0,unary_844_inst_ack_0,unary_844_inst_req_1,unary_844_inst_ack_1,sl_one,"unary_844_inst",false,exitcond1_841,
    false,unary_844_wire);
    -- shared split operator group (11) : unary_844_inst 
    ApIntNot_group_11: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      -- 
    begin -- 
      data_in <= exitcond1_841;
      unary_844_wire <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL(0) <= unary_844_inst_req_0;
      reqR(0) <= unary_844_inst_req_1;
      unary_844_inst_ack_0 <= ackL(0); 
      unary_844_inst_ack_1 <= ackR(0); 
      UnsharedOperator: UnsharedOperatorBase -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_667_load_0_req_0,ptr_deref_667_load_0_ack_0,ptr_deref_667_load_0_req_1,ptr_deref_667_load_0_ack_1,sl_one,"ptr_deref_667_load_0",false,ptr_deref_667_word_address_0,
    false,ptr_deref_667_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_576_load_0_req_0,ptr_deref_576_load_0_ack_0,ptr_deref_576_load_0_req_1,ptr_deref_576_load_0_ack_1,sl_one,"ptr_deref_576_load_0",false,ptr_deref_576_word_address_0,
    false,ptr_deref_576_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_589_load_0_req_0,ptr_deref_589_load_0_ack_0,ptr_deref_589_load_0_req_1,ptr_deref_589_load_0_ack_1,sl_one,"ptr_deref_589_load_0",false,ptr_deref_589_word_address_0,
    false,ptr_deref_589_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_602_load_0_req_0,ptr_deref_602_load_0_ack_0,ptr_deref_602_load_0_req_1,ptr_deref_602_load_0_ack_1,sl_one,"ptr_deref_602_load_0",false,ptr_deref_602_word_address_0,
    false,ptr_deref_602_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_615_load_0_req_0,ptr_deref_615_load_0_ack_0,ptr_deref_615_load_0_req_1,ptr_deref_615_load_0_ack_1,sl_one,"ptr_deref_615_load_0",false,ptr_deref_615_word_address_0,
    false,ptr_deref_615_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_628_load_0_req_0,ptr_deref_628_load_0_ack_0,ptr_deref_628_load_0_req_1,ptr_deref_628_load_0_ack_1,sl_one,"ptr_deref_628_load_0",false,ptr_deref_628_word_address_0,
    false,ptr_deref_628_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_641_load_0_req_0,ptr_deref_641_load_0_ack_0,ptr_deref_641_load_0_req_1,ptr_deref_641_load_0_ack_1,sl_one,"ptr_deref_641_load_0",false,ptr_deref_641_word_address_0,
    false,ptr_deref_641_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_654_load_0_req_0,ptr_deref_654_load_0_ack_0,ptr_deref_654_load_0_req_1,ptr_deref_654_load_0_ack_1,sl_one,"ptr_deref_654_load_0",false,ptr_deref_654_word_address_0,
    false,ptr_deref_654_data_0);
    -- shared load operator group (0) : ptr_deref_667_load_0 ptr_deref_576_load_0 ptr_deref_589_load_0 ptr_deref_602_load_0 ptr_deref_615_load_0 ptr_deref_628_load_0 ptr_deref_641_load_0 ptr_deref_654_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_667_load_0_req_0,
        ptr_deref_667_load_0_ack_0,
        ptr_deref_667_load_0_req_1,
        ptr_deref_667_load_0_ack_1,
        "ptr_deref_667_load_0",
        "memory_space_0" ,
        ptr_deref_667_data_0,
        ptr_deref_667_word_address_0,
        "ptr_deref_667_data_0",
        "ptr_deref_667_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_576_load_0_req_0,
        ptr_deref_576_load_0_ack_0,
        ptr_deref_576_load_0_req_1,
        ptr_deref_576_load_0_ack_1,
        "ptr_deref_576_load_0",
        "memory_space_0" ,
        ptr_deref_576_data_0,
        ptr_deref_576_word_address_0,
        "ptr_deref_576_data_0",
        "ptr_deref_576_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_589_load_0_req_0,
        ptr_deref_589_load_0_ack_0,
        ptr_deref_589_load_0_req_1,
        ptr_deref_589_load_0_ack_1,
        "ptr_deref_589_load_0",
        "memory_space_0" ,
        ptr_deref_589_data_0,
        ptr_deref_589_word_address_0,
        "ptr_deref_589_data_0",
        "ptr_deref_589_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_602_load_0_req_0,
        ptr_deref_602_load_0_ack_0,
        ptr_deref_602_load_0_req_1,
        ptr_deref_602_load_0_ack_1,
        "ptr_deref_602_load_0",
        "memory_space_0" ,
        ptr_deref_602_data_0,
        ptr_deref_602_word_address_0,
        "ptr_deref_602_data_0",
        "ptr_deref_602_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_615_load_0_req_0,
        ptr_deref_615_load_0_ack_0,
        ptr_deref_615_load_0_req_1,
        ptr_deref_615_load_0_ack_1,
        "ptr_deref_615_load_0",
        "memory_space_0" ,
        ptr_deref_615_data_0,
        ptr_deref_615_word_address_0,
        "ptr_deref_615_data_0",
        "ptr_deref_615_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_628_load_0_req_0,
        ptr_deref_628_load_0_ack_0,
        ptr_deref_628_load_0_req_1,
        ptr_deref_628_load_0_ack_1,
        "ptr_deref_628_load_0",
        "memory_space_0" ,
        ptr_deref_628_data_0,
        ptr_deref_628_word_address_0,
        "ptr_deref_628_data_0",
        "ptr_deref_628_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_641_load_0_req_0,
        ptr_deref_641_load_0_ack_0,
        ptr_deref_641_load_0_req_1,
        ptr_deref_641_load_0_ack_1,
        "ptr_deref_641_load_0",
        "memory_space_0" ,
        ptr_deref_641_data_0,
        ptr_deref_641_word_address_0,
        "ptr_deref_641_data_0",
        "ptr_deref_641_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_654_load_0_req_0,
        ptr_deref_654_load_0_ack_0,
        ptr_deref_654_load_0_req_1,
        ptr_deref_654_load_0_ack_1,
        "ptr_deref_654_load_0",
        "memory_space_0" ,
        ptr_deref_654_data_0,
        ptr_deref_654_word_address_0,
        "ptr_deref_654_data_0",
        "ptr_deref_654_word_address_0" -- 
      );
      reqL_unguarded(7) <= ptr_deref_667_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_576_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_589_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_602_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_615_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_628_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_641_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_654_load_0_req_0;
      ptr_deref_667_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_576_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_589_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_602_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_615_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_628_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_641_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_654_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_667_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_576_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_589_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_602_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_615_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_628_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_641_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_654_load_0_req_1;
      ptr_deref_667_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_576_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_589_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_602_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_615_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_628_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_641_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_654_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_667_word_address_0 & ptr_deref_576_word_address_0 & ptr_deref_589_word_address_0 & ptr_deref_602_word_address_0 & ptr_deref_615_word_address_0 & ptr_deref_628_word_address_0 & ptr_deref_641_word_address_0 & ptr_deref_654_word_address_0;
      ptr_deref_667_data_0 <= data_out(255 downto 224);
      ptr_deref_576_data_0 <= data_out(223 downto 192);
      ptr_deref_589_data_0 <= data_out(191 downto 160);
      ptr_deref_602_data_0 <= data_out(159 downto 128);
      ptr_deref_615_data_0 <= data_out(127 downto 96);
      ptr_deref_628_data_0 <= data_out(95 downto 64);
      ptr_deref_641_data_0 <= data_out(63 downto 32);
      ptr_deref_654_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_0_lr_req(0),
          mack => memory_space_0_lr_ack(0),
          maddr => memory_space_0_lr_addr(6 downto 0),
          mtag => memory_space_0_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 8,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_0_lc_req(0),
          mack => memory_space_0_lc_ack(0),
          mdata => memory_space_0_lc_data(31 downto 0),
          mtag => memory_space_0_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_658_load_0_req_0,ptr_deref_658_load_0_ack_0,ptr_deref_658_load_0_req_1,ptr_deref_658_load_0_ack_1,sl_one,"ptr_deref_658_load_0",false,ptr_deref_658_word_address_0,
    false,ptr_deref_658_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_671_load_0_req_0,ptr_deref_671_load_0_ack_0,ptr_deref_671_load_0_req_1,ptr_deref_671_load_0_ack_1,sl_one,"ptr_deref_671_load_0",false,ptr_deref_671_word_address_0,
    false,ptr_deref_671_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_580_load_0_req_0,ptr_deref_580_load_0_ack_0,ptr_deref_580_load_0_req_1,ptr_deref_580_load_0_ack_1,sl_one,"ptr_deref_580_load_0",false,ptr_deref_580_word_address_0,
    false,ptr_deref_580_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_593_load_0_req_0,ptr_deref_593_load_0_ack_0,ptr_deref_593_load_0_req_1,ptr_deref_593_load_0_ack_1,sl_one,"ptr_deref_593_load_0",false,ptr_deref_593_word_address_0,
    false,ptr_deref_593_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_606_load_0_req_0,ptr_deref_606_load_0_ack_0,ptr_deref_606_load_0_req_1,ptr_deref_606_load_0_ack_1,sl_one,"ptr_deref_606_load_0",false,ptr_deref_606_word_address_0,
    false,ptr_deref_606_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_619_load_0_req_0,ptr_deref_619_load_0_ack_0,ptr_deref_619_load_0_req_1,ptr_deref_619_load_0_ack_1,sl_one,"ptr_deref_619_load_0",false,ptr_deref_619_word_address_0,
    false,ptr_deref_619_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_632_load_0_req_0,ptr_deref_632_load_0_ack_0,ptr_deref_632_load_0_req_1,ptr_deref_632_load_0_ack_1,sl_one,"ptr_deref_632_load_0",false,ptr_deref_632_word_address_0,
    false,ptr_deref_632_data_0);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_645_load_0_req_0,ptr_deref_645_load_0_ack_0,ptr_deref_645_load_0_req_1,ptr_deref_645_load_0_ack_1,sl_one,"ptr_deref_645_load_0",false,ptr_deref_645_word_address_0,
    false,ptr_deref_645_data_0);
    -- shared load operator group (1) : ptr_deref_658_load_0 ptr_deref_671_load_0 ptr_deref_580_load_0 ptr_deref_593_load_0 ptr_deref_606_load_0 ptr_deref_619_load_0 ptr_deref_632_load_0 ptr_deref_645_load_0 
    LoadGroup1: Block -- 
      signal data_in: std_logic_vector(55 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      -- logging on!
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_658_load_0_req_0,
        ptr_deref_658_load_0_ack_0,
        ptr_deref_658_load_0_req_1,
        ptr_deref_658_load_0_ack_1,
        "ptr_deref_658_load_0",
        "memory_space_1" ,
        ptr_deref_658_data_0,
        ptr_deref_658_word_address_0,
        "ptr_deref_658_data_0",
        "ptr_deref_658_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_671_load_0_req_0,
        ptr_deref_671_load_0_ack_0,
        ptr_deref_671_load_0_req_1,
        ptr_deref_671_load_0_ack_1,
        "ptr_deref_671_load_0",
        "memory_space_1" ,
        ptr_deref_671_data_0,
        ptr_deref_671_word_address_0,
        "ptr_deref_671_data_0",
        "ptr_deref_671_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_580_load_0_req_0,
        ptr_deref_580_load_0_ack_0,
        ptr_deref_580_load_0_req_1,
        ptr_deref_580_load_0_ack_1,
        "ptr_deref_580_load_0",
        "memory_space_1" ,
        ptr_deref_580_data_0,
        ptr_deref_580_word_address_0,
        "ptr_deref_580_data_0",
        "ptr_deref_580_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_593_load_0_req_0,
        ptr_deref_593_load_0_ack_0,
        ptr_deref_593_load_0_req_1,
        ptr_deref_593_load_0_ack_1,
        "ptr_deref_593_load_0",
        "memory_space_1" ,
        ptr_deref_593_data_0,
        ptr_deref_593_word_address_0,
        "ptr_deref_593_data_0",
        "ptr_deref_593_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_606_load_0_req_0,
        ptr_deref_606_load_0_ack_0,
        ptr_deref_606_load_0_req_1,
        ptr_deref_606_load_0_ack_1,
        "ptr_deref_606_load_0",
        "memory_space_1" ,
        ptr_deref_606_data_0,
        ptr_deref_606_word_address_0,
        "ptr_deref_606_data_0",
        "ptr_deref_606_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_619_load_0_req_0,
        ptr_deref_619_load_0_ack_0,
        ptr_deref_619_load_0_req_1,
        ptr_deref_619_load_0_ack_1,
        "ptr_deref_619_load_0",
        "memory_space_1" ,
        ptr_deref_619_data_0,
        ptr_deref_619_word_address_0,
        "ptr_deref_619_data_0",
        "ptr_deref_619_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_632_load_0_req_0,
        ptr_deref_632_load_0_ack_0,
        ptr_deref_632_load_0_req_1,
        ptr_deref_632_load_0_ack_1,
        "ptr_deref_632_load_0",
        "memory_space_1" ,
        ptr_deref_632_data_0,
        ptr_deref_632_word_address_0,
        "ptr_deref_632_data_0",
        "ptr_deref_632_word_address_0" -- 
      );
      LogMemRead(clk, reset, global_clock_cycle_count,-- 
        ptr_deref_645_load_0_req_0,
        ptr_deref_645_load_0_ack_0,
        ptr_deref_645_load_0_req_1,
        ptr_deref_645_load_0_ack_1,
        "ptr_deref_645_load_0",
        "memory_space_1" ,
        ptr_deref_645_data_0,
        ptr_deref_645_word_address_0,
        "ptr_deref_645_data_0",
        "ptr_deref_645_word_address_0" -- 
      );
      reqL_unguarded(7) <= ptr_deref_658_load_0_req_0;
      reqL_unguarded(6) <= ptr_deref_671_load_0_req_0;
      reqL_unguarded(5) <= ptr_deref_580_load_0_req_0;
      reqL_unguarded(4) <= ptr_deref_593_load_0_req_0;
      reqL_unguarded(3) <= ptr_deref_606_load_0_req_0;
      reqL_unguarded(2) <= ptr_deref_619_load_0_req_0;
      reqL_unguarded(1) <= ptr_deref_632_load_0_req_0;
      reqL_unguarded(0) <= ptr_deref_645_load_0_req_0;
      ptr_deref_658_load_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_671_load_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_580_load_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_593_load_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_606_load_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_619_load_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_632_load_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_645_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_658_load_0_req_1;
      reqR_unguarded(6) <= ptr_deref_671_load_0_req_1;
      reqR_unguarded(5) <= ptr_deref_580_load_0_req_1;
      reqR_unguarded(4) <= ptr_deref_593_load_0_req_1;
      reqR_unguarded(3) <= ptr_deref_606_load_0_req_1;
      reqR_unguarded(2) <= ptr_deref_619_load_0_req_1;
      reqR_unguarded(1) <= ptr_deref_632_load_0_req_1;
      reqR_unguarded(0) <= ptr_deref_645_load_0_req_1;
      ptr_deref_658_load_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_671_load_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_580_load_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_593_load_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_606_load_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_619_load_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_632_load_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_645_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      data_in <= ptr_deref_658_word_address_0 & ptr_deref_671_word_address_0 & ptr_deref_580_word_address_0 & ptr_deref_593_word_address_0 & ptr_deref_606_word_address_0 & ptr_deref_619_word_address_0 & ptr_deref_632_word_address_0 & ptr_deref_645_word_address_0;
      ptr_deref_658_data_0 <= data_out(255 downto 224);
      ptr_deref_671_data_0 <= data_out(223 downto 192);
      ptr_deref_580_data_0 <= data_out(191 downto 160);
      ptr_deref_593_data_0 <= data_out(159 downto 128);
      ptr_deref_606_data_0 <= data_out(127 downto 96);
      ptr_deref_619_data_0 <= data_out(95 downto 64);
      ptr_deref_632_data_0 <= data_out(63 downto 32);
      ptr_deref_645_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqShared -- 
        generic map (addr_width => 7,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_1_lr_req(0),
          mack => memory_space_1_lr_ack(0),
          maddr => memory_space_1_lr_addr(6 downto 0),
          mtag => memory_space_1_lr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( data_width => 32,  num_reqs => 8,  tag_length => 4,  no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_1_lc_req(0),
          mack => memory_space_1_lc_ack(0),
          mdata => memory_space_1_lc_data(31 downto 0),
          mtag => memory_space_1_lc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 1
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_713_store_0_req_0,ptr_deref_713_store_0_ack_0,ptr_deref_713_store_0_req_1,ptr_deref_713_store_0_ack_1,sl_one,"ptr_deref_713_store_0",false,ptr_deref_713_word_address_0 & ptr_deref_713_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_827_store_0_req_0,ptr_deref_827_store_0_ack_0,ptr_deref_827_store_0_req_1,ptr_deref_827_store_0_ack_1,sl_one,"ptr_deref_827_store_0",false,ptr_deref_827_word_address_0 & ptr_deref_827_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_732_store_0_req_0,ptr_deref_732_store_0_ack_0,ptr_deref_732_store_0_req_1,ptr_deref_732_store_0_ack_1,sl_one,"ptr_deref_732_store_0",false,ptr_deref_732_word_address_0 & ptr_deref_732_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_770_store_0_req_0,ptr_deref_770_store_0_ack_0,ptr_deref_770_store_0_req_1,ptr_deref_770_store_0_ack_1,sl_one,"ptr_deref_770_store_0",false,ptr_deref_770_word_address_0 & ptr_deref_770_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_694_store_0_req_0,ptr_deref_694_store_0_ack_0,ptr_deref_694_store_0_req_1,ptr_deref_694_store_0_ack_1,sl_one,"ptr_deref_694_store_0",false,ptr_deref_694_word_address_0 & ptr_deref_694_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_751_store_0_req_0,ptr_deref_751_store_0_ack_0,ptr_deref_751_store_0_req_1,ptr_deref_751_store_0_ack_1,sl_one,"ptr_deref_751_store_0",false,ptr_deref_751_word_address_0 & ptr_deref_751_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_789_store_0_req_0,ptr_deref_789_store_0_ack_0,ptr_deref_789_store_0_req_1,ptr_deref_789_store_0_ack_1,sl_one,"ptr_deref_789_store_0",false,ptr_deref_789_word_address_0 & ptr_deref_789_data_0,
    true, slv_zero);
    LogSplitOperator(clk,reset,global_clock_cycle_count,ptr_deref_808_store_0_req_0,ptr_deref_808_store_0_ack_0,ptr_deref_808_store_0_req_1,ptr_deref_808_store_0_ack_1,sl_one,"ptr_deref_808_store_0",false,ptr_deref_808_word_address_0 & ptr_deref_808_data_0,
    true, slv_zero);
    -- logging on!
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_713_store_0_req_0,
      ptr_deref_713_store_0_ack_0,
      ptr_deref_713_store_0_req_1,
      ptr_deref_713_store_0_ack_1,
      "ptr_deref_713_store_0",
      "memory_space_2" ,
      ptr_deref_713_data_0,
      ptr_deref_713_word_address_0,
      "ptr_deref_713_data_0",
      "ptr_deref_713_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_827_store_0_req_0,
      ptr_deref_827_store_0_ack_0,
      ptr_deref_827_store_0_req_1,
      ptr_deref_827_store_0_ack_1,
      "ptr_deref_827_store_0",
      "memory_space_2" ,
      ptr_deref_827_data_0,
      ptr_deref_827_word_address_0,
      "ptr_deref_827_data_0",
      "ptr_deref_827_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_732_store_0_req_0,
      ptr_deref_732_store_0_ack_0,
      ptr_deref_732_store_0_req_1,
      ptr_deref_732_store_0_ack_1,
      "ptr_deref_732_store_0",
      "memory_space_2" ,
      ptr_deref_732_data_0,
      ptr_deref_732_word_address_0,
      "ptr_deref_732_data_0",
      "ptr_deref_732_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_770_store_0_req_0,
      ptr_deref_770_store_0_ack_0,
      ptr_deref_770_store_0_req_1,
      ptr_deref_770_store_0_ack_1,
      "ptr_deref_770_store_0",
      "memory_space_2" ,
      ptr_deref_770_data_0,
      ptr_deref_770_word_address_0,
      "ptr_deref_770_data_0",
      "ptr_deref_770_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_694_store_0_req_0,
      ptr_deref_694_store_0_ack_0,
      ptr_deref_694_store_0_req_1,
      ptr_deref_694_store_0_ack_1,
      "ptr_deref_694_store_0",
      "memory_space_2" ,
      ptr_deref_694_data_0,
      ptr_deref_694_word_address_0,
      "ptr_deref_694_data_0",
      "ptr_deref_694_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_751_store_0_req_0,
      ptr_deref_751_store_0_ack_0,
      ptr_deref_751_store_0_req_1,
      ptr_deref_751_store_0_ack_1,
      "ptr_deref_751_store_0",
      "memory_space_2" ,
      ptr_deref_751_data_0,
      ptr_deref_751_word_address_0,
      "ptr_deref_751_data_0",
      "ptr_deref_751_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_789_store_0_req_0,
      ptr_deref_789_store_0_ack_0,
      ptr_deref_789_store_0_req_1,
      ptr_deref_789_store_0_ack_1,
      "ptr_deref_789_store_0",
      "memory_space_2" ,
      ptr_deref_789_data_0,
      ptr_deref_789_word_address_0,
      "ptr_deref_789_data_0",
      "ptr_deref_789_word_address_0" -- 
    );
    LogMemWrite(clk, reset,global_clock_cycle_count,  -- 
      ptr_deref_808_store_0_req_0,
      ptr_deref_808_store_0_ack_0,
      ptr_deref_808_store_0_req_1,
      ptr_deref_808_store_0_ack_1,
      "ptr_deref_808_store_0",
      "memory_space_2" ,
      ptr_deref_808_data_0,
      ptr_deref_808_word_address_0,
      "ptr_deref_808_data_0",
      "ptr_deref_808_word_address_0" -- 
    );
    -- shared store operator group (0) : ptr_deref_713_store_0 ptr_deref_827_store_0 ptr_deref_732_store_0 ptr_deref_770_store_0 ptr_deref_694_store_0 ptr_deref_751_store_0 ptr_deref_789_store_0 ptr_deref_808_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(55 downto 0);
      signal data_in: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 7 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 7 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 7 downto 0);
      signal guard_vector : std_logic_vector( 7 downto 0);
      -- 
    begin -- 
      reqL_unguarded(7) <= ptr_deref_713_store_0_req_0;
      reqL_unguarded(6) <= ptr_deref_827_store_0_req_0;
      reqL_unguarded(5) <= ptr_deref_732_store_0_req_0;
      reqL_unguarded(4) <= ptr_deref_770_store_0_req_0;
      reqL_unguarded(3) <= ptr_deref_694_store_0_req_0;
      reqL_unguarded(2) <= ptr_deref_751_store_0_req_0;
      reqL_unguarded(1) <= ptr_deref_789_store_0_req_0;
      reqL_unguarded(0) <= ptr_deref_808_store_0_req_0;
      ptr_deref_713_store_0_ack_0 <= ackL_unguarded(7);
      ptr_deref_827_store_0_ack_0 <= ackL_unguarded(6);
      ptr_deref_732_store_0_ack_0 <= ackL_unguarded(5);
      ptr_deref_770_store_0_ack_0 <= ackL_unguarded(4);
      ptr_deref_694_store_0_ack_0 <= ackL_unguarded(3);
      ptr_deref_751_store_0_ack_0 <= ackL_unguarded(2);
      ptr_deref_789_store_0_ack_0 <= ackL_unguarded(1);
      ptr_deref_808_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(7) <= ptr_deref_713_store_0_req_1;
      reqR_unguarded(6) <= ptr_deref_827_store_0_req_1;
      reqR_unguarded(5) <= ptr_deref_732_store_0_req_1;
      reqR_unguarded(4) <= ptr_deref_770_store_0_req_1;
      reqR_unguarded(3) <= ptr_deref_694_store_0_req_1;
      reqR_unguarded(2) <= ptr_deref_751_store_0_req_1;
      reqR_unguarded(1) <= ptr_deref_789_store_0_req_1;
      reqR_unguarded(0) <= ptr_deref_808_store_0_req_1;
      ptr_deref_713_store_0_ack_1 <= ackR_unguarded(7);
      ptr_deref_827_store_0_ack_1 <= ackR_unguarded(6);
      ptr_deref_732_store_0_ack_1 <= ackR_unguarded(5);
      ptr_deref_770_store_0_ack_1 <= ackR_unguarded(4);
      ptr_deref_694_store_0_ack_1 <= ackR_unguarded(3);
      ptr_deref_751_store_0_ack_1 <= ackR_unguarded(2);
      ptr_deref_789_store_0_ack_1 <= ackR_unguarded(1);
      ptr_deref_808_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      guard_vector(4)  <=  '1';
      guard_vector(5)  <=  '1';
      guard_vector(6)  <=  '1';
      guard_vector(7)  <=  '1';
      gI0: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqL_unguarded,
        ackL => ackL_unguarded,
        reqR => reqL_unregulated,
        ackR => ackL_unregulated,
        guards => guard_vector); -- 
      accessRegulator_0: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessRegulator_1: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessRegulator_2: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessRegulator_3: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessRegulator_4: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      accessRegulator_5: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      accessRegulator_6: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(6), -- 
          ack => ackL_unregulated(6),
          regulated_req => reqL(6),
          regulated_ack => ackL(6),
          release_req => reqR(6),
          release_ack => ackR(6),
          clk => clk, reset => reset); -- 
      accessRegulator_7: access_regulator_base generic map (num_slots => 1) -- 
        port map (req => reqL_unregulated(7), -- 
          ack => ackL_unregulated(7),
          regulated_req => reqL(7),
          regulated_ack => ackL(7),
          release_req => reqR(7),
          release_ack => ackR(7),
          clk => clk, reset => reset); -- 
      gI1: GuardInterface generic map(nreqs => 8) -- 
        port map(reqL => reqR_unguarded,
        ackL => ackR_unguarded,
        reqR => reqR,
        ackR => ackR,
        guards => guard_vector); -- 
      addr_in <= ptr_deref_713_word_address_0 & ptr_deref_827_word_address_0 & ptr_deref_732_word_address_0 & ptr_deref_770_word_address_0 & ptr_deref_694_word_address_0 & ptr_deref_751_word_address_0 & ptr_deref_789_word_address_0 & ptr_deref_808_word_address_0;
      data_in <= ptr_deref_713_data_0 & ptr_deref_827_data_0 & ptr_deref_732_data_0 & ptr_deref_770_data_0 & ptr_deref_694_data_0 & ptr_deref_751_data_0 & ptr_deref_789_data_0 & ptr_deref_808_data_0;
      StoreReq: StoreReqShared -- 
        generic map ( addr_width => 7,
        data_width => 32,
        num_reqs => 8,
        tag_length => 4,
        time_stamp_width => 3,
        min_clock_period => false,
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(6 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(6 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          num_reqs => 8,
          tag_length => 4 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(3 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end Default;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library work;
use work.ahir_system_global_package.all;
entity ahir_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    in_data_pipe_pipe_write_data: in std_logic_vector(31 downto 0);
    in_data_pipe_pipe_write_req : in std_logic_vector(0 downto 0);
    in_data_pipe_pipe_write_ack : out std_logic_vector(0 downto 0);
    out_data_pipe_pipe_read_data: out std_logic_vector(31 downto 0);
    out_data_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    out_data_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture Default of ahir_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  signal memory_space_0_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_0_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_0_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_0_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_0_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_0_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_0_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_0_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_0_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_0_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_0_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_1
  signal memory_space_1_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_1_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_1_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_1_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_1_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_1_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_1_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_1_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_1_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_1_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_1_sc_tag :  std_logic_vector(3 downto 0);
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(31 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(3 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(0 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(0 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(6 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(31 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(6 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(0 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(0 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(3 downto 0);
  -- declarations related to module vectorSum
  component vectorSum is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_1_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_1_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_1_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_sc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_0_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_0_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_sc_tag :  in  std_logic_vector(3 downto 0);
      in_data_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      in_data_pipe_pipe_read_data : in   std_logic_vector(31 downto 0);
      out_data_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
      out_data_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
      out_data_pipe_pipe_write_data : out  std_logic_vector(31 downto 0);
      x_vectorSum_x_call_reqs : out  std_logic_vector(0 downto 0);
      x_vectorSum_x_call_acks : in   std_logic_vector(0 downto 0);
      x_vectorSum_x_call_tag  :  out  std_logic_vector(0 downto 0);
      x_vectorSum_x_return_reqs : out  std_logic_vector(0 downto 0);
      x_vectorSum_x_return_acks : in   std_logic_vector(0 downto 0);
      x_vectorSum_x_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module vectorSum
  signal vectorSum_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal vectorSum_tag_out   : std_logic_vector(1 downto 0);
  signal vectorSum_start_req : std_logic;
  signal vectorSum_start_ack : std_logic;
  signal vectorSum_fin_req   : std_logic;
  signal vectorSum_fin_ack : std_logic;
  -- declarations related to module x_vectorSum_x
  component x_vectorSum_x is -- 
    generic (tag_length : integer); 
    port ( -- 
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      memory_space_1_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_1_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_1_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_1_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_1_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_1_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_0_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lr_addr : out  std_logic_vector(6 downto 0);
      memory_space_0_lr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_0_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_0_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_0_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_0_lc_tag :  in  std_logic_vector(3 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(6 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(6 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
    -- 
  end component;
  -- argument signals for module x_vectorSum_x
  signal x_vectorSum_x_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal x_vectorSum_x_tag_out   : std_logic_vector(1 downto 0);
  signal x_vectorSum_x_start_req : std_logic;
  signal x_vectorSum_x_start_ack : std_logic;
  signal x_vectorSum_x_fin_req   : std_logic;
  signal x_vectorSum_x_fin_ack : std_logic;
  -- caller side aggregated signals for module x_vectorSum_x
  signal x_vectorSum_x_call_reqs: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_call_acks: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_reqs: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_acks: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_call_tag: std_logic_vector(0 downto 0);
  signal x_vectorSum_x_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe in_data_pipe
  signal in_data_pipe_pipe_read_data: std_logic_vector(31 downto 0);
  signal in_data_pipe_pipe_read_req: std_logic_vector(0 downto 0);
  signal in_data_pipe_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe out_data_pipe
  signal out_data_pipe_pipe_write_data: std_logic_vector(31 downto 0);
  signal out_data_pipe_pipe_write_req: std_logic_vector(0 downto 0);
  signal out_data_pipe_pipe_write_ack: std_logic_vector(0 downto 0);
  -- 
begin -- 
  -- module vectorSum
  vectorSum_instance:vectorSum-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => vectorSum_start_req,
      start_ack => vectorSum_start_ack,
      fin_req => vectorSum_fin_req,
      fin_ack => vectorSum_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(6 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(6 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(3 downto 0),
      memory_space_0_sr_req => memory_space_0_sr_req(0 downto 0),
      memory_space_0_sr_ack => memory_space_0_sr_ack(0 downto 0),
      memory_space_0_sr_addr => memory_space_0_sr_addr(6 downto 0),
      memory_space_0_sr_data => memory_space_0_sr_data(31 downto 0),
      memory_space_0_sr_tag => memory_space_0_sr_tag(6 downto 0),
      memory_space_0_sc_req => memory_space_0_sc_req(0 downto 0),
      memory_space_0_sc_ack => memory_space_0_sc_ack(0 downto 0),
      memory_space_0_sc_tag => memory_space_0_sc_tag(3 downto 0),
      memory_space_1_sr_req => memory_space_1_sr_req(0 downto 0),
      memory_space_1_sr_ack => memory_space_1_sr_ack(0 downto 0),
      memory_space_1_sr_addr => memory_space_1_sr_addr(6 downto 0),
      memory_space_1_sr_data => memory_space_1_sr_data(31 downto 0),
      memory_space_1_sr_tag => memory_space_1_sr_tag(6 downto 0),
      memory_space_1_sc_req => memory_space_1_sc_req(0 downto 0),
      memory_space_1_sc_ack => memory_space_1_sc_ack(0 downto 0),
      memory_space_1_sc_tag => memory_space_1_sc_tag(3 downto 0),
      in_data_pipe_pipe_read_req => in_data_pipe_pipe_read_req(0 downto 0),
      in_data_pipe_pipe_read_ack => in_data_pipe_pipe_read_ack(0 downto 0),
      in_data_pipe_pipe_read_data => in_data_pipe_pipe_read_data(31 downto 0),
      out_data_pipe_pipe_write_req => out_data_pipe_pipe_write_req(0 downto 0),
      out_data_pipe_pipe_write_ack => out_data_pipe_pipe_write_ack(0 downto 0),
      out_data_pipe_pipe_write_data => out_data_pipe_pipe_write_data(31 downto 0),
      x_vectorSum_x_call_reqs => x_vectorSum_x_call_reqs(0 downto 0),
      x_vectorSum_x_call_acks => x_vectorSum_x_call_acks(0 downto 0),
      x_vectorSum_x_call_tag => x_vectorSum_x_call_tag(0 downto 0),
      x_vectorSum_x_return_reqs => x_vectorSum_x_return_reqs(0 downto 0),
      x_vectorSum_x_return_acks => x_vectorSum_x_return_acks(0 downto 0),
      x_vectorSum_x_return_tag => x_vectorSum_x_return_tag(0 downto 0),
      tag_in => vectorSum_tag_in,
      tag_out => vectorSum_tag_out-- 
    ); -- 
  -- module will be run forever 
  vectorSum_tag_in <= (others => '0');
  vectorSum_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => vectorSum_start_req, start_ack => vectorSum_start_ack,  fin_req => vectorSum_fin_req,  fin_ack => vectorSum_fin_ack);
  -- module x_vectorSum_x
  -- call arbiter for module x_vectorSum_x
  x_vectorSum_x_arbiter: SplitCallArbiterNoInargsNoOutargs -- 
    generic map( --
      num_reqs => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => x_vectorSum_x_call_reqs,
      call_acks => x_vectorSum_x_call_acks,
      return_reqs => x_vectorSum_x_return_reqs,
      return_acks => x_vectorSum_x_return_acks,
      call_tag  => x_vectorSum_x_call_tag,
      return_tag  => x_vectorSum_x_return_tag,
      call_mtag => x_vectorSum_x_tag_in,
      return_mtag => x_vectorSum_x_tag_out,
      call_mreq => x_vectorSum_x_start_req,
      call_mack => x_vectorSum_x_start_ack,
      return_mreq => x_vectorSum_x_fin_req,
      return_mack => x_vectorSum_x_fin_ack,
      clk => clk, 
      reset => reset --
    ); --
  x_vectorSum_x_instance:x_vectorSum_x-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => x_vectorSum_x_start_req,
      start_ack => x_vectorSum_x_start_ack,
      fin_req => x_vectorSum_x_fin_req,
      fin_ack => x_vectorSum_x_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_0_lr_req => memory_space_0_lr_req(0 downto 0),
      memory_space_0_lr_ack => memory_space_0_lr_ack(0 downto 0),
      memory_space_0_lr_addr => memory_space_0_lr_addr(6 downto 0),
      memory_space_0_lr_tag => memory_space_0_lr_tag(6 downto 0),
      memory_space_0_lc_req => memory_space_0_lc_req(0 downto 0),
      memory_space_0_lc_ack => memory_space_0_lc_ack(0 downto 0),
      memory_space_0_lc_data => memory_space_0_lc_data(31 downto 0),
      memory_space_0_lc_tag => memory_space_0_lc_tag(3 downto 0),
      memory_space_1_lr_req => memory_space_1_lr_req(0 downto 0),
      memory_space_1_lr_ack => memory_space_1_lr_ack(0 downto 0),
      memory_space_1_lr_addr => memory_space_1_lr_addr(6 downto 0),
      memory_space_1_lr_tag => memory_space_1_lr_tag(6 downto 0),
      memory_space_1_lc_req => memory_space_1_lc_req(0 downto 0),
      memory_space_1_lc_ack => memory_space_1_lc_ack(0 downto 0),
      memory_space_1_lc_data => memory_space_1_lc_data(31 downto 0),
      memory_space_1_lc_tag => memory_space_1_lc_tag(3 downto 0),
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(6 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(6 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(3 downto 0),
      tag_in => x_vectorSum_x_tag_in,
      tag_out => x_vectorSum_x_tag_out-- 
    ); -- 
  in_data_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => in_data_pipe_pipe_read_req,
      read_ack => in_data_pipe_pipe_read_ack,
      read_data => in_data_pipe_pipe_read_data,
      write_req => in_data_pipe_pipe_write_req,
      write_ack => in_data_pipe_pipe_write_ack,
      write_data => in_data_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  out_data_pipe_Pipe: PipeBase -- 
    generic map( -- 
      num_reads => 1,
      num_writes => 1,
      data_width => 32,
      lifo_mode => false,
      depth => 1 --
    )
    port map( -- 
      read_req => out_data_pipe_pipe_read_req,
      read_ack => out_data_pipe_pipe_read_ack,
      read_data => out_data_pipe_pipe_read_data,
      write_req => out_data_pipe_pipe_write_req,
      write_ack => out_data_pipe_pipe_write_ack,
      write_data => out_data_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MemorySpace_memory_space_0: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_0_lr_addr,
      lr_req_in => memory_space_0_lr_req,
      lr_ack_out => memory_space_0_lr_ack,
      lr_tag_in => memory_space_0_lr_tag,
      lc_req_in => memory_space_0_lc_req,
      lc_ack_out => memory_space_0_lc_ack,
      lc_data_out => memory_space_0_lc_data,
      lc_tag_out => memory_space_0_lc_tag,
      sr_addr_in => memory_space_0_sr_addr,
      sr_data_in => memory_space_0_sr_data,
      sr_req_in => memory_space_0_sr_req,
      sr_ack_out => memory_space_0_sr_ack,
      sr_tag_in => memory_space_0_sr_tag,
      sc_req_in=> memory_space_0_sc_req,
      sc_ack_out => memory_space_0_sc_ack,
      sc_tag_out => memory_space_0_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_1: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_1_lr_addr,
      lr_req_in => memory_space_1_lr_req,
      lr_ack_out => memory_space_1_lr_ack,
      lr_tag_in => memory_space_1_lr_tag,
      lc_req_in => memory_space_1_lc_req,
      lc_ack_out => memory_space_1_lc_ack,
      lc_data_out => memory_space_1_lc_data,
      lc_tag_out => memory_space_1_lc_tag,
      sr_addr_in => memory_space_1_sr_addr,
      sr_data_in => memory_space_1_sr_data,
      sr_req_in => memory_space_1_sr_req,
      sr_ack_out => memory_space_1_sr_ack,
      sr_tag_in => memory_space_1_sr_tag,
      sc_req_in=> memory_space_1_sc_req,
      sc_ack_out => memory_space_1_sc_ack,
      sc_tag_out => memory_space_1_sc_tag,
      clock => clk,
      reset => reset); -- 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      num_loads => 1,
      num_stores => 1,
      addr_width => 7,
      data_width => 32,
      tag_width => 4,
      time_stamp_width => 3,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 7,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end Default;
