-- $Header: /devl/xcs/repo/env/Databases/CAEInterfaces/vhdsclibs/data/simprims/fuji/VITAL/X_USR_ACCESSE2.vhd,v 1.2 2010/05/27 23:13:00 yanx Exp $
-------------------------------------------------------
--  Copyright (c) 2009 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : X_USR_ACCESSE2.vhd
-- \   \  /  \      
--  \__ \/\__ \                   
--                                 
--  Generated by    : /home/chen/xfoundry/HEAD/env/Databases/CAEInterfaces/LibraryWriters/bin/ltw.pl
--  Revision: 1.0
-------------------------------------------------------

----- CELL X_USR_ACCESSE2 -----

library IEEE;
use IEEE.STD_LOGIC_arith.all;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

library simprim;
use simprim.VCOMPONENTS.all;
use simprim.VPACKAGE.all;

  entity X_USR_ACCESSE2 is
    generic (
      TimingChecksOn : boolean := TRUE;
      InstancePath   : string  := "*";
      Xon            : boolean := TRUE;
      MsgOn          : boolean := FALSE;
      LOC            : string  := "UNPLACED"
    );

    port (
      CFGCLK               : out std_ulogic;
      DATA                 : out std_logic_vector(31 downto 0);
      DATAVALID            : out std_ulogic
    );
    attribute VITAL_LEVEL0 of X_USR_ACCESSE2 :     entity is true;
  end X_USR_ACCESSE2;

  architecture X_USR_ACCESSE2_V of X_USR_ACCESSE2 is
    TYPE VitalTimingDataArrayType IS ARRAY (NATURAL RANGE <>) OF VitalTimingDataType;
    
    constant IN_DELAY : time := 0 ps;
    constant OUT_DELAY : time := 0 ps;
    constant INCLK_DELAY : time := 0 ps;
    constant OUTCLK_DELAY : time := 0 ps;

    function SUL_TO_STR (sul : std_ulogic)
    return string is
    begin
      if sul = '0' then
        return "0";
      else
        return "1";
      end if;
    end SUL_TO_STR;

    function boolean_to_string(bool: boolean)
    return string is
    begin
      if bool then
        return "TRUE";
      else
        return "FALSE";
      end if;
    end boolean_to_string;

    function getstrlength(in_vec : std_logic_vector)
    return integer is
      variable string_length : integer;
    begin
      if ((in_vec'length mod 4) = 0) then
        string_length := in_vec'length/4;
      elsif ((in_vec'length mod 4) > 0) then
        string_length := in_vec'length/4 + 1;
      end if;
      return string_length;
    end getstrlength;

    signal CFGCLK_out : std_ulogic;
    signal DATAVALID_out : std_ulogic;
    signal DATA_out : std_logic_vector(31 downto 0);
    
    signal CFGCLK_outdelay : std_ulogic;
    signal DATAVALID_outdelay : std_ulogic;
    signal DATA_outdelay : std_logic_vector(31 downto 0);
    
    begin
    
    WireDelay : block
    begin
    end block;
    
    SignalDelay : block
    begin
    end block;
    CFGCLK_out <= CFGCLK_outdelay after OUT_DELAY;
    DATAVALID_out <= DATAVALID_outdelay after OUT_DELAY;
    DATA_out <= DATA_outdelay after OUT_DELAY;
    
    
    TIMING : process

      begin

      wait on
        CFGCLK_out,
        DATAVALID_out,
        DATA_out;
    end process TIMING;
    CFGCLK <= CFGCLK_out;
    DATA <= DATA_out;
    DATAVALID <= DATAVALID_out;
  end X_USR_ACCESSE2_V;
