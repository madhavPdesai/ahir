library work;
use work.cpath_components.all;

entity start_cp is
  port (

    ip    : in bit_vector(27 downto 1);
    op    : out bit_vector(32 downto 1) := (others => '0');
    reset : in bit;
    clk   : in bit);
end start_cp;

architecture behavioral of start_cp is

  signal place_1_tip : bit_vector(0 downto 0);
  signal place_1_rst : bit_vector(0 downto 0);
  signal place_1_top : bit;
  signal place_10_tip : bit_vector(0 downto 0);
  signal place_10_rst : bit_vector(0 downto 0);
  signal place_10_top : bit;
  signal place_12_tip : bit_vector(0 downto 0);
  signal place_12_rst : bit_vector(0 downto 0);
  signal place_12_top : bit;
  signal place_13_tip : bit_vector(0 downto 0);
  signal place_13_rst : bit_vector(0 downto 0);
  signal place_13_top : bit;
  signal place_14_tip : bit_vector(0 downto 0);
  signal place_14_rst : bit_vector(0 downto 0);
  signal place_14_top : bit;
  signal place_15_tip : bit_vector(0 downto 0);
  signal place_15_rst : bit_vector(0 downto 0);
  signal place_15_top : bit;
  signal place_16_tip : bit_vector(0 downto 0);
  signal place_16_rst : bit_vector(0 downto 0);
  signal place_16_top : bit;
  signal place_18_tip : bit_vector(0 downto 0);
  signal place_18_rst : bit_vector(0 downto 0);
  signal place_18_top : bit;
  signal place_19_tip : bit_vector(0 downto 0);
  signal place_19_rst : bit_vector(1 downto 0);
  signal place_19_top : bit;
  signal place_2_tip : bit_vector(0 downto 0);
  signal place_2_rst : bit_vector(0 downto 0);
  signal place_2_top : bit;
  signal place_20_tip : bit_vector(0 downto 0);
  signal place_20_rst : bit_vector(0 downto 0);
  signal place_20_top : bit;
  signal place_21_tip : bit_vector(1 downto 0);
  signal place_21_rst : bit_vector(0 downto 0);
  signal place_21_top : bit;
  signal place_22_tip : bit_vector(0 downto 0);
  signal place_22_rst : bit_vector(0 downto 0);
  signal place_22_top : bit;
  signal place_23_tip : bit_vector(0 downto 0);
  signal place_23_rst : bit_vector(0 downto 0);
  signal place_23_top : bit;
  signal place_24_tip : bit_vector(0 downto 0);
  signal place_24_rst : bit_vector(0 downto 0);
  signal place_24_top : bit;
  signal place_25_tip : bit_vector(0 downto 0);
  signal place_25_rst : bit_vector(0 downto 0);
  signal place_25_top : bit;
  signal place_26_tip : bit_vector(1 downto 0);
  signal place_26_rst : bit_vector(0 downto 0);
  signal place_26_top : bit;
  signal place_27_tip : bit_vector(0 downto 0);
  signal place_27_rst : bit_vector(0 downto 0);
  signal place_27_top : bit;
  signal place_28_tip : bit_vector(0 downto 0);
  signal place_28_rst : bit_vector(0 downto 0);
  signal place_28_top : bit;
  signal place_29_tip : bit_vector(0 downto 0);
  signal place_29_rst : bit_vector(0 downto 0);
  signal place_29_top : bit;
  signal place_3_tip : bit_vector(0 downto 0);
  signal place_3_rst : bit_vector(0 downto 0);
  signal place_3_top : bit;
  signal place_30_tip : bit_vector(0 downto 0);
  signal place_30_rst : bit_vector(0 downto 0);
  signal place_30_top : bit;
  signal place_31_tip : bit_vector(1 downto 0);
  signal place_31_rst : bit_vector(0 downto 0);
  signal place_31_top : bit;
  signal place_32_tip : bit_vector(0 downto 0);
  signal place_32_rst : bit_vector(0 downto 0);
  signal place_32_top : bit;
  signal place_33_tip : bit_vector(0 downto 0);
  signal place_33_rst : bit_vector(0 downto 0);
  signal place_33_top : bit;
  signal place_34_tip : bit_vector(0 downto 0);
  signal place_34_rst : bit_vector(0 downto 0);
  signal place_34_top : bit;
  signal place_35_tip : bit_vector(0 downto 0);
  signal place_35_rst : bit_vector(0 downto 0);
  signal place_35_top : bit;
  signal place_36_tip : bit_vector(1 downto 0);
  signal place_36_rst : bit_vector(0 downto 0);
  signal place_36_top : bit;
  signal place_37_tip : bit_vector(0 downto 0);
  signal place_37_rst : bit_vector(0 downto 0);
  signal place_37_top : bit;
  signal place_38_tip : bit_vector(0 downto 0);
  signal place_38_rst : bit_vector(0 downto 0);
  signal place_38_top : bit;
  signal place_39_tip : bit_vector(0 downto 0);
  signal place_39_rst : bit_vector(0 downto 0);
  signal place_39_top : bit;
  signal place_40_tip : bit_vector(0 downto 0);
  signal place_40_rst : bit_vector(0 downto 0);
  signal place_40_top : bit;
  signal place_41_tip : bit_vector(0 downto 0);
  signal place_41_rst : bit_vector(0 downto 0);
  signal place_41_top : bit;
  signal place_42_tip : bit_vector(0 downto 0);
  signal place_42_rst : bit_vector(1 downto 0);
  signal place_42_top : bit;
  signal place_43_tip : bit_vector(0 downto 0);
  signal place_43_rst : bit_vector(0 downto 0);
  signal place_43_top : bit;
  signal place_44_tip : bit_vector(1 downto 0);
  signal place_44_rst : bit_vector(0 downto 0);
  signal place_44_top : bit;
  signal place_45_tip : bit_vector(0 downto 0);
  signal place_45_rst : bit_vector(0 downto 0);
  signal place_45_top : bit;
  signal place_46_tip : bit_vector(0 downto 0);
  signal place_46_rst : bit_vector(0 downto 0);
  signal place_46_top : bit;
  signal place_47_tip : bit_vector(0 downto 0);
  signal place_47_rst : bit_vector(0 downto 0);
  signal place_47_top : bit;
  signal place_48_tip : bit_vector(1 downto 0);
  signal place_48_rst : bit_vector(0 downto 0);
  signal place_48_top : bit;
  signal place_49_tip : bit_vector(0 downto 0);
  signal place_49_rst : bit_vector(0 downto 0);
  signal place_49_top : bit;
  signal place_5_tip : bit_vector(0 downto 0);
  signal place_5_rst : bit_vector(0 downto 0);
  signal place_5_top : bit;
  signal place_50_tip : bit_vector(0 downto 0);
  signal place_50_rst : bit_vector(0 downto 0);
  signal place_50_top : bit;
  signal place_51_tip : bit_vector(0 downto 0);
  signal place_51_rst : bit_vector(0 downto 0);
  signal place_51_top : bit;
  signal place_52_tip : bit_vector(1 downto 0);
  signal place_52_rst : bit_vector(0 downto 0);
  signal place_52_top : bit;
  signal place_53_tip : bit_vector(0 downto 0);
  signal place_53_rst : bit_vector(0 downto 0);
  signal place_53_top : bit;
  signal place_54_tip : bit_vector(0 downto 0);
  signal place_54_rst : bit_vector(0 downto 0);
  signal place_54_top : bit;
  signal place_55_tip : bit_vector(0 downto 0);
  signal place_55_rst : bit_vector(0 downto 0);
  signal place_55_top : bit;
  signal place_56_tip : bit_vector(0 downto 0);
  signal place_56_rst : bit_vector(0 downto 0);
  signal place_56_top : bit;
  signal place_57_tip : bit_vector(0 downto 0);
  signal place_57_rst : bit_vector(0 downto 0);
  signal place_57_top : bit;
  signal place_58_tip : bit_vector(0 downto 0);
  signal place_58_rst : bit_vector(0 downto 0);
  signal place_58_top : bit;
  signal place_59_tip : bit_vector(0 downto 0);
  signal place_59_rst : bit_vector(0 downto 0);
  signal place_59_top : bit;
  signal place_60_tip : bit_vector(0 downto 0);
  signal place_60_rst : bit_vector(0 downto 0);
  signal place_60_top : bit;
  signal place_61_tip : bit_vector(0 downto 0);
  signal place_61_rst : bit_vector(0 downto 0);
  signal place_61_top : bit;
  signal place_62_tip : bit_vector(0 downto 0);
  signal place_62_rst : bit_vector(0 downto 0);
  signal place_62_top : bit;
  signal place_63_tip : bit_vector(0 downto 0);
  signal place_63_rst : bit_vector(0 downto 0);
  signal place_63_top : bit;
  signal place_64_tip : bit_vector(0 downto 0);
  signal place_64_rst : bit_vector(0 downto 0);
  signal place_64_top : bit;
  signal place_65_tip : bit_vector(0 downto 0);
  signal place_65_rst : bit_vector(0 downto 0);
  signal place_65_top : bit;
  signal place_66_tip : bit_vector(0 downto 0);
  signal place_66_rst : bit_vector(1 downto 0);
  signal place_66_top : bit;
  signal place_68_tip : bit_vector(0 downto 0);
  signal place_68_rst : bit_vector(0 downto 0);
  signal place_68_top : bit;
  signal place_69_tip : bit_vector(1 downto 0);
  signal place_69_rst : bit_vector(0 downto 0);
  signal place_69_top : bit;
  signal place_7_tip : bit_vector(0 downto 0);
  signal place_7_rst : bit_vector(0 downto 0);
  signal place_7_top : bit;
  signal place_70_tip : bit_vector(0 downto 0);
  signal place_70_rst : bit_vector(0 downto 0);
  signal place_70_top : bit;
  signal place_72_tip : bit_vector(0 downto 0);
  signal place_72_rst : bit_vector(0 downto 0);
  signal place_72_top : bit;
  signal place_73_tip : bit_vector(0 downto 0);
  signal place_73_rst : bit_vector(0 downto 0);
  signal place_73_top : bit;
  signal place_74_tip : bit_vector(0 downto 0);
  signal place_74_rst : bit_vector(1 downto 0);
  signal place_74_top : bit;
  signal place_76_tip : bit_vector(0 downto 0);
  signal place_76_rst : bit_vector(0 downto 0);
  signal place_76_top : bit;
  signal place_77_tip : bit_vector(1 downto 0);
  signal place_77_rst : bit_vector(0 downto 0);
  signal place_77_top : bit;
  signal place_78_tip : bit_vector(0 downto 0);
  signal place_78_rst : bit_vector(0 downto 0);
  signal place_78_top : bit;
  signal place_80_tip : bit_vector(0 downto 0);
  signal place_80_rst : bit_vector(0 downto 0);
  signal place_80_top : bit;
  signal place_81_tip : bit_vector(0 downto 0);
  signal place_81_rst : bit_vector(0 downto 0);
  signal place_81_top : bit;
  signal place_82_tip : bit_vector(0 downto 0);
  signal place_82_rst : bit_vector(0 downto 0);
  signal place_82_top : bit;
  signal place_83_tip : bit_vector(0 downto 0);
  signal place_83_rst : bit_vector(0 downto 0);
  signal place_83_top : bit;
  signal place_84_tip : bit_vector(0 downto 0);
  signal place_84_rst : bit_vector(0 downto 0);
  signal place_84_top : bit;

  signal cbr_4_oper_tmp_d_1_d_i_bool_d_req_tip : bit_vector(0 downto 0);
  signal cbr_4_oper_tmp_d_1_d_i_bool_d_req_ge : bit;
  signal cbr_4_oper_tmp_d_1_d_i_bool_d_req_top : bit;
  signal cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip : bit_vector(3 downto 0);
  signal cbr_5_oper_tmp_d_6_d_i_bool_d_req_ge : bit;
  signal cbr_5_oper_tmp_d_6_d_i_bool_d_req_top : bit;
  signal cbr_6_oper_tmp_d_17_d_i_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_6_oper_tmp_d_17_d_i_bool_d_req_ge : bit;
  signal cbr_6_oper_tmp_d_17_d_i_bool_d_req_top : bit;
  signal cbr_7_oper_tmp_d_17_d_i_bool_d_req_tip : bit_vector(1 downto 0);
  signal cbr_7_oper_tmp_d_17_d_i_bool_d_req_ge : bit;
  signal cbr_7_oper_tmp_d_17_d_i_bool_d_req_top : bit;
  signal entry_to_loopentry_d_i_src_tip : bit_vector(0 downto 0);
  signal entry_to_loopentry_d_i_src_ge : bit;
  signal entry_to_loopentry_d_i_src_top : bit;
  signal entry_to_no_exit_d_i_src_tip : bit_vector(0 downto 0);
  signal entry_to_no_exit_d_i_src_ge : bit;
  signal entry_to_no_exit_d_i_src_top : bit;
  signal fin_tip : bit_vector(0 downto 0);
  signal fin_ge : bit;
  signal fin_top : bit;
  signal i_d_0_d_i_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_d_0_mux_1_d_ack_ge : bit;
  signal i_d_0_d_i_d_0_mux_1_d_ack_top : bit;
  signal i_d_0_d_i_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_d_0_mux_1_d_req0_ge : bit;
  signal i_d_0_d_i_d_0_mux_1_d_req0_top : bit;
  signal i_d_0_d_i_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_d_0_mux_1_d_req1_ge : bit;
  signal i_d_0_d_i_d_0_mux_1_d_req1_top : bit;
  signal i_d_0_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_mux_1_d_ack_ge : bit;
  signal i_d_0_d_i_mux_1_d_ack_top : bit;
  signal i_d_0_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_mux_1_d_req0_ge : bit;
  signal i_d_0_d_i_mux_1_d_req0_top : bit;
  signal i_d_0_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal i_d_0_d_i_mux_1_d_req1_ge : bit;
  signal i_d_0_d_i_mux_1_d_req1_top : bit;
  signal init_tip : bit_vector(0 downto 0);
  signal init_ge : bit;
  signal init_top : bit;
  signal llimit_d_1_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal llimit_d_1_d_i_mux_1_d_ack_ge : bit;
  signal llimit_d_1_d_i_mux_1_d_ack_top : bit;
  signal llimit_d_1_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal llimit_d_1_d_i_mux_1_d_req0_ge : bit;
  signal llimit_d_1_d_i_mux_1_d_req0_top : bit;
  signal llimit_d_1_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal llimit_d_1_d_i_mux_1_d_req1_ge : bit;
  signal llimit_d_1_d_i_mux_1_d_req1_top : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_d_0_mux_1_d_ack_ge : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_ack_top : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_d_0_mux_1_d_req0_ge : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_req0_top : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_d_0_mux_1_d_req1_ge : bit;
  signal llimit_d_2_d_i_d_0_mux_1_d_req1_top : bit;
  signal llimit_d_2_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_mux_1_d_ack_ge : bit;
  signal llimit_d_2_d_i_mux_1_d_ack_top : bit;
  signal llimit_d_2_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_mux_1_d_req0_ge : bit;
  signal llimit_d_2_d_i_mux_1_d_req0_top : bit;
  signal llimit_d_2_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal llimit_d_2_d_i_mux_1_d_req1_ge : bit;
  signal llimit_d_2_d_i_mux_1_d_req1_top : bit;
  signal load_number_d_ack_tip : bit_vector(0 downto 0);
  signal load_number_d_ack_ge : bit;
  signal load_number_d_ack_top : bit;
  signal load_number_d_req_tip : bit_vector(0 downto 0);
  signal load_number_d_req_ge : bit;
  signal load_number_d_req_top : bit;
  signal loopentry_d_i_d_entry_tip : bit_vector(0 downto 0);
  signal loopentry_d_i_d_entry_ge : bit;
  signal loopentry_d_i_d_entry_top : bit;
  signal loopentry_d_i_d_pre_tip : bit_vector(3 downto 0);
  signal loopentry_d_i_d_pre_ge : bit;
  signal loopentry_d_i_d_pre_top : bit;
  signal loopentry_d_i_to_no_exit_d_i_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_i_to_no_exit_d_i_src_ge : bit;
  signal loopentry_d_i_to_no_exit_d_i_src_top : bit;
  signal loopentry_d_i_to_sqroot_d_exit_src_tip : bit_vector(0 downto 0);
  signal loopentry_d_i_to_sqroot_d_exit_src_ge : bit;
  signal loopentry_d_i_to_sqroot_d_exit_src_top : bit;
  signal mid_d_0_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal mid_d_0_d_i_mux_1_d_ack_ge : bit;
  signal mid_d_0_d_i_mux_1_d_ack_top : bit;
  signal mid_d_0_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal mid_d_0_d_i_mux_1_d_req0_ge : bit;
  signal mid_d_0_d_i_mux_1_d_req0_top : bit;
  signal mid_d_0_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal mid_d_0_d_i_mux_1_d_req1_ge : bit;
  signal mid_d_0_d_i_mux_1_d_req1_top : bit;
  signal no_exit_d_i_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_d_entry_ge : bit;
  signal no_exit_d_i_d_entry_top : bit;
  signal no_exit_d_i_d_pre_tip : bit_vector(2 downto 0);
  signal no_exit_d_i_d_pre_ge : bit;
  signal no_exit_d_i_d_pre_top : bit;
  signal no_exit_d_i_d_selectcont_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_d_selectcont_d_entry_ge : bit;
  signal no_exit_d_i_d_selectcont_d_entry_top : bit;
  signal no_exit_d_i_d_selectcont_d_selectcont_d_entry_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_d_selectcont_d_selectcont_d_entry_ge : bit;
  signal no_exit_d_i_d_selectcont_d_selectcont_d_entry_top : bit;
  signal no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_tip : bit_vector(1 downto 0);
  signal no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_ge : bit;
  signal no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top : bit;
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_ge : bit;
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_top : bit;
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_ge : bit;
  signal no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_top : bit;
  signal no_exit_d_i_to_no_exit_d_i_d_selectcont_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_to_no_exit_d_i_d_selectcont_src_ge : bit;
  signal no_exit_d_i_to_no_exit_d_i_d_selectcont_src_top : bit;
  signal no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_tip : bit_vector(0 downto 0);
  signal no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_ge : bit;
  signal no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_top : bit;
  signal oper_inc_d_i_int_d_ack_tip : bit_vector(0 downto 0);
  signal oper_inc_d_i_int_d_ack_ge : bit;
  signal oper_inc_d_i_int_d_ack_top : bit;
  signal oper_inc_d_i_int_d_req_tip : bit_vector(0 downto 0);
  signal oper_inc_d_i_int_d_req_ge : bit;
  signal oper_inc_d_i_int_d_req_top : bit;
  signal oper_tmp_d_10_d_i_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_10_d_i_float_d_ack_ge : bit;
  signal oper_tmp_d_10_d_i_float_d_ack_top : bit;
  signal oper_tmp_d_10_d_i_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_10_d_i_float_d_req_ge : bit;
  signal oper_tmp_d_10_d_i_float_d_req_top : bit;
  signal oper_tmp_d_11_d_i_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_i_float_d_ack_ge : bit;
  signal oper_tmp_d_11_d_i_float_d_ack_top : bit;
  signal oper_tmp_d_11_d_i_float_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_11_d_i_float_d_req_ge : bit;
  signal oper_tmp_d_11_d_i_float_d_req_top : bit;
  signal oper_tmp_d_14_d_i_float_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_14_d_i_float_d_ack_ge : bit;
  signal oper_tmp_d_14_d_i_float_d_ack_top : bit;
  signal oper_tmp_d_14_d_i_float_d_req_tip : bit_vector(1 downto 0);
  signal oper_tmp_d_14_d_i_float_d_req_ge : bit;
  signal oper_tmp_d_14_d_i_float_d_req_top : bit;
  signal oper_tmp_d_17_d_i_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_17_d_i_bool_d_ack_ge : bit;
  signal oper_tmp_d_17_d_i_bool_d_ack_top : bit;
  signal oper_tmp_d_17_d_i_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_17_d_i_bool_d_req_ge : bit;
  signal oper_tmp_d_17_d_i_bool_d_req_top : bit;
  signal oper_tmp_d_1_d_i_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1_d_i_bool_d_ack_ge : bit;
  signal oper_tmp_d_1_d_i_bool_d_ack_top : bit;
  signal oper_tmp_d_1_d_i_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_1_d_i_bool_d_req_ge : bit;
  signal oper_tmp_d_1_d_i_bool_d_req_top : bit;
  signal oper_tmp_d_6_d_i_bool_d_ack_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_6_d_i_bool_d_ack_ge : bit;
  signal oper_tmp_d_6_d_i_bool_d_ack_top : bit;
  signal oper_tmp_d_6_d_i_bool_d_req_tip : bit_vector(0 downto 0);
  signal oper_tmp_d_6_d_i_bool_d_req_ge : bit;
  signal oper_tmp_d_6_d_i_bool_d_req_top : bit;
  signal store_location_start_return_d_ack_tip : bit_vector(0 downto 0);
  signal store_location_start_return_d_ack_ge : bit;
  signal store_location_start_return_d_ack_top : bit;
  signal store_location_start_return_d_req_tip : bit_vector(0 downto 0);
  signal store_location_start_return_d_req_ge : bit;
  signal store_location_start_return_d_req_top : bit;
  signal ulimit_d_1_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ulimit_d_1_d_i_mux_1_d_ack_ge : bit;
  signal ulimit_d_1_d_i_mux_1_d_ack_top : bit;
  signal ulimit_d_1_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ulimit_d_1_d_i_mux_1_d_req0_ge : bit;
  signal ulimit_d_1_d_i_mux_1_d_req0_top : bit;
  signal ulimit_d_1_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ulimit_d_1_d_i_mux_1_d_req1_ge : bit;
  signal ulimit_d_1_d_i_mux_1_d_req1_top : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_d_0_mux_1_d_ack_ge : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_ack_top : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_d_0_mux_1_d_req0_ge : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_req0_top : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_d_0_mux_1_d_req1_ge : bit;
  signal ulimit_d_2_d_i_d_0_mux_1_d_req1_top : bit;
  signal ulimit_d_2_d_i_mux_1_d_ack_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_mux_1_d_ack_ge : bit;
  signal ulimit_d_2_d_i_mux_1_d_ack_top : bit;
  signal ulimit_d_2_d_i_mux_1_d_req0_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_mux_1_d_req0_ge : bit;
  signal ulimit_d_2_d_i_mux_1_d_req0_top : bit;
  signal ulimit_d_2_d_i_mux_1_d_req1_tip : bit_vector(0 downto 0);
  signal ulimit_d_2_d_i_mux_1_d_req1_ge : bit;
  signal ulimit_d_2_d_i_mux_1_d_req1_top : bit;

begin


  place_1 : place
  generic map(1, 1, '0')
  port map(place_1_tip, place_1_rst, place_1_top, reset, clk);

  place_10 : place
  generic map(1, 1, '0')
  port map(place_10_tip, place_10_rst, place_10_top, reset, clk);

  place_12 : place
  generic map(1, 1, '1')
  port map(place_12_tip, place_12_rst, place_12_top, reset, clk);

  place_13 : place
  generic map(1, 1, '0')
  port map(place_13_tip, place_13_rst, place_13_top, reset, clk);

  place_14 : place
  generic map(1, 1, '0')
  port map(place_14_tip, place_14_rst, place_14_top, reset, clk);

  place_15 : place
  generic map(1, 1, '0')
  port map(place_15_tip, place_15_rst, place_15_top, reset, clk);

  place_16 : place
  generic map(1, 1, '0')
  port map(place_16_tip, place_16_rst, place_16_top, reset, clk);

  place_18 : place
  generic map(1, 1, '0')
  port map(place_18_tip, place_18_rst, place_18_top, reset, clk);

  place_19 : place
  generic map(1, 2, '0')
  port map(place_19_tip, place_19_rst, place_19_top, reset, clk);

  place_2 : place
  generic map(1, 1, '0')
  port map(place_2_tip, place_2_rst, place_2_top, reset, clk);

  place_20 : place
  generic map(1, 1, '0')
  port map(place_20_tip, place_20_rst, place_20_top, reset, clk);

  place_21 : place
  generic map(2, 1, '0')
  port map(place_21_tip, place_21_rst, place_21_top, reset, clk);

  place_22 : place
  generic map(1, 1, '0')
  port map(place_22_tip, place_22_rst, place_22_top, reset, clk);

  place_23 : place
  generic map(1, 1, '0')
  port map(place_23_tip, place_23_rst, place_23_top, reset, clk);

  place_24 : place
  generic map(1, 1, '0')
  port map(place_24_tip, place_24_rst, place_24_top, reset, clk);

  place_25 : place
  generic map(1, 1, '0')
  port map(place_25_tip, place_25_rst, place_25_top, reset, clk);

  place_26 : place
  generic map(2, 1, '0')
  port map(place_26_tip, place_26_rst, place_26_top, reset, clk);

  place_27 : place
  generic map(1, 1, '0')
  port map(place_27_tip, place_27_rst, place_27_top, reset, clk);

  place_28 : place
  generic map(1, 1, '0')
  port map(place_28_tip, place_28_rst, place_28_top, reset, clk);

  place_29 : place
  generic map(1, 1, '0')
  port map(place_29_tip, place_29_rst, place_29_top, reset, clk);

  place_3 : place
  generic map(1, 1, '0')
  port map(place_3_tip, place_3_rst, place_3_top, reset, clk);

  place_30 : place
  generic map(1, 1, '0')
  port map(place_30_tip, place_30_rst, place_30_top, reset, clk);

  place_31 : place
  generic map(2, 1, '0')
  port map(place_31_tip, place_31_rst, place_31_top, reset, clk);

  place_32 : place
  generic map(1, 1, '0')
  port map(place_32_tip, place_32_rst, place_32_top, reset, clk);

  place_33 : place
  generic map(1, 1, '0')
  port map(place_33_tip, place_33_rst, place_33_top, reset, clk);

  place_34 : place
  generic map(1, 1, '0')
  port map(place_34_tip, place_34_rst, place_34_top, reset, clk);

  place_35 : place
  generic map(1, 1, '0')
  port map(place_35_tip, place_35_rst, place_35_top, reset, clk);

  place_36 : place
  generic map(2, 1, '0')
  port map(place_36_tip, place_36_rst, place_36_top, reset, clk);

  place_37 : place
  generic map(1, 1, '0')
  port map(place_37_tip, place_37_rst, place_37_top, reset, clk);

  place_38 : place
  generic map(1, 1, '0')
  port map(place_38_tip, place_38_rst, place_38_top, reset, clk);

  place_39 : place
  generic map(1, 1, '0')
  port map(place_39_tip, place_39_rst, place_39_top, reset, clk);

  place_40 : place
  generic map(1, 1, '0')
  port map(place_40_tip, place_40_rst, place_40_top, reset, clk);

  place_41 : place
  generic map(1, 1, '0')
  port map(place_41_tip, place_41_rst, place_41_top, reset, clk);

  place_42 : place
  generic map(1, 2, '0')
  port map(place_42_tip, place_42_rst, place_42_top, reset, clk);

  place_43 : place
  generic map(1, 1, '0')
  port map(place_43_tip, place_43_rst, place_43_top, reset, clk);

  place_44 : place
  generic map(2, 1, '0')
  port map(place_44_tip, place_44_rst, place_44_top, reset, clk);

  place_45 : place
  generic map(1, 1, '0')
  port map(place_45_tip, place_45_rst, place_45_top, reset, clk);

  place_46 : place
  generic map(1, 1, '0')
  port map(place_46_tip, place_46_rst, place_46_top, reset, clk);

  place_47 : place
  generic map(1, 1, '0')
  port map(place_47_tip, place_47_rst, place_47_top, reset, clk);

  place_48 : place
  generic map(2, 1, '0')
  port map(place_48_tip, place_48_rst, place_48_top, reset, clk);

  place_49 : place
  generic map(1, 1, '0')
  port map(place_49_tip, place_49_rst, place_49_top, reset, clk);

  place_5 : place
  generic map(1, 1, '0')
  port map(place_5_tip, place_5_rst, place_5_top, reset, clk);

  place_50 : place
  generic map(1, 1, '0')
  port map(place_50_tip, place_50_rst, place_50_top, reset, clk);

  place_51 : place
  generic map(1, 1, '0')
  port map(place_51_tip, place_51_rst, place_51_top, reset, clk);

  place_52 : place
  generic map(2, 1, '0')
  port map(place_52_tip, place_52_rst, place_52_top, reset, clk);

  place_53 : place
  generic map(1, 1, '0')
  port map(place_53_tip, place_53_rst, place_53_top, reset, clk);

  place_54 : place
  generic map(1, 1, '0')
  port map(place_54_tip, place_54_rst, place_54_top, reset, clk);

  place_55 : place
  generic map(1, 1, '0')
  port map(place_55_tip, place_55_rst, place_55_top, reset, clk);

  place_56 : place
  generic map(1, 1, '0')
  port map(place_56_tip, place_56_rst, place_56_top, reset, clk);

  place_57 : place
  generic map(1, 1, '0')
  port map(place_57_tip, place_57_rst, place_57_top, reset, clk);

  place_58 : place
  generic map(1, 1, '0')
  port map(place_58_tip, place_58_rst, place_58_top, reset, clk);

  place_59 : place
  generic map(1, 1, '0')
  port map(place_59_tip, place_59_rst, place_59_top, reset, clk);

  place_60 : place
  generic map(1, 1, '0')
  port map(place_60_tip, place_60_rst, place_60_top, reset, clk);

  place_61 : place
  generic map(1, 1, '0')
  port map(place_61_tip, place_61_rst, place_61_top, reset, clk);

  place_62 : place
  generic map(1, 1, '0')
  port map(place_62_tip, place_62_rst, place_62_top, reset, clk);

  place_63 : place
  generic map(1, 1, '0')
  port map(place_63_tip, place_63_rst, place_63_top, reset, clk);

  place_64 : place
  generic map(1, 1, '0')
  port map(place_64_tip, place_64_rst, place_64_top, reset, clk);

  place_65 : place
  generic map(1, 1, '0')
  port map(place_65_tip, place_65_rst, place_65_top, reset, clk);

  place_66 : place
  generic map(1, 2, '0')
  port map(place_66_tip, place_66_rst, place_66_top, reset, clk);

  place_68 : place
  generic map(1, 1, '0')
  port map(place_68_tip, place_68_rst, place_68_top, reset, clk);

  place_69 : place
  generic map(2, 1, '0')
  port map(place_69_tip, place_69_rst, place_69_top, reset, clk);

  place_7 : place
  generic map(1, 1, '0')
  port map(place_7_tip, place_7_rst, place_7_top, reset, clk);

  place_70 : place
  generic map(1, 1, '0')
  port map(place_70_tip, place_70_rst, place_70_top, reset, clk);

  place_72 : place
  generic map(1, 1, '0')
  port map(place_72_tip, place_72_rst, place_72_top, reset, clk);

  place_73 : place
  generic map(1, 1, '0')
  port map(place_73_tip, place_73_rst, place_73_top, reset, clk);

  place_74 : place
  generic map(1, 2, '0')
  port map(place_74_tip, place_74_rst, place_74_top, reset, clk);

  place_76 : place
  generic map(1, 1, '0')
  port map(place_76_tip, place_76_rst, place_76_top, reset, clk);

  place_77 : place
  generic map(2, 1, '0')
  port map(place_77_tip, place_77_rst, place_77_top, reset, clk);

  place_78 : place
  generic map(1, 1, '0')
  port map(place_78_tip, place_78_rst, place_78_top, reset, clk);

  place_80 : place
  generic map(1, 1, '0')
  port map(place_80_tip, place_80_rst, place_80_top, reset, clk);

  place_81 : place
  generic map(1, 1, '0')
  port map(place_81_tip, place_81_rst, place_81_top, reset, clk);

  place_82 : place
  generic map(1, 1, '0')
  port map(place_82_tip, place_82_rst, place_82_top, reset, clk);

  place_83 : place
  generic map(1, 1, '0')
  port map(place_83_tip, place_83_rst, place_83_top, reset, clk);

  place_84 : place
  generic map(1, 1, '0')
  port map(place_84_tip, place_84_rst, place_84_top, reset, clk);


  cbr_4_oper_tmp_d_1_d_i_bool_d_req : transition
  generic map(1)
  port map(cbr_4_oper_tmp_d_1_d_i_bool_d_req_tip, cbr_4_oper_tmp_d_1_d_i_bool_d_req_ge, cbr_4_oper_tmp_d_1_d_i_bool_d_req_top);

  cbr_5_oper_tmp_d_6_d_i_bool_d_req : transition
  generic map(4)
  port map(cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip, cbr_5_oper_tmp_d_6_d_i_bool_d_req_ge, cbr_5_oper_tmp_d_6_d_i_bool_d_req_top);

  cbr_6_oper_tmp_d_17_d_i_bool_d_req : transition
  generic map(2)
  port map(cbr_6_oper_tmp_d_17_d_i_bool_d_req_tip, cbr_6_oper_tmp_d_17_d_i_bool_d_req_ge, cbr_6_oper_tmp_d_17_d_i_bool_d_req_top);

  cbr_7_oper_tmp_d_17_d_i_bool_d_req : transition
  generic map(2)
  port map(cbr_7_oper_tmp_d_17_d_i_bool_d_req_tip, cbr_7_oper_tmp_d_17_d_i_bool_d_req_ge, cbr_7_oper_tmp_d_17_d_i_bool_d_req_top);

  entry_to_loopentry_d_i_src : transition
  generic map(1)
  port map(entry_to_loopentry_d_i_src_tip, entry_to_loopentry_d_i_src_ge, entry_to_loopentry_d_i_src_top);

  entry_to_no_exit_d_i_src : transition
  generic map(1)
  port map(entry_to_no_exit_d_i_src_tip, entry_to_no_exit_d_i_src_ge, entry_to_no_exit_d_i_src_top);

  fin : transition
  generic map(1)
  port map(fin_tip, fin_ge, fin_top);

  i_d_0_d_i_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(i_d_0_d_i_d_0_mux_1_d_ack_tip, i_d_0_d_i_d_0_mux_1_d_ack_ge, i_d_0_d_i_d_0_mux_1_d_ack_top);

  i_d_0_d_i_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(i_d_0_d_i_d_0_mux_1_d_req0_tip, i_d_0_d_i_d_0_mux_1_d_req0_ge, i_d_0_d_i_d_0_mux_1_d_req0_top);

  i_d_0_d_i_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(i_d_0_d_i_d_0_mux_1_d_req1_tip, i_d_0_d_i_d_0_mux_1_d_req1_ge, i_d_0_d_i_d_0_mux_1_d_req1_top);

  i_d_0_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(i_d_0_d_i_mux_1_d_ack_tip, i_d_0_d_i_mux_1_d_ack_ge, i_d_0_d_i_mux_1_d_ack_top);

  i_d_0_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(i_d_0_d_i_mux_1_d_req0_tip, i_d_0_d_i_mux_1_d_req0_ge, i_d_0_d_i_mux_1_d_req0_top);

  i_d_0_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(i_d_0_d_i_mux_1_d_req1_tip, i_d_0_d_i_mux_1_d_req1_ge, i_d_0_d_i_mux_1_d_req1_top);

  init : transition
  generic map(1)
  port map(init_tip, init_ge, init_top);

  llimit_d_1_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(llimit_d_1_d_i_mux_1_d_ack_tip, llimit_d_1_d_i_mux_1_d_ack_ge, llimit_d_1_d_i_mux_1_d_ack_top);

  llimit_d_1_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(llimit_d_1_d_i_mux_1_d_req0_tip, llimit_d_1_d_i_mux_1_d_req0_ge, llimit_d_1_d_i_mux_1_d_req0_top);

  llimit_d_1_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(llimit_d_1_d_i_mux_1_d_req1_tip, llimit_d_1_d_i_mux_1_d_req1_ge, llimit_d_1_d_i_mux_1_d_req1_top);

  llimit_d_2_d_i_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(llimit_d_2_d_i_d_0_mux_1_d_ack_tip, llimit_d_2_d_i_d_0_mux_1_d_ack_ge, llimit_d_2_d_i_d_0_mux_1_d_ack_top);

  llimit_d_2_d_i_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(llimit_d_2_d_i_d_0_mux_1_d_req0_tip, llimit_d_2_d_i_d_0_mux_1_d_req0_ge, llimit_d_2_d_i_d_0_mux_1_d_req0_top);

  llimit_d_2_d_i_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(llimit_d_2_d_i_d_0_mux_1_d_req1_tip, llimit_d_2_d_i_d_0_mux_1_d_req1_ge, llimit_d_2_d_i_d_0_mux_1_d_req1_top);

  llimit_d_2_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(llimit_d_2_d_i_mux_1_d_ack_tip, llimit_d_2_d_i_mux_1_d_ack_ge, llimit_d_2_d_i_mux_1_d_ack_top);

  llimit_d_2_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(llimit_d_2_d_i_mux_1_d_req0_tip, llimit_d_2_d_i_mux_1_d_req0_ge, llimit_d_2_d_i_mux_1_d_req0_top);

  llimit_d_2_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(llimit_d_2_d_i_mux_1_d_req1_tip, llimit_d_2_d_i_mux_1_d_req1_ge, llimit_d_2_d_i_mux_1_d_req1_top);

  load_number_d_ack : transition
  generic map(1)
  port map(load_number_d_ack_tip, load_number_d_ack_ge, load_number_d_ack_top);

  load_number_d_req : transition
  generic map(1)
  port map(load_number_d_req_tip, load_number_d_req_ge, load_number_d_req_top);

  loopentry_d_i_d_entry : transition
  generic map(1)
  port map(loopentry_d_i_d_entry_tip, loopentry_d_i_d_entry_ge, loopentry_d_i_d_entry_top);

  loopentry_d_i_d_pre : transition
  generic map(4)
  port map(loopentry_d_i_d_pre_tip, loopentry_d_i_d_pre_ge, loopentry_d_i_d_pre_top);

  loopentry_d_i_to_no_exit_d_i_src : transition
  generic map(1)
  port map(loopentry_d_i_to_no_exit_d_i_src_tip, loopentry_d_i_to_no_exit_d_i_src_ge, loopentry_d_i_to_no_exit_d_i_src_top);

  loopentry_d_i_to_sqroot_d_exit_src : transition
  generic map(1)
  port map(loopentry_d_i_to_sqroot_d_exit_src_tip, loopentry_d_i_to_sqroot_d_exit_src_ge, loopentry_d_i_to_sqroot_d_exit_src_top);

  mid_d_0_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(mid_d_0_d_i_mux_1_d_ack_tip, mid_d_0_d_i_mux_1_d_ack_ge, mid_d_0_d_i_mux_1_d_ack_top);

  mid_d_0_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(mid_d_0_d_i_mux_1_d_req0_tip, mid_d_0_d_i_mux_1_d_req0_ge, mid_d_0_d_i_mux_1_d_req0_top);

  mid_d_0_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(mid_d_0_d_i_mux_1_d_req1_tip, mid_d_0_d_i_mux_1_d_req1_ge, mid_d_0_d_i_mux_1_d_req1_top);

  no_exit_d_i_d_entry : transition
  generic map(1)
  port map(no_exit_d_i_d_entry_tip, no_exit_d_i_d_entry_ge, no_exit_d_i_d_entry_top);

  no_exit_d_i_d_pre : transition
  generic map(3)
  port map(no_exit_d_i_d_pre_tip, no_exit_d_i_d_pre_ge, no_exit_d_i_d_pre_top);

  no_exit_d_i_d_selectcont_d_entry : transition
  generic map(1)
  port map(no_exit_d_i_d_selectcont_d_entry_tip, no_exit_d_i_d_selectcont_d_entry_ge, no_exit_d_i_d_selectcont_d_entry_top);

  no_exit_d_i_d_selectcont_d_selectcont_d_entry : transition
  generic map(1)
  port map(no_exit_d_i_d_selectcont_d_selectcont_d_entry_tip, no_exit_d_i_d_selectcont_d_selectcont_d_entry_ge, no_exit_d_i_d_selectcont_d_selectcont_d_entry_top);

  no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src : transition
  generic map(2)
  port map(no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_tip, no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_ge, no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top);

  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src : transition
  generic map(1)
  port map(no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_tip, no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_ge, no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_top);

  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src : transition
  generic map(1)
  port map(no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_tip, no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_ge, no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_top);

  no_exit_d_i_to_no_exit_d_i_d_selectcont_src : transition
  generic map(1)
  port map(no_exit_d_i_to_no_exit_d_i_d_selectcont_src_tip, no_exit_d_i_to_no_exit_d_i_d_selectcont_src_ge, no_exit_d_i_to_no_exit_d_i_d_selectcont_src_top);

  no_exit_d_i_to_no_exit_d_i_d_selecttrue_src : transition
  generic map(1)
  port map(no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_tip, no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_ge, no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_top);

  oper_inc_d_i_int_d_ack : transition
  generic map(1)
  port map(oper_inc_d_i_int_d_ack_tip, oper_inc_d_i_int_d_ack_ge, oper_inc_d_i_int_d_ack_top);

  oper_inc_d_i_int_d_req : transition
  generic map(1)
  port map(oper_inc_d_i_int_d_req_tip, oper_inc_d_i_int_d_req_ge, oper_inc_d_i_int_d_req_top);

  oper_tmp_d_10_d_i_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_10_d_i_float_d_ack_tip, oper_tmp_d_10_d_i_float_d_ack_ge, oper_tmp_d_10_d_i_float_d_ack_top);

  oper_tmp_d_10_d_i_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_10_d_i_float_d_req_tip, oper_tmp_d_10_d_i_float_d_req_ge, oper_tmp_d_10_d_i_float_d_req_top);

  oper_tmp_d_11_d_i_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_11_d_i_float_d_ack_tip, oper_tmp_d_11_d_i_float_d_ack_ge, oper_tmp_d_11_d_i_float_d_ack_top);

  oper_tmp_d_11_d_i_float_d_req : transition
  generic map(1)
  port map(oper_tmp_d_11_d_i_float_d_req_tip, oper_tmp_d_11_d_i_float_d_req_ge, oper_tmp_d_11_d_i_float_d_req_top);

  oper_tmp_d_14_d_i_float_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_14_d_i_float_d_ack_tip, oper_tmp_d_14_d_i_float_d_ack_ge, oper_tmp_d_14_d_i_float_d_ack_top);

  oper_tmp_d_14_d_i_float_d_req : transition
  generic map(2)
  port map(oper_tmp_d_14_d_i_float_d_req_tip, oper_tmp_d_14_d_i_float_d_req_ge, oper_tmp_d_14_d_i_float_d_req_top);

  oper_tmp_d_17_d_i_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_17_d_i_bool_d_ack_tip, oper_tmp_d_17_d_i_bool_d_ack_ge, oper_tmp_d_17_d_i_bool_d_ack_top);

  oper_tmp_d_17_d_i_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_17_d_i_bool_d_req_tip, oper_tmp_d_17_d_i_bool_d_req_ge, oper_tmp_d_17_d_i_bool_d_req_top);

  oper_tmp_d_1_d_i_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_1_d_i_bool_d_ack_tip, oper_tmp_d_1_d_i_bool_d_ack_ge, oper_tmp_d_1_d_i_bool_d_ack_top);

  oper_tmp_d_1_d_i_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_1_d_i_bool_d_req_tip, oper_tmp_d_1_d_i_bool_d_req_ge, oper_tmp_d_1_d_i_bool_d_req_top);

  oper_tmp_d_6_d_i_bool_d_ack : transition
  generic map(1)
  port map(oper_tmp_d_6_d_i_bool_d_ack_tip, oper_tmp_d_6_d_i_bool_d_ack_ge, oper_tmp_d_6_d_i_bool_d_ack_top);

  oper_tmp_d_6_d_i_bool_d_req : transition
  generic map(1)
  port map(oper_tmp_d_6_d_i_bool_d_req_tip, oper_tmp_d_6_d_i_bool_d_req_ge, oper_tmp_d_6_d_i_bool_d_req_top);

  store_location_start_return_d_ack : transition
  generic map(1)
  port map(store_location_start_return_d_ack_tip, store_location_start_return_d_ack_ge, store_location_start_return_d_ack_top);

  store_location_start_return_d_req : transition
  generic map(1)
  port map(store_location_start_return_d_req_tip, store_location_start_return_d_req_ge, store_location_start_return_d_req_top);

  ulimit_d_1_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(ulimit_d_1_d_i_mux_1_d_ack_tip, ulimit_d_1_d_i_mux_1_d_ack_ge, ulimit_d_1_d_i_mux_1_d_ack_top);

  ulimit_d_1_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(ulimit_d_1_d_i_mux_1_d_req0_tip, ulimit_d_1_d_i_mux_1_d_req0_ge, ulimit_d_1_d_i_mux_1_d_req0_top);

  ulimit_d_1_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(ulimit_d_1_d_i_mux_1_d_req1_tip, ulimit_d_1_d_i_mux_1_d_req1_ge, ulimit_d_1_d_i_mux_1_d_req1_top);

  ulimit_d_2_d_i_d_0_mux_1_d_ack : transition
  generic map(1)
  port map(ulimit_d_2_d_i_d_0_mux_1_d_ack_tip, ulimit_d_2_d_i_d_0_mux_1_d_ack_ge, ulimit_d_2_d_i_d_0_mux_1_d_ack_top);

  ulimit_d_2_d_i_d_0_mux_1_d_req0 : transition
  generic map(1)
  port map(ulimit_d_2_d_i_d_0_mux_1_d_req0_tip, ulimit_d_2_d_i_d_0_mux_1_d_req0_ge, ulimit_d_2_d_i_d_0_mux_1_d_req0_top);

  ulimit_d_2_d_i_d_0_mux_1_d_req1 : transition
  generic map(1)
  port map(ulimit_d_2_d_i_d_0_mux_1_d_req1_tip, ulimit_d_2_d_i_d_0_mux_1_d_req1_ge, ulimit_d_2_d_i_d_0_mux_1_d_req1_top);

  ulimit_d_2_d_i_mux_1_d_ack : transition
  generic map(1)
  port map(ulimit_d_2_d_i_mux_1_d_ack_tip, ulimit_d_2_d_i_mux_1_d_ack_ge, ulimit_d_2_d_i_mux_1_d_ack_top);

  ulimit_d_2_d_i_mux_1_d_req0 : transition
  generic map(1)
  port map(ulimit_d_2_d_i_mux_1_d_req0_tip, ulimit_d_2_d_i_mux_1_d_req0_ge, ulimit_d_2_d_i_mux_1_d_req0_top);

  ulimit_d_2_d_i_mux_1_d_req1 : transition
  generic map(1)
  port map(ulimit_d_2_d_i_mux_1_d_req1_tip, ulimit_d_2_d_i_mux_1_d_req1_ge, ulimit_d_2_d_i_mux_1_d_req1_top);

  place_1_tip(0) <= load_number_d_ack_top;
  place_1_rst(0) <= oper_tmp_d_1_d_i_bool_d_req_top;
  place_10_tip(0) <= no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_top;
  place_10_rst(0) <= ulimit_d_1_d_i_mux_1_d_req0_top;
  place_12_tip(0) <= fin_top;
  place_12_rst(0) <= init_top;
  place_13_tip(0) <= store_location_start_return_d_ack_top;
  place_13_rst(0) <= fin_top;
  place_14_tip(0) <= init_top;
  place_14_rst(0) <= load_number_d_req_top;
  place_15_tip(0) <= load_number_d_req_top;
  place_15_rst(0) <= load_number_d_ack_top;
  place_16_tip(0) <= oper_tmp_d_1_d_i_bool_d_req_top;
  place_16_rst(0) <= oper_tmp_d_1_d_i_bool_d_ack_top;
  place_18_tip(0) <= oper_tmp_d_1_d_i_bool_d_ack_top;
  place_18_rst(0) <= cbr_4_oper_tmp_d_1_d_i_bool_d_req_top;
  place_19_tip(0) <= cbr_4_oper_tmp_d_1_d_i_bool_d_req_top;
  place_19_rst(0) <= entry_to_loopentry_d_i_src_top;
  place_19_rst(1) <= entry_to_no_exit_d_i_src_top;
  place_2_tip(0) <= loopentry_d_i_d_pre_top;
  place_2_rst(0) <= loopentry_d_i_d_entry_top;
  place_20_tip(0) <= entry_to_loopentry_d_i_src_top;
  place_20_rst(0) <= mid_d_0_d_i_mux_1_d_req1_top;
  place_21_tip(0) <= mid_d_0_d_i_mux_1_d_req0_top;
  place_21_tip(1) <= mid_d_0_d_i_mux_1_d_req1_top;
  place_21_rst(0) <= mid_d_0_d_i_mux_1_d_ack_top;
  place_22_tip(0) <= mid_d_0_d_i_mux_1_d_ack_top;
  place_22_rst(0) <= loopentry_d_i_d_pre_top;
  place_23_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_23_rst(0) <= mid_d_0_d_i_mux_1_d_req0_top;
  place_24_tip(0) <= loopentry_d_i_d_entry_top;
  place_24_rst(0) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  place_25_tip(0) <= entry_to_loopentry_d_i_src_top;
  place_25_rst(0) <= llimit_d_2_d_i_mux_1_d_req1_top;
  place_26_tip(0) <= llimit_d_2_d_i_mux_1_d_req0_top;
  place_26_tip(1) <= llimit_d_2_d_i_mux_1_d_req1_top;
  place_26_rst(0) <= llimit_d_2_d_i_mux_1_d_ack_top;
  place_27_tip(0) <= llimit_d_2_d_i_mux_1_d_ack_top;
  place_27_rst(0) <= loopentry_d_i_d_pre_top;
  place_28_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_28_rst(0) <= llimit_d_2_d_i_mux_1_d_req0_top;
  place_29_tip(0) <= loopentry_d_i_d_entry_top;
  place_29_rst(0) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  place_3_tip(0) <= no_exit_d_i_d_pre_top;
  place_3_rst(0) <= no_exit_d_i_d_entry_top;
  place_30_tip(0) <= entry_to_loopentry_d_i_src_top;
  place_30_rst(0) <= ulimit_d_2_d_i_mux_1_d_req1_top;
  place_31_tip(0) <= ulimit_d_2_d_i_mux_1_d_req0_top;
  place_31_tip(1) <= ulimit_d_2_d_i_mux_1_d_req1_top;
  place_31_rst(0) <= ulimit_d_2_d_i_mux_1_d_ack_top;
  place_32_tip(0) <= ulimit_d_2_d_i_mux_1_d_ack_top;
  place_32_rst(0) <= loopentry_d_i_d_pre_top;
  place_33_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_33_rst(0) <= ulimit_d_2_d_i_mux_1_d_req0_top;
  place_34_tip(0) <= loopentry_d_i_d_entry_top;
  place_34_rst(0) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  place_35_tip(0) <= entry_to_loopentry_d_i_src_top;
  place_35_rst(0) <= i_d_0_d_i_mux_1_d_req1_top;
  place_36_tip(0) <= i_d_0_d_i_mux_1_d_req0_top;
  place_36_tip(1) <= i_d_0_d_i_mux_1_d_req1_top;
  place_36_rst(0) <= i_d_0_d_i_mux_1_d_ack_top;
  place_37_tip(0) <= i_d_0_d_i_mux_1_d_ack_top;
  place_37_rst(0) <= loopentry_d_i_d_pre_top;
  place_38_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_38_rst(0) <= i_d_0_d_i_mux_1_d_req0_top;
  place_39_tip(0) <= oper_tmp_d_6_d_i_bool_d_req_top;
  place_39_rst(0) <= oper_tmp_d_6_d_i_bool_d_ack_top;
  place_40_tip(0) <= loopentry_d_i_d_entry_top;
  place_40_rst(0) <= oper_tmp_d_6_d_i_bool_d_req_top;
  place_41_tip(0) <= oper_tmp_d_6_d_i_bool_d_ack_top;
  place_41_rst(0) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  place_42_tip(0) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  place_42_rst(0) <= loopentry_d_i_to_no_exit_d_i_src_top;
  place_42_rst(1) <= loopentry_d_i_to_sqroot_d_exit_src_top;
  place_43_tip(0) <= loopentry_d_i_to_no_exit_d_i_src_top;
  place_43_rst(0) <= llimit_d_2_d_i_d_0_mux_1_d_req1_top;
  place_44_tip(0) <= llimit_d_2_d_i_d_0_mux_1_d_req0_top;
  place_44_tip(1) <= llimit_d_2_d_i_d_0_mux_1_d_req1_top;
  place_44_rst(0) <= llimit_d_2_d_i_d_0_mux_1_d_ack_top;
  place_45_tip(0) <= llimit_d_2_d_i_d_0_mux_1_d_ack_top;
  place_45_rst(0) <= no_exit_d_i_d_pre_top;
  place_46_tip(0) <= entry_to_no_exit_d_i_src_top;
  place_46_rst(0) <= llimit_d_2_d_i_d_0_mux_1_d_req0_top;
  place_47_tip(0) <= loopentry_d_i_to_no_exit_d_i_src_top;
  place_47_rst(0) <= ulimit_d_2_d_i_d_0_mux_1_d_req1_top;
  place_48_tip(0) <= ulimit_d_2_d_i_d_0_mux_1_d_req0_top;
  place_48_tip(1) <= ulimit_d_2_d_i_d_0_mux_1_d_req1_top;
  place_48_rst(0) <= ulimit_d_2_d_i_d_0_mux_1_d_ack_top;
  place_49_tip(0) <= ulimit_d_2_d_i_d_0_mux_1_d_ack_top;
  place_49_rst(0) <= no_exit_d_i_d_pre_top;
  place_5_tip(0) <= loopentry_d_i_to_sqroot_d_exit_src_top;
  place_5_rst(0) <= store_location_start_return_d_req_top;
  place_50_tip(0) <= entry_to_no_exit_d_i_src_top;
  place_50_rst(0) <= ulimit_d_2_d_i_d_0_mux_1_d_req0_top;
  place_51_tip(0) <= loopentry_d_i_to_no_exit_d_i_src_top;
  place_51_rst(0) <= i_d_0_d_i_d_0_mux_1_d_req1_top;
  place_52_tip(0) <= i_d_0_d_i_d_0_mux_1_d_req0_top;
  place_52_tip(1) <= i_d_0_d_i_d_0_mux_1_d_req1_top;
  place_52_rst(0) <= i_d_0_d_i_d_0_mux_1_d_ack_top;
  place_53_tip(0) <= i_d_0_d_i_d_0_mux_1_d_ack_top;
  place_53_rst(0) <= no_exit_d_i_d_pre_top;
  place_54_tip(0) <= entry_to_no_exit_d_i_src_top;
  place_54_rst(0) <= i_d_0_d_i_d_0_mux_1_d_req0_top;
  place_55_tip(0) <= no_exit_d_i_d_entry_top;
  place_55_rst(0) <= cbr_6_oper_tmp_d_17_d_i_bool_d_req_top;
  place_56_tip(0) <= oper_tmp_d_10_d_i_float_d_req_top;
  place_56_rst(0) <= oper_tmp_d_10_d_i_float_d_ack_top;
  place_57_tip(0) <= no_exit_d_i_d_entry_top;
  place_57_rst(0) <= oper_tmp_d_10_d_i_float_d_req_top;
  place_58_tip(0) <= oper_tmp_d_11_d_i_float_d_req_top;
  place_58_rst(0) <= oper_tmp_d_11_d_i_float_d_ack_top;
  place_59_tip(0) <= oper_tmp_d_10_d_i_float_d_ack_top;
  place_59_rst(0) <= oper_tmp_d_11_d_i_float_d_req_top;
  place_60_tip(0) <= oper_tmp_d_14_d_i_float_d_req_top;
  place_60_rst(0) <= oper_tmp_d_14_d_i_float_d_ack_top;
  place_61_tip(0) <= oper_tmp_d_11_d_i_float_d_ack_top;
  place_61_rst(0) <= oper_tmp_d_14_d_i_float_d_req_top;
  place_62_tip(0) <= oper_tmp_d_11_d_i_float_d_ack_top;
  place_62_rst(0) <= oper_tmp_d_14_d_i_float_d_req_top;
  place_63_tip(0) <= oper_tmp_d_17_d_i_bool_d_req_top;
  place_63_rst(0) <= oper_tmp_d_17_d_i_bool_d_ack_top;
  place_64_tip(0) <= oper_tmp_d_14_d_i_float_d_ack_top;
  place_64_rst(0) <= oper_tmp_d_17_d_i_bool_d_req_top;
  place_65_tip(0) <= oper_tmp_d_17_d_i_bool_d_ack_top;
  place_65_rst(0) <= cbr_6_oper_tmp_d_17_d_i_bool_d_req_top;
  place_66_tip(0) <= cbr_6_oper_tmp_d_17_d_i_bool_d_req_top;
  place_66_rst(0) <= no_exit_d_i_to_no_exit_d_i_d_selectcont_src_top;
  place_66_rst(1) <= no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_top;
  place_68_tip(0) <= no_exit_d_i_to_no_exit_d_i_d_selectcont_src_top;
  place_68_rst(0) <= llimit_d_1_d_i_mux_1_d_req1_top;
  place_69_tip(0) <= llimit_d_1_d_i_mux_1_d_req0_top;
  place_69_tip(1) <= llimit_d_1_d_i_mux_1_d_req1_top;
  place_69_rst(0) <= llimit_d_1_d_i_mux_1_d_ack_top;
  place_7_tip(0) <= no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_top;
  place_7_rst(0) <= llimit_d_1_d_i_mux_1_d_req0_top;
  place_70_tip(0) <= llimit_d_1_d_i_mux_1_d_ack_top;
  place_70_rst(0) <= no_exit_d_i_d_selectcont_d_entry_top;
  place_72_tip(0) <= no_exit_d_i_d_selectcont_d_entry_top;
  place_72_rst(0) <= cbr_7_oper_tmp_d_17_d_i_bool_d_req_top;
  place_73_tip(0) <= no_exit_d_i_d_selectcont_d_entry_top;
  place_73_rst(0) <= cbr_7_oper_tmp_d_17_d_i_bool_d_req_top;
  place_74_tip(0) <= cbr_7_oper_tmp_d_17_d_i_bool_d_req_top;
  place_74_rst(0) <= no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_top;
  place_74_rst(1) <= no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_top;
  place_76_tip(0) <= no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_top;
  place_76_rst(0) <= ulimit_d_1_d_i_mux_1_d_req1_top;
  place_77_tip(0) <= ulimit_d_1_d_i_mux_1_d_req0_top;
  place_77_tip(1) <= ulimit_d_1_d_i_mux_1_d_req1_top;
  place_77_rst(0) <= ulimit_d_1_d_i_mux_1_d_ack_top;
  place_78_tip(0) <= ulimit_d_1_d_i_mux_1_d_ack_top;
  place_78_rst(0) <= no_exit_d_i_d_selectcont_d_selectcont_d_entry_top;
  place_80_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_d_entry_top;
  place_80_rst(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_81_tip(0) <= oper_inc_d_i_int_d_req_top;
  place_81_rst(0) <= oper_inc_d_i_int_d_ack_top;
  place_82_tip(0) <= no_exit_d_i_d_selectcont_d_selectcont_d_entry_top;
  place_82_rst(0) <= oper_inc_d_i_int_d_req_top;
  place_83_tip(0) <= oper_inc_d_i_int_d_ack_top;
  place_83_rst(0) <= no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_top;
  place_84_tip(0) <= store_location_start_return_d_req_top;
  place_84_rst(0) <= store_location_start_return_d_ack_top;

  cbr_4_oper_tmp_d_1_d_i_bool_d_req_tip(0) <= place_18_top;
  cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip(0) <= place_24_top;
  cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip(1) <= place_29_top;
  cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip(2) <= place_34_top;
  cbr_5_oper_tmp_d_6_d_i_bool_d_req_tip(3) <= place_41_top;
  cbr_6_oper_tmp_d_17_d_i_bool_d_req_tip(0) <= place_55_top;
  cbr_6_oper_tmp_d_17_d_i_bool_d_req_tip(1) <= place_65_top;
  cbr_7_oper_tmp_d_17_d_i_bool_d_req_tip(0) <= place_72_top;
  cbr_7_oper_tmp_d_17_d_i_bool_d_req_tip(1) <= place_73_top;
  entry_to_loopentry_d_i_src_tip(0) <= place_19_top;
  entry_to_no_exit_d_i_src_tip(0) <= place_19_top;
  fin_tip(0) <= place_13_top;
  i_d_0_d_i_d_0_mux_1_d_ack_tip(0) <= place_52_top;
  i_d_0_d_i_d_0_mux_1_d_req0_tip(0) <= place_54_top;
  i_d_0_d_i_d_0_mux_1_d_req1_tip(0) <= place_51_top;
  i_d_0_d_i_mux_1_d_ack_tip(0) <= place_36_top;
  i_d_0_d_i_mux_1_d_req0_tip(0) <= place_38_top;
  i_d_0_d_i_mux_1_d_req1_tip(0) <= place_35_top;
  init_tip(0) <= place_12_top;
  llimit_d_1_d_i_mux_1_d_ack_tip(0) <= place_69_top;
  llimit_d_1_d_i_mux_1_d_req0_tip(0) <= place_7_top;
  llimit_d_1_d_i_mux_1_d_req1_tip(0) <= place_68_top;
  llimit_d_2_d_i_d_0_mux_1_d_ack_tip(0) <= place_44_top;
  llimit_d_2_d_i_d_0_mux_1_d_req0_tip(0) <= place_46_top;
  llimit_d_2_d_i_d_0_mux_1_d_req1_tip(0) <= place_43_top;
  llimit_d_2_d_i_mux_1_d_ack_tip(0) <= place_26_top;
  llimit_d_2_d_i_mux_1_d_req0_tip(0) <= place_28_top;
  llimit_d_2_d_i_mux_1_d_req1_tip(0) <= place_25_top;
  load_number_d_ack_tip(0) <= place_15_top;
  load_number_d_req_tip(0) <= place_14_top;
  loopentry_d_i_d_entry_tip(0) <= place_2_top;
  loopentry_d_i_d_pre_tip(0) <= place_22_top;
  loopentry_d_i_d_pre_tip(1) <= place_27_top;
  loopentry_d_i_d_pre_tip(2) <= place_32_top;
  loopentry_d_i_d_pre_tip(3) <= place_37_top;
  loopentry_d_i_to_no_exit_d_i_src_tip(0) <= place_42_top;
  loopentry_d_i_to_sqroot_d_exit_src_tip(0) <= place_42_top;
  mid_d_0_d_i_mux_1_d_ack_tip(0) <= place_21_top;
  mid_d_0_d_i_mux_1_d_req0_tip(0) <= place_23_top;
  mid_d_0_d_i_mux_1_d_req1_tip(0) <= place_20_top;
  no_exit_d_i_d_entry_tip(0) <= place_3_top;
  no_exit_d_i_d_pre_tip(0) <= place_45_top;
  no_exit_d_i_d_pre_tip(1) <= place_49_top;
  no_exit_d_i_d_pre_tip(2) <= place_53_top;
  no_exit_d_i_d_selectcont_d_entry_tip(0) <= place_70_top;
  no_exit_d_i_d_selectcont_d_selectcont_d_entry_tip(0) <= place_78_top;
  no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_tip(0) <= place_80_top;
  no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_tip(1) <= place_83_top;
  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_tip(0) <= place_74_top;
  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_tip(0) <= place_74_top;
  no_exit_d_i_to_no_exit_d_i_d_selectcont_src_tip(0) <= place_66_top;
  no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_tip(0) <= place_66_top;
  oper_inc_d_i_int_d_ack_tip(0) <= place_81_top;
  oper_inc_d_i_int_d_req_tip(0) <= place_82_top;
  oper_tmp_d_10_d_i_float_d_ack_tip(0) <= place_56_top;
  oper_tmp_d_10_d_i_float_d_req_tip(0) <= place_57_top;
  oper_tmp_d_11_d_i_float_d_ack_tip(0) <= place_58_top;
  oper_tmp_d_11_d_i_float_d_req_tip(0) <= place_59_top;
  oper_tmp_d_14_d_i_float_d_ack_tip(0) <= place_60_top;
  oper_tmp_d_14_d_i_float_d_req_tip(0) <= place_61_top;
  oper_tmp_d_14_d_i_float_d_req_tip(1) <= place_62_top;
  oper_tmp_d_17_d_i_bool_d_ack_tip(0) <= place_63_top;
  oper_tmp_d_17_d_i_bool_d_req_tip(0) <= place_64_top;
  oper_tmp_d_1_d_i_bool_d_ack_tip(0) <= place_16_top;
  oper_tmp_d_1_d_i_bool_d_req_tip(0) <= place_1_top;
  oper_tmp_d_6_d_i_bool_d_ack_tip(0) <= place_39_top;
  oper_tmp_d_6_d_i_bool_d_req_tip(0) <= place_40_top;
  store_location_start_return_d_ack_tip(0) <= place_84_top;
  store_location_start_return_d_req_tip(0) <= place_5_top;
  ulimit_d_1_d_i_mux_1_d_ack_tip(0) <= place_77_top;
  ulimit_d_1_d_i_mux_1_d_req0_tip(0) <= place_10_top;
  ulimit_d_1_d_i_mux_1_d_req1_tip(0) <= place_76_top;
  ulimit_d_2_d_i_d_0_mux_1_d_ack_tip(0) <= place_48_top;
  ulimit_d_2_d_i_d_0_mux_1_d_req0_tip(0) <= place_50_top;
  ulimit_d_2_d_i_d_0_mux_1_d_req1_tip(0) <= place_47_top;
  ulimit_d_2_d_i_mux_1_d_ack_tip(0) <= place_31_top;
  ulimit_d_2_d_i_mux_1_d_req0_tip(0) <= place_33_top;
  ulimit_d_2_d_i_mux_1_d_req1_tip(0) <= place_30_top;

  cbr_4_oper_tmp_d_1_d_i_bool_d_req_ge <= '1';
  op(4) <= cbr_4_oper_tmp_d_1_d_i_bool_d_req_top;
  cbr_5_oper_tmp_d_6_d_i_bool_d_req_ge <= '1';
  op(14) <= cbr_5_oper_tmp_d_6_d_i_bool_d_req_top;
  cbr_6_oper_tmp_d_17_d_i_bool_d_req_ge <= '1';
  op(25) <= cbr_6_oper_tmp_d_17_d_i_bool_d_req_top;
  cbr_7_oper_tmp_d_17_d_i_bool_d_req_ge <= '1';
  op(28) <= cbr_7_oper_tmp_d_17_d_i_bool_d_req_top;
  entry_to_loopentry_d_i_src_ge <= ip(4);
  entry_to_no_exit_d_i_src_ge <= ip(5);
  fin_ge <= '1';
  op(1) <= fin_top;
  i_d_0_d_i_d_0_mux_1_d_ack_ge <= ip(15);
  i_d_0_d_i_d_0_mux_1_d_req0_ge <= '1';
  op(20) <= i_d_0_d_i_d_0_mux_1_d_req0_top;
  i_d_0_d_i_d_0_mux_1_d_req1_ge <= '1';
  op(19) <= i_d_0_d_i_d_0_mux_1_d_req1_top;
  i_d_0_d_i_mux_1_d_ack_ge <= ip(9);
  i_d_0_d_i_mux_1_d_req0_ge <= '1';
  op(12) <= i_d_0_d_i_mux_1_d_req0_top;
  i_d_0_d_i_mux_1_d_req1_ge <= '1';
  op(11) <= i_d_0_d_i_mux_1_d_req1_top;
  init_ge <= ip(1);
  llimit_d_1_d_i_mux_1_d_ack_ge <= ip(22);
  llimit_d_1_d_i_mux_1_d_req0_ge <= '1';
  op(27) <= llimit_d_1_d_i_mux_1_d_req0_top;
  llimit_d_1_d_i_mux_1_d_req1_ge <= '1';
  op(26) <= llimit_d_1_d_i_mux_1_d_req1_top;
  llimit_d_2_d_i_d_0_mux_1_d_ack_ge <= ip(13);
  llimit_d_2_d_i_d_0_mux_1_d_req0_ge <= '1';
  op(16) <= llimit_d_2_d_i_d_0_mux_1_d_req0_top;
  llimit_d_2_d_i_d_0_mux_1_d_req1_ge <= '1';
  op(15) <= llimit_d_2_d_i_d_0_mux_1_d_req1_top;
  llimit_d_2_d_i_mux_1_d_ack_ge <= ip(7);
  llimit_d_2_d_i_mux_1_d_req0_ge <= '1';
  op(8) <= llimit_d_2_d_i_mux_1_d_req0_top;
  llimit_d_2_d_i_mux_1_d_req1_ge <= '1';
  op(7) <= llimit_d_2_d_i_mux_1_d_req1_top;
  load_number_d_ack_ge <= ip(2);
  load_number_d_req_ge <= '1';
  op(2) <= load_number_d_req_top;
  loopentry_d_i_d_entry_ge <= '1';
  loopentry_d_i_d_pre_ge <= '1';
  loopentry_d_i_to_no_exit_d_i_src_ge <= ip(11);
  loopentry_d_i_to_sqroot_d_exit_src_ge <= ip(12);
  mid_d_0_d_i_mux_1_d_ack_ge <= ip(6);
  mid_d_0_d_i_mux_1_d_req0_ge <= '1';
  op(6) <= mid_d_0_d_i_mux_1_d_req0_top;
  mid_d_0_d_i_mux_1_d_req1_ge <= '1';
  op(5) <= mid_d_0_d_i_mux_1_d_req1_top;
  no_exit_d_i_d_entry_ge <= '1';
  no_exit_d_i_d_pre_ge <= '1';
  no_exit_d_i_d_selectcont_d_entry_ge <= '1';
  no_exit_d_i_d_selectcont_d_selectcont_d_entry_ge <= '1';
  no_exit_d_i_d_selectcont_d_selectcont_to_loopentry_d_i_src_ge <= '1';
  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selectcont_src_ge <= ip(24);
  no_exit_d_i_d_selectcont_to_no_exit_d_i_d_selectcont_d_selecttrue_src_ge <= ip(23);
  no_exit_d_i_to_no_exit_d_i_d_selectcont_src_ge <= ip(21);
  no_exit_d_i_to_no_exit_d_i_d_selecttrue_src_ge <= ip(20);
  oper_inc_d_i_int_d_ack_ge <= ip(26);
  oper_inc_d_i_int_d_req_ge <= '1';
  op(31) <= oper_inc_d_i_int_d_req_top;
  oper_tmp_d_10_d_i_float_d_ack_ge <= ip(16);
  oper_tmp_d_10_d_i_float_d_req_ge <= '1';
  op(21) <= oper_tmp_d_10_d_i_float_d_req_top;
  oper_tmp_d_11_d_i_float_d_ack_ge <= ip(17);
  oper_tmp_d_11_d_i_float_d_req_ge <= '1';
  op(22) <= oper_tmp_d_11_d_i_float_d_req_top;
  oper_tmp_d_14_d_i_float_d_ack_ge <= ip(18);
  oper_tmp_d_14_d_i_float_d_req_ge <= '1';
  op(23) <= oper_tmp_d_14_d_i_float_d_req_top;
  oper_tmp_d_17_d_i_bool_d_ack_ge <= ip(19);
  oper_tmp_d_17_d_i_bool_d_req_ge <= '1';
  op(24) <= oper_tmp_d_17_d_i_bool_d_req_top;
  oper_tmp_d_1_d_i_bool_d_ack_ge <= ip(3);
  oper_tmp_d_1_d_i_bool_d_req_ge <= '1';
  op(3) <= oper_tmp_d_1_d_i_bool_d_req_top;
  oper_tmp_d_6_d_i_bool_d_ack_ge <= ip(10);
  oper_tmp_d_6_d_i_bool_d_req_ge <= '1';
  op(13) <= oper_tmp_d_6_d_i_bool_d_req_top;
  store_location_start_return_d_ack_ge <= ip(27);
  store_location_start_return_d_req_ge <= '1';
  op(32) <= store_location_start_return_d_req_top;
  ulimit_d_1_d_i_mux_1_d_ack_ge <= ip(25);
  ulimit_d_1_d_i_mux_1_d_req0_ge <= '1';
  op(30) <= ulimit_d_1_d_i_mux_1_d_req0_top;
  ulimit_d_1_d_i_mux_1_d_req1_ge <= '1';
  op(29) <= ulimit_d_1_d_i_mux_1_d_req1_top;
  ulimit_d_2_d_i_d_0_mux_1_d_ack_ge <= ip(14);
  ulimit_d_2_d_i_d_0_mux_1_d_req0_ge <= '1';
  op(18) <= ulimit_d_2_d_i_d_0_mux_1_d_req0_top;
  ulimit_d_2_d_i_d_0_mux_1_d_req1_ge <= '1';
  op(17) <= ulimit_d_2_d_i_d_0_mux_1_d_req1_top;
  ulimit_d_2_d_i_mux_1_d_ack_ge <= ip(8);
  ulimit_d_2_d_i_mux_1_d_req0_ge <= '1';
  op(10) <= ulimit_d_2_d_i_mux_1_d_req0_top;
  ulimit_d_2_d_i_mux_1_d_req1_ge <= '1';
  op(9) <= ulimit_d_2_d_i_mux_1_d_req1_top;

end behavioral;
