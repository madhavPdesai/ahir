
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;

entity start_ln is
  port(
    clk : in std_logic;
    reset : in std_logic;
    start_cp_LambdaIn : out BooleanArray(292 downto 1);
    start_cp_LambdaOut : in BooleanArray(294 downto 1);
    start_dp_SigmaIn : out BooleanArray(294 downto 1);
    start_dp_SigmaOut : in BooleanArray(292 downto 1));
end start_ln;

architecture default_arch of start_ln is
begin
  start_cp_LambdaIn(1) <= start_dp_SigmaOut(1);
  start_cp_LambdaIn(2) <= start_dp_SigmaOut(2);
  start_cp_LambdaIn(3) <= start_dp_SigmaOut(3);
  start_cp_LambdaIn(4) <= start_dp_SigmaOut(4);
  start_cp_LambdaIn(5) <= start_dp_SigmaOut(5);
  start_cp_LambdaIn(6) <= start_dp_SigmaOut(6);
  start_cp_LambdaIn(7) <= start_dp_SigmaOut(7);
  start_cp_LambdaIn(8) <= start_dp_SigmaOut(8);
  start_cp_LambdaIn(9) <= start_dp_SigmaOut(9);
  start_cp_LambdaIn(10) <= start_dp_SigmaOut(10);
  start_cp_LambdaIn(11) <= start_dp_SigmaOut(11);
  start_cp_LambdaIn(12) <= start_dp_SigmaOut(12);
  start_cp_LambdaIn(13) <= start_dp_SigmaOut(13);
  start_cp_LambdaIn(14) <= start_dp_SigmaOut(14);
  start_cp_LambdaIn(15) <= start_dp_SigmaOut(15);
  start_cp_LambdaIn(16) <= start_dp_SigmaOut(16);
  start_cp_LambdaIn(17) <= start_dp_SigmaOut(17);
  start_cp_LambdaIn(18) <= start_dp_SigmaOut(18);
  start_cp_LambdaIn(19) <= start_dp_SigmaOut(19);
  start_cp_LambdaIn(20) <= start_dp_SigmaOut(20);
  start_cp_LambdaIn(21) <= start_dp_SigmaOut(21);
  start_cp_LambdaIn(22) <= start_dp_SigmaOut(22);
  start_cp_LambdaIn(23) <= start_dp_SigmaOut(23);
  start_cp_LambdaIn(24) <= start_dp_SigmaOut(24);
  start_cp_LambdaIn(25) <= start_dp_SigmaOut(25);
  start_cp_LambdaIn(26) <= start_dp_SigmaOut(26);
  start_cp_LambdaIn(27) <= start_dp_SigmaOut(27);
  start_cp_LambdaIn(28) <= start_dp_SigmaOut(28);
  start_cp_LambdaIn(29) <= start_dp_SigmaOut(29);
  start_cp_LambdaIn(30) <= start_dp_SigmaOut(30);
  start_cp_LambdaIn(31) <= start_dp_SigmaOut(31);
  start_cp_LambdaIn(32) <= start_dp_SigmaOut(32);
  start_cp_LambdaIn(33) <= start_dp_SigmaOut(33);
  start_cp_LambdaIn(34) <= start_dp_SigmaOut(34);
  start_cp_LambdaIn(35) <= start_dp_SigmaOut(35);
  start_cp_LambdaIn(36) <= start_dp_SigmaOut(36);
  start_cp_LambdaIn(37) <= start_dp_SigmaOut(37);
  start_cp_LambdaIn(38) <= start_dp_SigmaOut(38);
  start_cp_LambdaIn(39) <= start_dp_SigmaOut(39);
  start_cp_LambdaIn(40) <= start_dp_SigmaOut(40);
  start_cp_LambdaIn(41) <= start_dp_SigmaOut(41);
  start_cp_LambdaIn(42) <= start_dp_SigmaOut(42);
  start_cp_LambdaIn(43) <= start_dp_SigmaOut(43);
  start_cp_LambdaIn(44) <= start_dp_SigmaOut(44);
  start_cp_LambdaIn(45) <= start_dp_SigmaOut(45);
  start_cp_LambdaIn(46) <= start_dp_SigmaOut(46);
  start_cp_LambdaIn(47) <= start_dp_SigmaOut(47);
  start_cp_LambdaIn(48) <= start_dp_SigmaOut(48);
  start_cp_LambdaIn(49) <= start_dp_SigmaOut(49);
  start_cp_LambdaIn(50) <= start_dp_SigmaOut(50);
  start_cp_LambdaIn(51) <= start_dp_SigmaOut(51);
  start_cp_LambdaIn(52) <= start_dp_SigmaOut(52);
  start_cp_LambdaIn(53) <= start_dp_SigmaOut(53);
  start_cp_LambdaIn(54) <= start_dp_SigmaOut(54);
  start_cp_LambdaIn(55) <= start_dp_SigmaOut(55);
  start_cp_LambdaIn(56) <= start_dp_SigmaOut(56);
  start_cp_LambdaIn(57) <= start_dp_SigmaOut(57);
  start_cp_LambdaIn(58) <= start_dp_SigmaOut(58);
  start_cp_LambdaIn(59) <= start_dp_SigmaOut(59);
  start_cp_LambdaIn(60) <= start_dp_SigmaOut(60);
  start_cp_LambdaIn(61) <= start_dp_SigmaOut(61);
  start_cp_LambdaIn(62) <= start_dp_SigmaOut(62);
  start_cp_LambdaIn(63) <= start_dp_SigmaOut(63);
  start_cp_LambdaIn(64) <= start_dp_SigmaOut(64);
  start_cp_LambdaIn(65) <= start_dp_SigmaOut(65);
  start_cp_LambdaIn(66) <= start_dp_SigmaOut(66);
  start_cp_LambdaIn(67) <= start_dp_SigmaOut(67);
  start_cp_LambdaIn(68) <= start_dp_SigmaOut(68);
  start_cp_LambdaIn(69) <= start_dp_SigmaOut(69);
  start_cp_LambdaIn(70) <= start_dp_SigmaOut(70);
  start_cp_LambdaIn(71) <= start_dp_SigmaOut(71);
  start_cp_LambdaIn(72) <= start_dp_SigmaOut(72);
  start_cp_LambdaIn(73) <= start_dp_SigmaOut(73);
  start_cp_LambdaIn(74) <= start_dp_SigmaOut(74);
  start_cp_LambdaIn(75) <= start_dp_SigmaOut(75);
  start_cp_LambdaIn(76) <= start_dp_SigmaOut(76);
  start_cp_LambdaIn(77) <= start_dp_SigmaOut(77);
  start_cp_LambdaIn(78) <= start_dp_SigmaOut(78);
  start_cp_LambdaIn(79) <= start_dp_SigmaOut(79);
  start_cp_LambdaIn(80) <= start_dp_SigmaOut(80);
  start_cp_LambdaIn(81) <= start_dp_SigmaOut(81);
  start_cp_LambdaIn(82) <= start_dp_SigmaOut(82);
  start_cp_LambdaIn(83) <= start_dp_SigmaOut(83);
  start_cp_LambdaIn(84) <= start_dp_SigmaOut(84);
  start_cp_LambdaIn(85) <= start_dp_SigmaOut(85);
  start_cp_LambdaIn(86) <= start_dp_SigmaOut(86);
  start_cp_LambdaIn(87) <= start_dp_SigmaOut(87);
  start_cp_LambdaIn(88) <= start_dp_SigmaOut(88);
  start_cp_LambdaIn(89) <= start_dp_SigmaOut(89);
  start_cp_LambdaIn(90) <= start_dp_SigmaOut(90);
  start_cp_LambdaIn(91) <= start_dp_SigmaOut(91);
  start_cp_LambdaIn(92) <= start_dp_SigmaOut(92);
  start_cp_LambdaIn(93) <= start_dp_SigmaOut(93);
  start_cp_LambdaIn(94) <= start_dp_SigmaOut(94);
  start_cp_LambdaIn(95) <= start_dp_SigmaOut(95);
  start_cp_LambdaIn(96) <= start_dp_SigmaOut(96);
  start_cp_LambdaIn(97) <= start_dp_SigmaOut(97);
  start_cp_LambdaIn(98) <= start_dp_SigmaOut(98);
  start_cp_LambdaIn(99) <= start_dp_SigmaOut(99);
  start_cp_LambdaIn(100) <= start_dp_SigmaOut(100);
  start_cp_LambdaIn(101) <= start_dp_SigmaOut(101);
  start_cp_LambdaIn(102) <= start_dp_SigmaOut(102);
  start_cp_LambdaIn(103) <= start_dp_SigmaOut(103);
  start_cp_LambdaIn(104) <= start_dp_SigmaOut(104);
  start_cp_LambdaIn(105) <= start_dp_SigmaOut(105);
  start_cp_LambdaIn(106) <= start_dp_SigmaOut(106);
  start_cp_LambdaIn(107) <= start_dp_SigmaOut(107);
  start_cp_LambdaIn(108) <= start_dp_SigmaOut(108);
  start_cp_LambdaIn(109) <= start_dp_SigmaOut(109);
  start_cp_LambdaIn(110) <= start_dp_SigmaOut(110);
  start_cp_LambdaIn(111) <= start_dp_SigmaOut(111);
  start_cp_LambdaIn(112) <= start_dp_SigmaOut(112);
  start_cp_LambdaIn(113) <= start_dp_SigmaOut(113);
  start_cp_LambdaIn(114) <= start_dp_SigmaOut(114);
  start_cp_LambdaIn(115) <= start_dp_SigmaOut(115);
  start_cp_LambdaIn(116) <= start_dp_SigmaOut(116);
  start_cp_LambdaIn(117) <= start_dp_SigmaOut(117);
  start_cp_LambdaIn(118) <= start_dp_SigmaOut(118);
  start_cp_LambdaIn(119) <= start_dp_SigmaOut(119);
  start_cp_LambdaIn(120) <= start_dp_SigmaOut(120);
  start_cp_LambdaIn(121) <= start_dp_SigmaOut(121);
  start_cp_LambdaIn(122) <= start_dp_SigmaOut(122);
  start_cp_LambdaIn(123) <= start_dp_SigmaOut(123);
  start_cp_LambdaIn(124) <= start_dp_SigmaOut(124);
  start_cp_LambdaIn(125) <= start_dp_SigmaOut(125);
  start_cp_LambdaIn(126) <= start_dp_SigmaOut(126);
  start_cp_LambdaIn(127) <= start_dp_SigmaOut(127);
  start_cp_LambdaIn(128) <= start_dp_SigmaOut(128);
  start_cp_LambdaIn(129) <= start_dp_SigmaOut(129);
  start_cp_LambdaIn(130) <= start_dp_SigmaOut(130);
  start_cp_LambdaIn(131) <= start_dp_SigmaOut(131);
  start_cp_LambdaIn(132) <= start_dp_SigmaOut(132);
  start_cp_LambdaIn(133) <= start_dp_SigmaOut(133);
  start_cp_LambdaIn(134) <= start_dp_SigmaOut(134);
  start_cp_LambdaIn(135) <= start_dp_SigmaOut(135);
  start_cp_LambdaIn(136) <= start_dp_SigmaOut(136);
  start_cp_LambdaIn(137) <= start_dp_SigmaOut(137);
  start_cp_LambdaIn(138) <= start_dp_SigmaOut(138);
  start_cp_LambdaIn(139) <= start_dp_SigmaOut(139);
  start_cp_LambdaIn(140) <= start_dp_SigmaOut(140);
  start_cp_LambdaIn(141) <= start_dp_SigmaOut(141);
  start_cp_LambdaIn(142) <= start_dp_SigmaOut(142);
  start_cp_LambdaIn(143) <= start_dp_SigmaOut(143);
  start_cp_LambdaIn(144) <= start_dp_SigmaOut(144);
  start_cp_LambdaIn(145) <= start_dp_SigmaOut(145);
  start_cp_LambdaIn(146) <= start_dp_SigmaOut(146);
  start_cp_LambdaIn(147) <= start_dp_SigmaOut(147);
  start_cp_LambdaIn(148) <= start_dp_SigmaOut(148);
  start_cp_LambdaIn(149) <= start_dp_SigmaOut(149);
  start_cp_LambdaIn(150) <= start_dp_SigmaOut(150);
  start_cp_LambdaIn(151) <= start_dp_SigmaOut(151);
  start_cp_LambdaIn(152) <= start_dp_SigmaOut(152);
  start_cp_LambdaIn(153) <= start_dp_SigmaOut(153);
  start_cp_LambdaIn(154) <= start_dp_SigmaOut(154);
  start_cp_LambdaIn(155) <= start_dp_SigmaOut(155);
  start_cp_LambdaIn(156) <= start_dp_SigmaOut(156);
  start_cp_LambdaIn(157) <= start_dp_SigmaOut(157);
  start_cp_LambdaIn(158) <= start_dp_SigmaOut(158);
  start_cp_LambdaIn(159) <= start_dp_SigmaOut(159);
  start_cp_LambdaIn(160) <= start_dp_SigmaOut(160);
  start_cp_LambdaIn(161) <= start_dp_SigmaOut(161);
  start_cp_LambdaIn(162) <= start_dp_SigmaOut(162);
  start_cp_LambdaIn(163) <= start_dp_SigmaOut(163);
  start_cp_LambdaIn(164) <= start_dp_SigmaOut(164);
  start_cp_LambdaIn(165) <= start_dp_SigmaOut(165);
  start_cp_LambdaIn(166) <= start_dp_SigmaOut(166);
  start_cp_LambdaIn(167) <= start_dp_SigmaOut(167);
  start_cp_LambdaIn(168) <= start_dp_SigmaOut(168);
  start_cp_LambdaIn(169) <= start_dp_SigmaOut(169);
  start_cp_LambdaIn(170) <= start_dp_SigmaOut(170);
  start_cp_LambdaIn(171) <= start_dp_SigmaOut(171);
  start_cp_LambdaIn(172) <= start_dp_SigmaOut(172);
  start_cp_LambdaIn(173) <= start_dp_SigmaOut(173);
  start_cp_LambdaIn(174) <= start_dp_SigmaOut(174);
  start_cp_LambdaIn(175) <= start_dp_SigmaOut(175);
  start_cp_LambdaIn(176) <= start_dp_SigmaOut(176);
  start_cp_LambdaIn(177) <= start_dp_SigmaOut(177);
  start_cp_LambdaIn(178) <= start_dp_SigmaOut(178);
  start_cp_LambdaIn(179) <= start_dp_SigmaOut(179);
  start_cp_LambdaIn(180) <= start_dp_SigmaOut(180);
  start_cp_LambdaIn(181) <= start_dp_SigmaOut(181);
  start_cp_LambdaIn(182) <= start_dp_SigmaOut(182);
  start_cp_LambdaIn(183) <= start_dp_SigmaOut(183);
  start_cp_LambdaIn(184) <= start_dp_SigmaOut(184);
  start_cp_LambdaIn(185) <= start_dp_SigmaOut(185);
  start_cp_LambdaIn(186) <= start_dp_SigmaOut(186);
  start_cp_LambdaIn(187) <= start_dp_SigmaOut(187);
  start_cp_LambdaIn(188) <= start_dp_SigmaOut(188);
  start_cp_LambdaIn(189) <= start_dp_SigmaOut(189);
  start_cp_LambdaIn(190) <= start_dp_SigmaOut(190);
  start_cp_LambdaIn(191) <= start_dp_SigmaOut(191);
  start_cp_LambdaIn(192) <= start_dp_SigmaOut(192);
  start_cp_LambdaIn(193) <= start_dp_SigmaOut(193);
  start_cp_LambdaIn(194) <= start_dp_SigmaOut(194);
  start_cp_LambdaIn(195) <= start_dp_SigmaOut(195);
  start_cp_LambdaIn(196) <= start_dp_SigmaOut(196);
  start_cp_LambdaIn(197) <= start_dp_SigmaOut(197);
  start_cp_LambdaIn(198) <= start_dp_SigmaOut(198);
  start_cp_LambdaIn(199) <= start_dp_SigmaOut(199);
  start_cp_LambdaIn(200) <= start_dp_SigmaOut(200);
  start_cp_LambdaIn(201) <= start_dp_SigmaOut(201);
  start_cp_LambdaIn(202) <= start_dp_SigmaOut(202);
  start_cp_LambdaIn(203) <= start_dp_SigmaOut(203);
  start_cp_LambdaIn(204) <= start_dp_SigmaOut(204);
  start_cp_LambdaIn(205) <= start_dp_SigmaOut(205);
  start_cp_LambdaIn(206) <= start_dp_SigmaOut(206);
  start_cp_LambdaIn(207) <= start_dp_SigmaOut(207);
  start_cp_LambdaIn(208) <= start_dp_SigmaOut(208);
  start_cp_LambdaIn(209) <= start_dp_SigmaOut(209);
  start_cp_LambdaIn(210) <= start_dp_SigmaOut(210);
  start_cp_LambdaIn(211) <= start_dp_SigmaOut(211);
  start_cp_LambdaIn(212) <= start_dp_SigmaOut(212);
  start_cp_LambdaIn(213) <= start_dp_SigmaOut(213);
  start_cp_LambdaIn(214) <= start_dp_SigmaOut(214);
  start_cp_LambdaIn(215) <= start_dp_SigmaOut(215);
  start_cp_LambdaIn(216) <= start_dp_SigmaOut(216);
  start_cp_LambdaIn(217) <= start_dp_SigmaOut(217);
  start_cp_LambdaIn(218) <= start_dp_SigmaOut(218);
  start_cp_LambdaIn(219) <= start_dp_SigmaOut(219);
  start_cp_LambdaIn(220) <= start_dp_SigmaOut(220);
  start_cp_LambdaIn(221) <= start_dp_SigmaOut(221);
  start_cp_LambdaIn(222) <= start_dp_SigmaOut(222);
  start_cp_LambdaIn(223) <= start_dp_SigmaOut(223);
  start_cp_LambdaIn(224) <= start_dp_SigmaOut(224);
  start_cp_LambdaIn(225) <= start_dp_SigmaOut(225);
  start_cp_LambdaIn(226) <= start_dp_SigmaOut(226);
  start_cp_LambdaIn(227) <= start_dp_SigmaOut(227);
  start_cp_LambdaIn(228) <= start_dp_SigmaOut(228);
  start_cp_LambdaIn(229) <= start_dp_SigmaOut(229);
  start_cp_LambdaIn(230) <= start_dp_SigmaOut(230);
  start_cp_LambdaIn(231) <= start_dp_SigmaOut(231);
  start_cp_LambdaIn(232) <= start_dp_SigmaOut(232);
  start_cp_LambdaIn(233) <= start_dp_SigmaOut(233);
  start_cp_LambdaIn(234) <= start_dp_SigmaOut(234);
  start_cp_LambdaIn(235) <= start_dp_SigmaOut(235);
  start_cp_LambdaIn(236) <= start_dp_SigmaOut(236);
  start_cp_LambdaIn(237) <= start_dp_SigmaOut(237);
  start_cp_LambdaIn(238) <= start_dp_SigmaOut(238);
  start_cp_LambdaIn(239) <= start_dp_SigmaOut(239);
  start_cp_LambdaIn(240) <= start_dp_SigmaOut(240);
  start_cp_LambdaIn(241) <= start_dp_SigmaOut(241);
  start_cp_LambdaIn(242) <= start_dp_SigmaOut(242);
  start_cp_LambdaIn(243) <= start_dp_SigmaOut(243);
  start_cp_LambdaIn(244) <= start_dp_SigmaOut(244);
  start_cp_LambdaIn(245) <= start_dp_SigmaOut(245);
  start_cp_LambdaIn(246) <= start_dp_SigmaOut(246);
  start_cp_LambdaIn(247) <= start_dp_SigmaOut(247);
  start_cp_LambdaIn(248) <= start_dp_SigmaOut(248);
  start_cp_LambdaIn(249) <= start_dp_SigmaOut(249);
  start_cp_LambdaIn(250) <= start_dp_SigmaOut(250);
  start_cp_LambdaIn(251) <= start_dp_SigmaOut(251);
  start_cp_LambdaIn(252) <= start_dp_SigmaOut(252);
  start_cp_LambdaIn(253) <= start_dp_SigmaOut(253);
  start_cp_LambdaIn(254) <= start_dp_SigmaOut(254);
  start_cp_LambdaIn(255) <= start_dp_SigmaOut(255);
  start_cp_LambdaIn(256) <= start_dp_SigmaOut(256);
  start_cp_LambdaIn(257) <= start_dp_SigmaOut(257);
  start_cp_LambdaIn(258) <= start_dp_SigmaOut(258);
  start_cp_LambdaIn(259) <= start_dp_SigmaOut(259);
  start_cp_LambdaIn(260) <= start_dp_SigmaOut(260);
  start_cp_LambdaIn(261) <= start_dp_SigmaOut(261);
  start_cp_LambdaIn(262) <= start_dp_SigmaOut(262);
  start_cp_LambdaIn(263) <= start_dp_SigmaOut(263);
  start_cp_LambdaIn(264) <= start_dp_SigmaOut(264);
  start_cp_LambdaIn(265) <= start_dp_SigmaOut(265);
  start_cp_LambdaIn(266) <= start_dp_SigmaOut(266);
  start_cp_LambdaIn(267) <= start_dp_SigmaOut(267);
  start_cp_LambdaIn(268) <= start_dp_SigmaOut(268);
  start_cp_LambdaIn(269) <= start_dp_SigmaOut(269);
  start_cp_LambdaIn(270) <= start_dp_SigmaOut(270);
  start_cp_LambdaIn(271) <= start_dp_SigmaOut(271);
  start_cp_LambdaIn(272) <= start_dp_SigmaOut(272);
  start_cp_LambdaIn(273) <= start_dp_SigmaOut(273);
  start_cp_LambdaIn(274) <= start_dp_SigmaOut(274);
  start_cp_LambdaIn(275) <= start_dp_SigmaOut(275);
  start_cp_LambdaIn(276) <= start_dp_SigmaOut(276);
  start_cp_LambdaIn(277) <= start_dp_SigmaOut(277);
  start_cp_LambdaIn(278) <= start_dp_SigmaOut(278);
  start_cp_LambdaIn(279) <= start_dp_SigmaOut(279);
  start_cp_LambdaIn(280) <= start_dp_SigmaOut(280);
  start_cp_LambdaIn(281) <= start_dp_SigmaOut(281);
  start_cp_LambdaIn(282) <= start_dp_SigmaOut(282);
  start_cp_LambdaIn(283) <= start_dp_SigmaOut(283);
  start_cp_LambdaIn(284) <= start_dp_SigmaOut(284);
  start_cp_LambdaIn(285) <= start_dp_SigmaOut(285);
  start_cp_LambdaIn(286) <= start_dp_SigmaOut(286);
  start_cp_LambdaIn(287) <= start_dp_SigmaOut(287);
  start_cp_LambdaIn(288) <= start_dp_SigmaOut(288);
  start_cp_LambdaIn(289) <= start_dp_SigmaOut(289);
  start_cp_LambdaIn(290) <= start_dp_SigmaOut(290);
  start_cp_LambdaIn(291) <= start_dp_SigmaOut(291);
  start_cp_LambdaIn(292) <= start_dp_SigmaOut(292);

  start_dp_SigmaIn(1) <= start_cp_LambdaOut(1);
  start_dp_SigmaIn(2) <= start_cp_LambdaOut(2);
  start_dp_SigmaIn(3) <= start_cp_LambdaOut(3);
  start_dp_SigmaIn(4) <= start_cp_LambdaOut(4);
  start_dp_SigmaIn(5) <= start_cp_LambdaOut(5);
  start_dp_SigmaIn(6) <= start_cp_LambdaOut(6);
  start_dp_SigmaIn(7) <= start_cp_LambdaOut(7);
  start_dp_SigmaIn(8) <= start_cp_LambdaOut(8);
  start_dp_SigmaIn(9) <= start_cp_LambdaOut(9);
  start_dp_SigmaIn(10) <= start_cp_LambdaOut(10);
  start_dp_SigmaIn(11) <= start_cp_LambdaOut(11);
  start_dp_SigmaIn(12) <= start_cp_LambdaOut(12);
  start_dp_SigmaIn(13) <= start_cp_LambdaOut(13);
  start_dp_SigmaIn(14) <= start_cp_LambdaOut(14);
  start_dp_SigmaIn(15) <= start_cp_LambdaOut(15);
  start_dp_SigmaIn(16) <= start_cp_LambdaOut(16);
  start_dp_SigmaIn(17) <= start_cp_LambdaOut(17);
  start_dp_SigmaIn(18) <= start_cp_LambdaOut(18);
  start_dp_SigmaIn(19) <= start_cp_LambdaOut(19);
  start_dp_SigmaIn(20) <= start_cp_LambdaOut(20);
  start_dp_SigmaIn(21) <= start_cp_LambdaOut(21);
  start_dp_SigmaIn(22) <= start_cp_LambdaOut(22);
  start_dp_SigmaIn(23) <= start_cp_LambdaOut(23);
  start_dp_SigmaIn(24) <= start_cp_LambdaOut(24);
  start_dp_SigmaIn(25) <= start_cp_LambdaOut(25);
  start_dp_SigmaIn(26) <= start_cp_LambdaOut(26);
  start_dp_SigmaIn(27) <= start_cp_LambdaOut(27);
  start_dp_SigmaIn(28) <= start_cp_LambdaOut(28);
  start_dp_SigmaIn(29) <= start_cp_LambdaOut(29);
  start_dp_SigmaIn(30) <= start_cp_LambdaOut(30);
  start_dp_SigmaIn(31) <= start_cp_LambdaOut(31);
  start_dp_SigmaIn(32) <= start_cp_LambdaOut(32);
  start_dp_SigmaIn(33) <= start_cp_LambdaOut(33);
  start_dp_SigmaIn(34) <= start_cp_LambdaOut(34);
  start_dp_SigmaIn(35) <= start_cp_LambdaOut(35);
  start_dp_SigmaIn(36) <= start_cp_LambdaOut(36);
  start_dp_SigmaIn(37) <= start_cp_LambdaOut(37);
  start_dp_SigmaIn(38) <= start_cp_LambdaOut(38);
  start_dp_SigmaIn(39) <= start_cp_LambdaOut(39);
  start_dp_SigmaIn(40) <= start_cp_LambdaOut(40);
  start_dp_SigmaIn(41) <= start_cp_LambdaOut(41);
  start_dp_SigmaIn(42) <= start_cp_LambdaOut(42);
  start_dp_SigmaIn(43) <= start_cp_LambdaOut(43);
  start_dp_SigmaIn(44) <= start_cp_LambdaOut(44);
  start_dp_SigmaIn(45) <= start_cp_LambdaOut(45);
  start_dp_SigmaIn(46) <= start_cp_LambdaOut(46);
  start_dp_SigmaIn(47) <= start_cp_LambdaOut(47);
  start_dp_SigmaIn(48) <= start_cp_LambdaOut(48);
  start_dp_SigmaIn(49) <= start_cp_LambdaOut(49);
  start_dp_SigmaIn(50) <= start_cp_LambdaOut(50);
  start_dp_SigmaIn(51) <= start_cp_LambdaOut(51);
  start_dp_SigmaIn(52) <= start_cp_LambdaOut(52);
  start_dp_SigmaIn(53) <= start_cp_LambdaOut(53);
  start_dp_SigmaIn(54) <= start_cp_LambdaOut(54);
  start_dp_SigmaIn(55) <= start_cp_LambdaOut(55);
  start_dp_SigmaIn(56) <= start_cp_LambdaOut(56);
  start_dp_SigmaIn(57) <= start_cp_LambdaOut(57);
  start_dp_SigmaIn(58) <= start_cp_LambdaOut(58);
  start_dp_SigmaIn(59) <= start_cp_LambdaOut(59);
  start_dp_SigmaIn(60) <= start_cp_LambdaOut(60);
  start_dp_SigmaIn(61) <= start_cp_LambdaOut(61);
  start_dp_SigmaIn(62) <= start_cp_LambdaOut(62);
  start_dp_SigmaIn(63) <= start_cp_LambdaOut(63);
  start_dp_SigmaIn(64) <= start_cp_LambdaOut(64);
  start_dp_SigmaIn(65) <= start_cp_LambdaOut(65);
  start_dp_SigmaIn(66) <= start_cp_LambdaOut(66);
  start_dp_SigmaIn(67) <= start_cp_LambdaOut(67);
  start_dp_SigmaIn(68) <= start_cp_LambdaOut(68);
  start_dp_SigmaIn(69) <= start_cp_LambdaOut(69);
  start_dp_SigmaIn(70) <= start_cp_LambdaOut(70);
  start_dp_SigmaIn(71) <= start_cp_LambdaOut(71);
  start_dp_SigmaIn(72) <= start_cp_LambdaOut(72);
  start_dp_SigmaIn(73) <= start_cp_LambdaOut(73);
  start_dp_SigmaIn(74) <= start_cp_LambdaOut(74);
  start_dp_SigmaIn(75) <= start_cp_LambdaOut(75);
  start_dp_SigmaIn(76) <= start_cp_LambdaOut(76);
  start_dp_SigmaIn(77) <= start_cp_LambdaOut(77);
  start_dp_SigmaIn(78) <= start_cp_LambdaOut(78);
  start_dp_SigmaIn(79) <= start_cp_LambdaOut(79);
  start_dp_SigmaIn(80) <= start_cp_LambdaOut(80);
  start_dp_SigmaIn(81) <= start_cp_LambdaOut(81);
  start_dp_SigmaIn(82) <= start_cp_LambdaOut(82);
  start_dp_SigmaIn(83) <= start_cp_LambdaOut(83);
  start_dp_SigmaIn(84) <= start_cp_LambdaOut(84);
  start_dp_SigmaIn(85) <= start_cp_LambdaOut(85);
  start_dp_SigmaIn(86) <= start_cp_LambdaOut(86);
  start_dp_SigmaIn(87) <= start_cp_LambdaOut(87);
  start_dp_SigmaIn(88) <= start_cp_LambdaOut(88);
  start_dp_SigmaIn(89) <= start_cp_LambdaOut(89);
  start_dp_SigmaIn(90) <= start_cp_LambdaOut(90);
  start_dp_SigmaIn(91) <= start_cp_LambdaOut(91);
  start_dp_SigmaIn(92) <= start_cp_LambdaOut(92);
  start_dp_SigmaIn(93) <= start_cp_LambdaOut(93);
  start_dp_SigmaIn(94) <= start_cp_LambdaOut(94);
  start_dp_SigmaIn(95) <= start_cp_LambdaOut(95);
  start_dp_SigmaIn(96) <= start_cp_LambdaOut(96);
  start_dp_SigmaIn(97) <= start_cp_LambdaOut(97);
  start_dp_SigmaIn(98) <= start_cp_LambdaOut(98);
  start_dp_SigmaIn(99) <= start_cp_LambdaOut(99);
  start_dp_SigmaIn(100) <= start_cp_LambdaOut(100);
  start_dp_SigmaIn(101) <= start_cp_LambdaOut(101);
  start_dp_SigmaIn(102) <= start_cp_LambdaOut(102);
  start_dp_SigmaIn(103) <= start_cp_LambdaOut(103);
  start_dp_SigmaIn(104) <= start_cp_LambdaOut(104);
  start_dp_SigmaIn(105) <= start_cp_LambdaOut(105);
  start_dp_SigmaIn(106) <= start_cp_LambdaOut(106);
  start_dp_SigmaIn(107) <= start_cp_LambdaOut(107);
  start_dp_SigmaIn(108) <= start_cp_LambdaOut(108);
  start_dp_SigmaIn(109) <= start_cp_LambdaOut(109);
  start_dp_SigmaIn(110) <= start_cp_LambdaOut(110);
  start_dp_SigmaIn(111) <= start_cp_LambdaOut(111);
  start_dp_SigmaIn(112) <= start_cp_LambdaOut(112);
  start_dp_SigmaIn(113) <= start_cp_LambdaOut(113);
  start_dp_SigmaIn(114) <= start_cp_LambdaOut(114);
  start_dp_SigmaIn(115) <= start_cp_LambdaOut(115);
  start_dp_SigmaIn(116) <= start_cp_LambdaOut(116);
  start_dp_SigmaIn(117) <= start_cp_LambdaOut(117);
  start_dp_SigmaIn(118) <= start_cp_LambdaOut(118);
  start_dp_SigmaIn(119) <= start_cp_LambdaOut(119);
  start_dp_SigmaIn(120) <= start_cp_LambdaOut(120);
  start_dp_SigmaIn(121) <= start_cp_LambdaOut(121);
  start_dp_SigmaIn(122) <= start_cp_LambdaOut(122);
  start_dp_SigmaIn(123) <= start_cp_LambdaOut(123);
  start_dp_SigmaIn(124) <= start_cp_LambdaOut(124);
  start_dp_SigmaIn(125) <= start_cp_LambdaOut(125);
  start_dp_SigmaIn(126) <= start_cp_LambdaOut(126);
  start_dp_SigmaIn(127) <= start_cp_LambdaOut(127);
  start_dp_SigmaIn(128) <= start_cp_LambdaOut(128);
  start_dp_SigmaIn(129) <= start_cp_LambdaOut(129);
  start_dp_SigmaIn(130) <= start_cp_LambdaOut(130);
  start_dp_SigmaIn(131) <= start_cp_LambdaOut(131);
  start_dp_SigmaIn(132) <= start_cp_LambdaOut(132);
  start_dp_SigmaIn(133) <= start_cp_LambdaOut(133);
  start_dp_SigmaIn(134) <= start_cp_LambdaOut(134);
  start_dp_SigmaIn(135) <= start_cp_LambdaOut(135);
  start_dp_SigmaIn(136) <= start_cp_LambdaOut(136);
  start_dp_SigmaIn(137) <= start_cp_LambdaOut(137);
  start_dp_SigmaIn(138) <= start_cp_LambdaOut(138);
  start_dp_SigmaIn(139) <= start_cp_LambdaOut(139);
  start_dp_SigmaIn(140) <= start_cp_LambdaOut(140);
  start_dp_SigmaIn(141) <= start_cp_LambdaOut(141);
  start_dp_SigmaIn(142) <= start_cp_LambdaOut(142);
  start_dp_SigmaIn(143) <= start_cp_LambdaOut(143);
  start_dp_SigmaIn(144) <= start_cp_LambdaOut(144);
  start_dp_SigmaIn(145) <= start_cp_LambdaOut(145);
  start_dp_SigmaIn(146) <= start_cp_LambdaOut(146);
  start_dp_SigmaIn(147) <= start_cp_LambdaOut(147);
  start_dp_SigmaIn(148) <= start_cp_LambdaOut(148);
  start_dp_SigmaIn(149) <= start_cp_LambdaOut(149);
  start_dp_SigmaIn(150) <= start_cp_LambdaOut(150);
  start_dp_SigmaIn(151) <= start_cp_LambdaOut(151);
  start_dp_SigmaIn(152) <= start_cp_LambdaOut(152);
  start_dp_SigmaIn(153) <= start_cp_LambdaOut(153);
  start_dp_SigmaIn(154) <= start_cp_LambdaOut(154);
  start_dp_SigmaIn(155) <= start_cp_LambdaOut(155);
  start_dp_SigmaIn(156) <= start_cp_LambdaOut(156);
  start_dp_SigmaIn(157) <= start_cp_LambdaOut(157);
  start_dp_SigmaIn(158) <= start_cp_LambdaOut(158);
  start_dp_SigmaIn(159) <= start_cp_LambdaOut(159);
  start_dp_SigmaIn(160) <= start_cp_LambdaOut(160);
  start_dp_SigmaIn(161) <= start_cp_LambdaOut(161);
  start_dp_SigmaIn(162) <= start_cp_LambdaOut(162);
  start_dp_SigmaIn(163) <= start_cp_LambdaOut(163);
  start_dp_SigmaIn(164) <= start_cp_LambdaOut(164);
  start_dp_SigmaIn(165) <= start_cp_LambdaOut(165);
  start_dp_SigmaIn(166) <= start_cp_LambdaOut(166);
  start_dp_SigmaIn(167) <= start_cp_LambdaOut(167);
  start_dp_SigmaIn(168) <= start_cp_LambdaOut(168);
  start_dp_SigmaIn(169) <= start_cp_LambdaOut(169);
  start_dp_SigmaIn(170) <= start_cp_LambdaOut(170);
  start_dp_SigmaIn(171) <= start_cp_LambdaOut(171);
  start_dp_SigmaIn(172) <= start_cp_LambdaOut(172);
  start_dp_SigmaIn(173) <= start_cp_LambdaOut(173);
  start_dp_SigmaIn(174) <= start_cp_LambdaOut(174);
  start_dp_SigmaIn(175) <= start_cp_LambdaOut(175);
  start_dp_SigmaIn(176) <= start_cp_LambdaOut(176);
  start_dp_SigmaIn(177) <= start_cp_LambdaOut(177);
  start_dp_SigmaIn(178) <= start_cp_LambdaOut(178);
  start_dp_SigmaIn(179) <= start_cp_LambdaOut(179);
  start_dp_SigmaIn(180) <= start_cp_LambdaOut(180);
  start_dp_SigmaIn(181) <= start_cp_LambdaOut(181);
  start_dp_SigmaIn(182) <= start_cp_LambdaOut(182);
  start_dp_SigmaIn(183) <= start_cp_LambdaOut(183);
  start_dp_SigmaIn(184) <= start_cp_LambdaOut(184);
  start_dp_SigmaIn(185) <= start_cp_LambdaOut(185);
  start_dp_SigmaIn(186) <= start_cp_LambdaOut(186);
  start_dp_SigmaIn(187) <= start_cp_LambdaOut(187);
  start_dp_SigmaIn(188) <= start_cp_LambdaOut(188);
  start_dp_SigmaIn(189) <= start_cp_LambdaOut(189);
  start_dp_SigmaIn(190) <= start_cp_LambdaOut(190);
  start_dp_SigmaIn(191) <= start_cp_LambdaOut(191);
  start_dp_SigmaIn(192) <= start_cp_LambdaOut(192);
  start_dp_SigmaIn(193) <= start_cp_LambdaOut(193);
  start_dp_SigmaIn(194) <= start_cp_LambdaOut(194);
  start_dp_SigmaIn(195) <= start_cp_LambdaOut(195);
  start_dp_SigmaIn(196) <= start_cp_LambdaOut(196);
  start_dp_SigmaIn(197) <= start_cp_LambdaOut(197);
  start_dp_SigmaIn(198) <= start_cp_LambdaOut(198);
  start_dp_SigmaIn(199) <= start_cp_LambdaOut(199);
  start_dp_SigmaIn(200) <= start_cp_LambdaOut(200);
  start_dp_SigmaIn(201) <= start_cp_LambdaOut(201);
  start_dp_SigmaIn(202) <= start_cp_LambdaOut(202);
  start_dp_SigmaIn(203) <= start_cp_LambdaOut(203);
  start_dp_SigmaIn(204) <= start_cp_LambdaOut(204);
  start_dp_SigmaIn(205) <= start_cp_LambdaOut(205);
  start_dp_SigmaIn(206) <= start_cp_LambdaOut(206);
  start_dp_SigmaIn(207) <= start_cp_LambdaOut(207);
  start_dp_SigmaIn(208) <= start_cp_LambdaOut(208);
  start_dp_SigmaIn(209) <= start_cp_LambdaOut(209);
  start_dp_SigmaIn(210) <= start_cp_LambdaOut(210);
  start_dp_SigmaIn(211) <= start_cp_LambdaOut(211);
  start_dp_SigmaIn(212) <= start_cp_LambdaOut(212);
  start_dp_SigmaIn(213) <= start_cp_LambdaOut(213);
  start_dp_SigmaIn(214) <= start_cp_LambdaOut(214);
  start_dp_SigmaIn(215) <= start_cp_LambdaOut(215);
  start_dp_SigmaIn(216) <= start_cp_LambdaOut(216);
  start_dp_SigmaIn(217) <= start_cp_LambdaOut(217);
  start_dp_SigmaIn(218) <= start_cp_LambdaOut(218);
  start_dp_SigmaIn(219) <= start_cp_LambdaOut(219);
  start_dp_SigmaIn(220) <= start_cp_LambdaOut(220);
  start_dp_SigmaIn(221) <= start_cp_LambdaOut(221);
  start_dp_SigmaIn(222) <= start_cp_LambdaOut(222);
  start_dp_SigmaIn(223) <= start_cp_LambdaOut(223);
  start_dp_SigmaIn(224) <= start_cp_LambdaOut(224);
  start_dp_SigmaIn(225) <= start_cp_LambdaOut(225);
  start_dp_SigmaIn(226) <= start_cp_LambdaOut(226);
  start_dp_SigmaIn(227) <= start_cp_LambdaOut(227);
  start_dp_SigmaIn(228) <= start_cp_LambdaOut(228);
  start_dp_SigmaIn(229) <= start_cp_LambdaOut(229);
  start_dp_SigmaIn(230) <= start_cp_LambdaOut(230);
  start_dp_SigmaIn(231) <= start_cp_LambdaOut(231);
  start_dp_SigmaIn(232) <= start_cp_LambdaOut(232);
  start_dp_SigmaIn(233) <= start_cp_LambdaOut(233);
  start_dp_SigmaIn(234) <= start_cp_LambdaOut(234);
  start_dp_SigmaIn(235) <= start_cp_LambdaOut(235);
  start_dp_SigmaIn(236) <= start_cp_LambdaOut(236);
  start_dp_SigmaIn(237) <= start_cp_LambdaOut(237);
  start_dp_SigmaIn(238) <= start_cp_LambdaOut(238);
  start_dp_SigmaIn(239) <= start_cp_LambdaOut(239);
  start_dp_SigmaIn(240) <= start_cp_LambdaOut(240);
  start_dp_SigmaIn(241) <= start_cp_LambdaOut(241);
  start_dp_SigmaIn(242) <= start_cp_LambdaOut(242);
  start_dp_SigmaIn(243) <= start_cp_LambdaOut(243);
  start_dp_SigmaIn(244) <= start_cp_LambdaOut(244);
  start_dp_SigmaIn(245) <= start_cp_LambdaOut(245);
  start_dp_SigmaIn(246) <= start_cp_LambdaOut(246);
  start_dp_SigmaIn(247) <= start_cp_LambdaOut(247);
  start_dp_SigmaIn(248) <= start_cp_LambdaOut(248);
  start_dp_SigmaIn(249) <= start_cp_LambdaOut(249);
  start_dp_SigmaIn(250) <= start_cp_LambdaOut(250);
  start_dp_SigmaIn(251) <= start_cp_LambdaOut(251);
  start_dp_SigmaIn(252) <= start_cp_LambdaOut(252);
  start_dp_SigmaIn(253) <= start_cp_LambdaOut(253);
  start_dp_SigmaIn(254) <= start_cp_LambdaOut(254);
  start_dp_SigmaIn(255) <= start_cp_LambdaOut(255);
  start_dp_SigmaIn(256) <= start_cp_LambdaOut(256);
  start_dp_SigmaIn(257) <= start_cp_LambdaOut(257);
  start_dp_SigmaIn(258) <= start_cp_LambdaOut(258);
  start_dp_SigmaIn(259) <= start_cp_LambdaOut(259);
  start_dp_SigmaIn(260) <= start_cp_LambdaOut(260);
  start_dp_SigmaIn(261) <= start_cp_LambdaOut(261);
  start_dp_SigmaIn(262) <= start_cp_LambdaOut(262);
  start_dp_SigmaIn(263) <= start_cp_LambdaOut(263);
  start_dp_SigmaIn(264) <= start_cp_LambdaOut(264);
  start_dp_SigmaIn(265) <= start_cp_LambdaOut(265);
  start_dp_SigmaIn(266) <= start_cp_LambdaOut(266);
  start_dp_SigmaIn(267) <= start_cp_LambdaOut(267);
  start_dp_SigmaIn(268) <= start_cp_LambdaOut(268);
  start_dp_SigmaIn(269) <= start_cp_LambdaOut(269);
  start_dp_SigmaIn(270) <= start_cp_LambdaOut(270);
  start_dp_SigmaIn(271) <= start_cp_LambdaOut(271);
  start_dp_SigmaIn(272) <= start_cp_LambdaOut(272);
  start_dp_SigmaIn(273) <= start_cp_LambdaOut(273);
  start_dp_SigmaIn(274) <= start_cp_LambdaOut(274);
  start_dp_SigmaIn(275) <= start_cp_LambdaOut(275);
  start_dp_SigmaIn(276) <= start_cp_LambdaOut(276);
  start_dp_SigmaIn(277) <= start_cp_LambdaOut(277);
  start_dp_SigmaIn(278) <= start_cp_LambdaOut(278);
  start_dp_SigmaIn(279) <= start_cp_LambdaOut(279);
  start_dp_SigmaIn(280) <= start_cp_LambdaOut(280);
  start_dp_SigmaIn(281) <= start_cp_LambdaOut(281);
  start_dp_SigmaIn(282) <= start_cp_LambdaOut(282);
  start_dp_SigmaIn(283) <= start_cp_LambdaOut(283);
  start_dp_SigmaIn(284) <= start_cp_LambdaOut(284);
  start_dp_SigmaIn(285) <= start_cp_LambdaOut(285);
  start_dp_SigmaIn(286) <= start_cp_LambdaOut(286);
  start_dp_SigmaIn(287) <= start_cp_LambdaOut(287);
  start_dp_SigmaIn(288) <= start_cp_LambdaOut(288);
  start_dp_SigmaIn(289) <= start_cp_LambdaOut(289);
  start_dp_SigmaIn(290) <= start_cp_LambdaOut(290);
  start_dp_SigmaIn(291) <= start_cp_LambdaOut(291);
  start_dp_SigmaIn(292) <= start_cp_LambdaOut(292);
  start_dp_SigmaIn(293) <= start_cp_LambdaOut(293);
  start_dp_SigmaIn(294) <= start_cp_LambdaOut(294);
end default_arch;