entity start_ln is
  port(

    omega_ip : in bit_vector(2 downto 1);
    start_cp_ip : in bit_vector(278 downto 1);
    start_dp_ip : in bit_vector(273 downto 1);
    omega_op : out bit_vector(2 downto 1) := (others => '0');
    start_cp_op : out bit_vector(275 downto 1) := (others => '0');
    start_dp_op : out bit_vector(276 downto 1) := (others => '0');

    reset : in bit;
    clk   : in bit);
end start_ln;

architecture Behavioral of start_ln is 

begin

  omega_op(1) <= start_cp_ip(1);
  omega_op(2) <= start_cp_ip(125);

  start_cp_op(1) <= omega_ip(1);
  start_cp_op(2) <= start_dp_ip(1);
  start_cp_op(3) <= start_dp_ip(2);
  start_cp_op(4) <= start_dp_ip(3);
  start_cp_op(5) <= start_dp_ip(4);
  start_cp_op(6) <= start_dp_ip(5);
  start_cp_op(7) <= start_dp_ip(6);
  start_cp_op(8) <= start_dp_ip(7);
  start_cp_op(9) <= start_dp_ip(8);
  start_cp_op(10) <= start_dp_ip(9);
  start_cp_op(11) <= start_dp_ip(10);
  start_cp_op(12) <= start_dp_ip(11);
  start_cp_op(13) <= start_dp_ip(12);
  start_cp_op(14) <= start_dp_ip(13);
  start_cp_op(15) <= start_dp_ip(14);
  start_cp_op(16) <= start_dp_ip(15);
  start_cp_op(17) <= start_dp_ip(16);
  start_cp_op(18) <= start_dp_ip(17);
  start_cp_op(19) <= start_dp_ip(18);
  start_cp_op(20) <= start_dp_ip(19);
  start_cp_op(21) <= start_dp_ip(20);
  start_cp_op(22) <= start_dp_ip(21);
  start_cp_op(23) <= start_dp_ip(22);
  start_cp_op(24) <= start_dp_ip(23);
  start_cp_op(25) <= start_dp_ip(24);
  start_cp_op(26) <= start_dp_ip(25);
  start_cp_op(27) <= start_dp_ip(26);
  start_cp_op(28) <= start_dp_ip(27);
  start_cp_op(29) <= start_dp_ip(28);
  start_cp_op(30) <= start_dp_ip(29);
  start_cp_op(31) <= start_dp_ip(30);
  start_cp_op(32) <= start_dp_ip(31);
  start_cp_op(33) <= start_dp_ip(32);
  start_cp_op(34) <= start_dp_ip(33);
  start_cp_op(35) <= start_dp_ip(34);
  start_cp_op(36) <= start_dp_ip(35);
  start_cp_op(37) <= start_dp_ip(36);
  start_cp_op(38) <= start_dp_ip(37);
  start_cp_op(39) <= start_dp_ip(38);
  start_cp_op(40) <= start_dp_ip(39);
  start_cp_op(41) <= start_dp_ip(40);
  start_cp_op(42) <= start_dp_ip(41);
  start_cp_op(43) <= start_dp_ip(42);
  start_cp_op(44) <= start_dp_ip(43);
  start_cp_op(45) <= start_dp_ip(44);
  start_cp_op(46) <= start_dp_ip(45);
  start_cp_op(47) <= start_dp_ip(46);
  start_cp_op(48) <= start_dp_ip(47);
  start_cp_op(49) <= start_dp_ip(48);
  start_cp_op(50) <= start_dp_ip(49);
  start_cp_op(51) <= start_dp_ip(50);
  start_cp_op(52) <= start_dp_ip(51);
  start_cp_op(53) <= start_dp_ip(52);
  start_cp_op(54) <= start_dp_ip(53);
  start_cp_op(55) <= start_dp_ip(54);
  start_cp_op(56) <= start_dp_ip(55);
  start_cp_op(57) <= start_dp_ip(56);
  start_cp_op(58) <= start_dp_ip(57);
  start_cp_op(59) <= start_dp_ip(58);
  start_cp_op(60) <= start_dp_ip(59);
  start_cp_op(61) <= start_dp_ip(60);
  start_cp_op(62) <= start_dp_ip(61);
  start_cp_op(63) <= start_dp_ip(62);
  start_cp_op(64) <= start_dp_ip(63);
  start_cp_op(65) <= start_dp_ip(64);
  start_cp_op(66) <= start_dp_ip(65);
  start_cp_op(67) <= start_dp_ip(66);
  start_cp_op(68) <= start_dp_ip(67);
  start_cp_op(69) <= start_dp_ip(68);
  start_cp_op(70) <= start_dp_ip(69);
  start_cp_op(71) <= start_dp_ip(70);
  start_cp_op(72) <= start_dp_ip(71);
  start_cp_op(73) <= start_dp_ip(72);
  start_cp_op(74) <= start_dp_ip(73);
  start_cp_op(75) <= start_dp_ip(74);
  start_cp_op(76) <= start_dp_ip(75);
  start_cp_op(77) <= start_dp_ip(76);
  start_cp_op(78) <= start_dp_ip(77);
  start_cp_op(79) <= start_dp_ip(78);
  start_cp_op(80) <= start_dp_ip(79);
  start_cp_op(81) <= start_dp_ip(80);
  start_cp_op(82) <= start_dp_ip(81);
  start_cp_op(83) <= start_dp_ip(82);
  start_cp_op(84) <= start_dp_ip(83);
  start_cp_op(85) <= start_dp_ip(84);
  start_cp_op(86) <= start_dp_ip(85);
  start_cp_op(87) <= start_dp_ip(86);
  start_cp_op(88) <= start_dp_ip(87);
  start_cp_op(89) <= start_dp_ip(88);
  start_cp_op(90) <= start_dp_ip(89);
  start_cp_op(91) <= start_dp_ip(90);
  start_cp_op(92) <= start_dp_ip(91);
  start_cp_op(93) <= start_dp_ip(92);
  start_cp_op(94) <= start_dp_ip(93);
  start_cp_op(95) <= start_dp_ip(94);
  start_cp_op(96) <= start_dp_ip(95);
  start_cp_op(97) <= start_dp_ip(96);
  start_cp_op(98) <= start_dp_ip(97);
  start_cp_op(99) <= start_dp_ip(98);
  start_cp_op(100) <= start_dp_ip(99);
  start_cp_op(101) <= start_dp_ip(100);
  start_cp_op(102) <= start_dp_ip(101);
  start_cp_op(103) <= start_dp_ip(102);
  start_cp_op(104) <= start_dp_ip(103);
  start_cp_op(105) <= start_dp_ip(104);
  start_cp_op(106) <= start_dp_ip(105);
  start_cp_op(107) <= start_dp_ip(106);
  start_cp_op(108) <= start_dp_ip(107);
  start_cp_op(109) <= start_dp_ip(108);
  start_cp_op(110) <= start_dp_ip(109);
  start_cp_op(111) <= start_dp_ip(110);
  start_cp_op(112) <= start_dp_ip(111);
  start_cp_op(113) <= start_dp_ip(112);
  start_cp_op(114) <= start_dp_ip(113);
  start_cp_op(115) <= start_dp_ip(114);
  start_cp_op(116) <= start_dp_ip(115);
  start_cp_op(117) <= start_dp_ip(116);
  start_cp_op(118) <= start_dp_ip(117);
  start_cp_op(119) <= start_dp_ip(118);
  start_cp_op(120) <= omega_ip(2);
  start_cp_op(121) <= start_dp_ip(119);
  start_cp_op(122) <= start_dp_ip(120);
  start_cp_op(123) <= start_dp_ip(121);
  start_cp_op(124) <= start_dp_ip(122);
  start_cp_op(125) <= start_dp_ip(123);
  start_cp_op(126) <= start_dp_ip(124);
  start_cp_op(127) <= start_dp_ip(125);
  start_cp_op(128) <= start_dp_ip(126);
  start_cp_op(129) <= start_dp_ip(127);
  start_cp_op(130) <= start_dp_ip(128);
  start_cp_op(131) <= start_dp_ip(129);
  start_cp_op(132) <= start_dp_ip(130);
  start_cp_op(133) <= start_dp_ip(131);
  start_cp_op(134) <= start_dp_ip(132);
  start_cp_op(135) <= start_dp_ip(133);
  start_cp_op(136) <= start_dp_ip(134);
  start_cp_op(137) <= start_dp_ip(135);
  start_cp_op(138) <= start_dp_ip(136);
  start_cp_op(139) <= start_dp_ip(137);
  start_cp_op(140) <= start_dp_ip(138);
  start_cp_op(141) <= start_dp_ip(139);
  start_cp_op(142) <= start_dp_ip(140);
  start_cp_op(143) <= start_dp_ip(141);
  start_cp_op(144) <= start_dp_ip(142);
  start_cp_op(145) <= start_dp_ip(143);
  start_cp_op(146) <= start_dp_ip(144);
  start_cp_op(147) <= start_dp_ip(145);
  start_cp_op(148) <= start_dp_ip(146);
  start_cp_op(149) <= start_dp_ip(147);
  start_cp_op(150) <= start_dp_ip(148);
  start_cp_op(151) <= start_dp_ip(149);
  start_cp_op(152) <= start_dp_ip(150);
  start_cp_op(153) <= start_dp_ip(151);
  start_cp_op(154) <= start_dp_ip(152);
  start_cp_op(155) <= start_dp_ip(153);
  start_cp_op(156) <= start_dp_ip(154);
  start_cp_op(157) <= start_dp_ip(155);
  start_cp_op(158) <= start_dp_ip(156);
  start_cp_op(159) <= start_dp_ip(157);
  start_cp_op(160) <= start_dp_ip(158);
  start_cp_op(161) <= start_dp_ip(159);
  start_cp_op(162) <= start_dp_ip(160);
  start_cp_op(163) <= start_dp_ip(161);
  start_cp_op(164) <= start_dp_ip(162);
  start_cp_op(165) <= start_dp_ip(163);
  start_cp_op(166) <= start_dp_ip(164);
  start_cp_op(167) <= start_dp_ip(165);
  start_cp_op(168) <= start_dp_ip(166);
  start_cp_op(169) <= start_dp_ip(167);
  start_cp_op(170) <= start_dp_ip(168);
  start_cp_op(171) <= start_dp_ip(169);
  start_cp_op(172) <= start_dp_ip(170);
  start_cp_op(173) <= start_dp_ip(171);
  start_cp_op(174) <= start_dp_ip(172);
  start_cp_op(175) <= start_dp_ip(173);
  start_cp_op(176) <= start_dp_ip(174);
  start_cp_op(177) <= start_dp_ip(175);
  start_cp_op(178) <= start_dp_ip(176);
  start_cp_op(179) <= start_dp_ip(177);
  start_cp_op(180) <= start_dp_ip(178);
  start_cp_op(181) <= start_dp_ip(179);
  start_cp_op(182) <= start_dp_ip(180);
  start_cp_op(183) <= start_dp_ip(181);
  start_cp_op(184) <= start_dp_ip(182);
  start_cp_op(185) <= start_dp_ip(183);
  start_cp_op(186) <= start_dp_ip(184);
  start_cp_op(187) <= start_dp_ip(185);
  start_cp_op(188) <= start_dp_ip(186);
  start_cp_op(189) <= start_dp_ip(187);
  start_cp_op(190) <= start_dp_ip(188);
  start_cp_op(191) <= start_dp_ip(189);
  start_cp_op(192) <= start_dp_ip(190);
  start_cp_op(193) <= start_dp_ip(191);
  start_cp_op(194) <= start_dp_ip(192);
  start_cp_op(195) <= start_dp_ip(193);
  start_cp_op(196) <= start_dp_ip(194);
  start_cp_op(197) <= start_dp_ip(195);
  start_cp_op(198) <= start_dp_ip(196);
  start_cp_op(199) <= start_dp_ip(197);
  start_cp_op(200) <= start_dp_ip(198);
  start_cp_op(201) <= start_dp_ip(199);
  start_cp_op(202) <= start_dp_ip(200);
  start_cp_op(203) <= start_dp_ip(201);
  start_cp_op(204) <= start_dp_ip(202);
  start_cp_op(205) <= start_dp_ip(203);
  start_cp_op(206) <= start_dp_ip(204);
  start_cp_op(207) <= start_dp_ip(205);
  start_cp_op(208) <= start_dp_ip(206);
  start_cp_op(209) <= start_dp_ip(207);
  start_cp_op(210) <= start_dp_ip(208);
  start_cp_op(211) <= start_dp_ip(209);
  start_cp_op(212) <= start_dp_ip(210);
  start_cp_op(213) <= start_dp_ip(211);
  start_cp_op(214) <= start_dp_ip(212);
  start_cp_op(215) <= start_dp_ip(213);
  start_cp_op(216) <= start_dp_ip(214);
  start_cp_op(217) <= start_dp_ip(215);
  start_cp_op(218) <= start_dp_ip(216);
  start_cp_op(219) <= start_dp_ip(217);
  start_cp_op(220) <= start_dp_ip(218);
  start_cp_op(221) <= start_dp_ip(219);
  start_cp_op(222) <= start_dp_ip(220);
  start_cp_op(223) <= start_dp_ip(221);
  start_cp_op(224) <= start_dp_ip(222);
  start_cp_op(225) <= start_dp_ip(223);
  start_cp_op(226) <= start_dp_ip(224);
  start_cp_op(227) <= start_dp_ip(225);
  start_cp_op(228) <= start_dp_ip(226);
  start_cp_op(229) <= start_dp_ip(227);
  start_cp_op(230) <= start_dp_ip(228);
  start_cp_op(231) <= start_dp_ip(229);
  start_cp_op(232) <= start_dp_ip(230);
  start_cp_op(233) <= start_dp_ip(231);
  start_cp_op(234) <= start_dp_ip(232);
  start_cp_op(235) <= start_dp_ip(233);
  start_cp_op(236) <= start_dp_ip(234);
  start_cp_op(237) <= start_dp_ip(235);
  start_cp_op(238) <= start_dp_ip(236);
  start_cp_op(239) <= start_dp_ip(237);
  start_cp_op(240) <= start_dp_ip(238);
  start_cp_op(241) <= start_dp_ip(239);
  start_cp_op(242) <= start_dp_ip(240);
  start_cp_op(243) <= start_dp_ip(241);
  start_cp_op(244) <= start_dp_ip(242);
  start_cp_op(245) <= start_dp_ip(243);
  start_cp_op(246) <= start_dp_ip(244);
  start_cp_op(247) <= start_dp_ip(245);
  start_cp_op(248) <= start_dp_ip(246);
  start_cp_op(249) <= start_dp_ip(247);
  start_cp_op(250) <= start_dp_ip(248);
  start_cp_op(251) <= start_dp_ip(249);
  start_cp_op(252) <= start_dp_ip(250);
  start_cp_op(253) <= start_dp_ip(251);
  start_cp_op(254) <= start_dp_ip(252);
  start_cp_op(255) <= start_dp_ip(253);
  start_cp_op(256) <= start_dp_ip(254);
  start_cp_op(257) <= start_dp_ip(255);
  start_cp_op(258) <= start_dp_ip(256);
  start_cp_op(259) <= start_dp_ip(257);
  start_cp_op(260) <= start_dp_ip(258);
  start_cp_op(261) <= start_dp_ip(259);
  start_cp_op(262) <= start_dp_ip(260);
  start_cp_op(263) <= start_dp_ip(261);
  start_cp_op(264) <= start_dp_ip(262);
  start_cp_op(265) <= start_dp_ip(263);
  start_cp_op(266) <= start_dp_ip(264);
  start_cp_op(267) <= start_dp_ip(265);
  start_cp_op(268) <= start_dp_ip(266);
  start_cp_op(269) <= start_dp_ip(267);
  start_cp_op(270) <= start_dp_ip(268);
  start_cp_op(271) <= start_dp_ip(269);
  start_cp_op(272) <= start_dp_ip(270);
  start_cp_op(273) <= start_dp_ip(271);
  start_cp_op(274) <= start_dp_ip(272);
  start_cp_op(275) <= start_dp_ip(273);

  start_dp_op(1) <= start_cp_ip(2);
  start_dp_op(2) <= start_cp_ip(3);
  start_dp_op(3) <= start_cp_ip(4);
  start_dp_op(4) <= start_cp_ip(5);
  start_dp_op(5) <= start_cp_ip(6);
  start_dp_op(6) <= start_cp_ip(7);
  start_dp_op(7) <= start_cp_ip(9);
  start_dp_op(8) <= start_cp_ip(8);
  start_dp_op(9) <= start_cp_ip(11);
  start_dp_op(10) <= start_cp_ip(10);
  start_dp_op(11) <= start_cp_ip(12);
  start_dp_op(12) <= start_cp_ip(13);
  start_dp_op(13) <= start_cp_ip(14);
  start_dp_op(14) <= start_cp_ip(15);
  start_dp_op(15) <= start_cp_ip(16);
  start_dp_op(16) <= start_cp_ip(17);
  start_dp_op(17) <= start_cp_ip(18);
  start_dp_op(18) <= start_cp_ip(19);
  start_dp_op(19) <= start_cp_ip(20);
  start_dp_op(20) <= start_cp_ip(21);
  start_dp_op(21) <= start_cp_ip(22);
  start_dp_op(22) <= start_cp_ip(23);
  start_dp_op(23) <= start_cp_ip(25);
  start_dp_op(24) <= start_cp_ip(24);
  start_dp_op(25) <= start_cp_ip(26);
  start_dp_op(26) <= start_cp_ip(27);
  start_dp_op(27) <= start_cp_ip(28);
  start_dp_op(28) <= start_cp_ip(29);
  start_dp_op(29) <= start_cp_ip(30);
  start_dp_op(30) <= start_cp_ip(31);
  start_dp_op(31) <= start_cp_ip(32);
  start_dp_op(32) <= start_cp_ip(33);
  start_dp_op(33) <= start_cp_ip(34);
  start_dp_op(34) <= start_cp_ip(35);
  start_dp_op(35) <= start_cp_ip(36);
  start_dp_op(36) <= start_cp_ip(37);
  start_dp_op(37) <= start_cp_ip(38);
  start_dp_op(38) <= start_cp_ip(39);
  start_dp_op(39) <= start_cp_ip(40);
  start_dp_op(40) <= start_cp_ip(41);
  start_dp_op(41) <= start_cp_ip(42);
  start_dp_op(42) <= start_cp_ip(44);
  start_dp_op(43) <= start_cp_ip(43);
  start_dp_op(44) <= start_cp_ip(46);
  start_dp_op(45) <= start_cp_ip(45);
  start_dp_op(46) <= start_cp_ip(48);
  start_dp_op(47) <= start_cp_ip(47);
  start_dp_op(48) <= start_cp_ip(49);
  start_dp_op(49) <= start_cp_ip(50);
  start_dp_op(50) <= start_cp_ip(51);
  start_dp_op(51) <= start_cp_ip(52);
  start_dp_op(52) <= start_cp_ip(54);
  start_dp_op(53) <= start_cp_ip(53);
  start_dp_op(54) <= start_cp_ip(56);
  start_dp_op(55) <= start_cp_ip(55);
  start_dp_op(56) <= start_cp_ip(57);
  start_dp_op(57) <= start_cp_ip(58);
  start_dp_op(58) <= start_cp_ip(59);
  start_dp_op(59) <= start_cp_ip(60);
  start_dp_op(60) <= start_cp_ip(61);
  start_dp_op(61) <= start_cp_ip(62);
  start_dp_op(62) <= start_cp_ip(64);
  start_dp_op(63) <= start_cp_ip(63);
  start_dp_op(64) <= start_cp_ip(66);
  start_dp_op(65) <= start_cp_ip(65);
  start_dp_op(66) <= start_cp_ip(67);
  start_dp_op(67) <= start_cp_ip(68);
  start_dp_op(68) <= start_cp_ip(69);
  start_dp_op(69) <= start_cp_ip(70);
  start_dp_op(70) <= start_cp_ip(71);
  start_dp_op(71) <= start_cp_ip(72);
  start_dp_op(72) <= start_cp_ip(73);
  start_dp_op(73) <= start_cp_ip(74);
  start_dp_op(74) <= start_cp_ip(75);
  start_dp_op(75) <= start_cp_ip(76);
  start_dp_op(76) <= start_cp_ip(77);
  start_dp_op(77) <= start_cp_ip(78);
  start_dp_op(78) <= start_cp_ip(80);
  start_dp_op(79) <= start_cp_ip(79);
  start_dp_op(80) <= start_cp_ip(82);
  start_dp_op(81) <= start_cp_ip(81);
  start_dp_op(82) <= start_cp_ip(83);
  start_dp_op(83) <= start_cp_ip(84);
  start_dp_op(84) <= start_cp_ip(85);
  start_dp_op(85) <= start_cp_ip(86);
  start_dp_op(86) <= start_cp_ip(87);
  start_dp_op(87) <= start_cp_ip(88);
  start_dp_op(88) <= start_cp_ip(89);
  start_dp_op(89) <= start_cp_ip(90);
  start_dp_op(90) <= start_cp_ip(91);
  start_dp_op(91) <= start_cp_ip(92);
  start_dp_op(92) <= start_cp_ip(93);
  start_dp_op(93) <= start_cp_ip(94);
  start_dp_op(94) <= start_cp_ip(95);
  start_dp_op(95) <= start_cp_ip(96);
  start_dp_op(96) <= start_cp_ip(97);
  start_dp_op(97) <= start_cp_ip(98);
  start_dp_op(98) <= start_cp_ip(99);
  start_dp_op(99) <= start_cp_ip(100);
  start_dp_op(100) <= start_cp_ip(102);
  start_dp_op(101) <= start_cp_ip(101);
  start_dp_op(102) <= start_cp_ip(104);
  start_dp_op(103) <= start_cp_ip(103);
  start_dp_op(104) <= start_cp_ip(105);
  start_dp_op(105) <= start_cp_ip(106);
  start_dp_op(106) <= start_cp_ip(107);
  start_dp_op(107) <= start_cp_ip(108);
  start_dp_op(108) <= start_cp_ip(109);
  start_dp_op(109) <= start_cp_ip(110);
  start_dp_op(110) <= start_cp_ip(111);
  start_dp_op(111) <= start_cp_ip(113);
  start_dp_op(112) <= start_cp_ip(112);
  start_dp_op(113) <= start_cp_ip(114);
  start_dp_op(114) <= start_cp_ip(115);
  start_dp_op(115) <= start_cp_ip(116);
  start_dp_op(116) <= start_cp_ip(117);
  start_dp_op(117) <= start_cp_ip(118);
  start_dp_op(118) <= start_cp_ip(119);
  start_dp_op(119) <= start_cp_ip(120);
  start_dp_op(120) <= start_cp_ip(121);
  start_dp_op(121) <= start_cp_ip(122);
  start_dp_op(122) <= start_cp_ip(123);
  start_dp_op(123) <= start_cp_ip(124);
  start_dp_op(124) <= start_cp_ip(126);
  start_dp_op(125) <= start_cp_ip(127);
  start_dp_op(126) <= start_cp_ip(128);
  start_dp_op(127) <= start_cp_ip(129);
  start_dp_op(128) <= start_cp_ip(130);
  start_dp_op(129) <= start_cp_ip(131);
  start_dp_op(130) <= start_cp_ip(133);
  start_dp_op(131) <= start_cp_ip(132);
  start_dp_op(132) <= start_cp_ip(134);
  start_dp_op(133) <= start_cp_ip(135);
  start_dp_op(134) <= start_cp_ip(136);
  start_dp_op(135) <= start_cp_ip(137);
  start_dp_op(136) <= start_cp_ip(138);
  start_dp_op(137) <= start_cp_ip(139);
  start_dp_op(138) <= start_cp_ip(140);
  start_dp_op(139) <= start_cp_ip(141);
  start_dp_op(140) <= start_cp_ip(142);
  start_dp_op(141) <= start_cp_ip(143);
  start_dp_op(142) <= start_cp_ip(144);
  start_dp_op(143) <= start_cp_ip(145);
  start_dp_op(144) <= start_cp_ip(146);
  start_dp_op(145) <= start_cp_ip(147);
  start_dp_op(146) <= start_cp_ip(148);
  start_dp_op(147) <= start_cp_ip(149);
  start_dp_op(148) <= start_cp_ip(150);
  start_dp_op(149) <= start_cp_ip(151);
  start_dp_op(150) <= start_cp_ip(152);
  start_dp_op(151) <= start_cp_ip(153);
  start_dp_op(152) <= start_cp_ip(154);
  start_dp_op(153) <= start_cp_ip(156);
  start_dp_op(154) <= start_cp_ip(155);
  start_dp_op(155) <= start_cp_ip(157);
  start_dp_op(156) <= start_cp_ip(159);
  start_dp_op(157) <= start_cp_ip(158);
  start_dp_op(158) <= start_cp_ip(160);
  start_dp_op(159) <= start_cp_ip(161);
  start_dp_op(160) <= start_cp_ip(162);
  start_dp_op(161) <= start_cp_ip(163);
  start_dp_op(162) <= start_cp_ip(164);
  start_dp_op(163) <= start_cp_ip(165);
  start_dp_op(164) <= start_cp_ip(166);
  start_dp_op(165) <= start_cp_ip(167);
  start_dp_op(166) <= start_cp_ip(168);
  start_dp_op(167) <= start_cp_ip(169);
  start_dp_op(168) <= start_cp_ip(170);
  start_dp_op(169) <= start_cp_ip(171);
  start_dp_op(170) <= start_cp_ip(172);
  start_dp_op(171) <= start_cp_ip(173);
  start_dp_op(172) <= start_cp_ip(174);
  start_dp_op(173) <= start_cp_ip(175);
  start_dp_op(174) <= start_cp_ip(176);
  start_dp_op(175) <= start_cp_ip(177);
  start_dp_op(176) <= start_cp_ip(178);
  start_dp_op(177) <= start_cp_ip(179);
  start_dp_op(178) <= start_cp_ip(181);
  start_dp_op(179) <= start_cp_ip(180);
  start_dp_op(180) <= start_cp_ip(183);
  start_dp_op(181) <= start_cp_ip(182);
  start_dp_op(182) <= start_cp_ip(184);
  start_dp_op(183) <= start_cp_ip(185);
  start_dp_op(184) <= start_cp_ip(186);
  start_dp_op(185) <= start_cp_ip(187);
  start_dp_op(186) <= start_cp_ip(188);
  start_dp_op(187) <= start_cp_ip(189);
  start_dp_op(188) <= start_cp_ip(190);
  start_dp_op(189) <= start_cp_ip(191);
  start_dp_op(190) <= start_cp_ip(192);
  start_dp_op(191) <= start_cp_ip(193);
  start_dp_op(192) <= start_cp_ip(194);
  start_dp_op(193) <= start_cp_ip(195);
  start_dp_op(194) <= start_cp_ip(196);
  start_dp_op(195) <= start_cp_ip(197);
  start_dp_op(196) <= start_cp_ip(198);
  start_dp_op(197) <= start_cp_ip(199);
  start_dp_op(198) <= start_cp_ip(200);
  start_dp_op(199) <= start_cp_ip(201);
  start_dp_op(200) <= start_cp_ip(202);
  start_dp_op(201) <= start_cp_ip(203);
  start_dp_op(202) <= start_cp_ip(204);
  start_dp_op(203) <= start_cp_ip(205);
  start_dp_op(204) <= start_cp_ip(206);
  start_dp_op(205) <= start_cp_ip(207);
  start_dp_op(206) <= start_cp_ip(208);
  start_dp_op(207) <= start_cp_ip(209);
  start_dp_op(208) <= start_cp_ip(210);
  start_dp_op(209) <= start_cp_ip(211);
  start_dp_op(210) <= start_cp_ip(212);
  start_dp_op(211) <= start_cp_ip(213);
  start_dp_op(212) <= start_cp_ip(214);
  start_dp_op(213) <= start_cp_ip(215);
  start_dp_op(214) <= start_cp_ip(216);
  start_dp_op(215) <= start_cp_ip(217);
  start_dp_op(216) <= start_cp_ip(218);
  start_dp_op(217) <= start_cp_ip(219);
  start_dp_op(218) <= start_cp_ip(220);
  start_dp_op(219) <= start_cp_ip(222);
  start_dp_op(220) <= start_cp_ip(221);
  start_dp_op(221) <= start_cp_ip(224);
  start_dp_op(222) <= start_cp_ip(223);
  start_dp_op(223) <= start_cp_ip(225);
  start_dp_op(224) <= start_cp_ip(226);
  start_dp_op(225) <= start_cp_ip(227);
  start_dp_op(226) <= start_cp_ip(229);
  start_dp_op(227) <= start_cp_ip(228);
  start_dp_op(228) <= start_cp_ip(230);
  start_dp_op(229) <= start_cp_ip(231);
  start_dp_op(230) <= start_cp_ip(232);
  start_dp_op(231) <= start_cp_ip(233);
  start_dp_op(232) <= start_cp_ip(234);
  start_dp_op(233) <= start_cp_ip(235);
  start_dp_op(234) <= start_cp_ip(236);
  start_dp_op(235) <= start_cp_ip(237);
  start_dp_op(236) <= start_cp_ip(238);
  start_dp_op(237) <= start_cp_ip(239);
  start_dp_op(238) <= start_cp_ip(240);
  start_dp_op(239) <= start_cp_ip(241);
  start_dp_op(240) <= start_cp_ip(242);
  start_dp_op(241) <= start_cp_ip(243);
  start_dp_op(242) <= start_cp_ip(245);
  start_dp_op(243) <= start_cp_ip(244);
  start_dp_op(244) <= start_cp_ip(246);
  start_dp_op(245) <= start_cp_ip(247);
  start_dp_op(246) <= start_cp_ip(248);
  start_dp_op(247) <= start_cp_ip(250);
  start_dp_op(248) <= start_cp_ip(249);
  start_dp_op(249) <= start_cp_ip(252);
  start_dp_op(250) <= start_cp_ip(251);
  start_dp_op(251) <= start_cp_ip(253);
  start_dp_op(252) <= start_cp_ip(254);
  start_dp_op(253) <= start_cp_ip(255);
  start_dp_op(254) <= start_cp_ip(257);
  start_dp_op(255) <= start_cp_ip(256);
  start_dp_op(256) <= start_cp_ip(258);
  start_dp_op(257) <= start_cp_ip(259);
  start_dp_op(258) <= start_cp_ip(260);
  start_dp_op(259) <= start_cp_ip(261);
  start_dp_op(260) <= start_cp_ip(262);
  start_dp_op(261) <= start_cp_ip(263);
  start_dp_op(262) <= start_cp_ip(264);
  start_dp_op(263) <= start_cp_ip(265);
  start_dp_op(264) <= start_cp_ip(266);
  start_dp_op(265) <= start_cp_ip(267);
  start_dp_op(266) <= start_cp_ip(268);
  start_dp_op(267) <= start_cp_ip(269);
  start_dp_op(268) <= start_cp_ip(270);
  start_dp_op(269) <= start_cp_ip(271);
  start_dp_op(270) <= start_cp_ip(272);
  start_dp_op(271) <= start_cp_ip(273);
  start_dp_op(272) <= start_cp_ip(275);
  start_dp_op(273) <= start_cp_ip(274);
  start_dp_op(274) <= start_cp_ip(276);
  start_dp_op(275) <= start_cp_ip(277);
  start_dp_op(276) <= start_cp_ip(278);

end Behavioral;
